module SEControl(
  input  [7:0] io_inst_in,
  output [2:0] io_fu_op,
  output [1:0] io_fu_type,
  output       io_signed
);
  wire  _ctrlSignals_T_1 = 8'h0 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_3 = 8'h4 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_5 = 8'h8 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_7 = 8'h20 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_9 = 8'h24 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_11 = 8'h28 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_13 = 8'h29 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_15 = 8'h80 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_17 = 8'h84 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_19 = 8'h88 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_21 = 8'h40 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_23 = 8'h41 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_25 = 8'h60 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_27 = 8'ha0 == io_inst_in; // @[Lookup.scala 31:38]
  wire  _ctrlSignals_T_29 = 8'hb0 == io_inst_in; // @[Lookup.scala 31:38]
  wire [2:0] _ctrlSignals_T_30 = _ctrlSignals_T_29 ? 3'h5 : 3'h6; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_31 = _ctrlSignals_T_27 ? 3'h5 : _ctrlSignals_T_30; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_32 = _ctrlSignals_T_25 ? 3'h3 : _ctrlSignals_T_31; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_33 = _ctrlSignals_T_23 ? 3'h2 : _ctrlSignals_T_32; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_34 = _ctrlSignals_T_21 ? 3'h2 : _ctrlSignals_T_33; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_35 = _ctrlSignals_T_19 ? 3'h4 : _ctrlSignals_T_34; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_36 = _ctrlSignals_T_17 ? 3'h4 : _ctrlSignals_T_35; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_37 = _ctrlSignals_T_15 ? 3'h4 : _ctrlSignals_T_36; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_38 = _ctrlSignals_T_13 ? 3'h1 : _ctrlSignals_T_37; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_39 = _ctrlSignals_T_11 ? 3'h1 : _ctrlSignals_T_38; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_40 = _ctrlSignals_T_9 ? 3'h1 : _ctrlSignals_T_39; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_41 = _ctrlSignals_T_7 ? 3'h1 : _ctrlSignals_T_40; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_42 = _ctrlSignals_T_5 ? 3'h0 : _ctrlSignals_T_41; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlSignals_T_43 = _ctrlSignals_T_3 ? 3'h0 : _ctrlSignals_T_42; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_44 = _ctrlSignals_T_29 ? 2'h1 : 2'h2; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_45 = _ctrlSignals_T_27 ? 2'h0 : _ctrlSignals_T_44; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_46 = _ctrlSignals_T_25 ? 2'h0 : _ctrlSignals_T_45; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_47 = _ctrlSignals_T_23 ? 2'h0 : _ctrlSignals_T_46; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_48 = _ctrlSignals_T_21 ? 2'h0 : _ctrlSignals_T_47; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_49 = _ctrlSignals_T_19 ? 2'h2 : _ctrlSignals_T_48; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_50 = _ctrlSignals_T_17 ? 2'h1 : _ctrlSignals_T_49; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_51 = _ctrlSignals_T_15 ? 2'h0 : _ctrlSignals_T_50; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_52 = _ctrlSignals_T_13 ? 2'h2 : _ctrlSignals_T_51; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_53 = _ctrlSignals_T_11 ? 2'h2 : _ctrlSignals_T_52; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_54 = _ctrlSignals_T_9 ? 2'h1 : _ctrlSignals_T_53; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_55 = _ctrlSignals_T_7 ? 2'h0 : _ctrlSignals_T_54; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_56 = _ctrlSignals_T_5 ? 2'h2 : _ctrlSignals_T_55; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlSignals_T_57 = _ctrlSignals_T_3 ? 2'h1 : _ctrlSignals_T_56; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_76 = _ctrlSignals_T_21 ? 1'h0 : _ctrlSignals_T_23; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_77 = _ctrlSignals_T_19 ? 1'h0 : _ctrlSignals_T_76; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_78 = _ctrlSignals_T_17 ? 1'h0 : _ctrlSignals_T_77; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_79 = _ctrlSignals_T_15 ? 1'h0 : _ctrlSignals_T_78; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_81 = _ctrlSignals_T_11 ? 1'h0 : _ctrlSignals_T_13 | _ctrlSignals_T_79; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_82 = _ctrlSignals_T_9 ? 1'h0 : _ctrlSignals_T_81; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_83 = _ctrlSignals_T_7 ? 1'h0 : _ctrlSignals_T_82; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_84 = _ctrlSignals_T_5 ? 1'h0 : _ctrlSignals_T_83; // @[Lookup.scala 34:39]
  wire  _ctrlSignals_T_85 = _ctrlSignals_T_3 ? 1'h0 : _ctrlSignals_T_84; // @[Lookup.scala 34:39]
  assign io_fu_op = _ctrlSignals_T_1 ? 3'h0 : _ctrlSignals_T_43; // @[Lookup.scala 34:39]
  assign io_fu_type = _ctrlSignals_T_1 ? 2'h0 : _ctrlSignals_T_57; // @[Lookup.scala 34:39]
  assign io_signed = _ctrlSignals_T_1 ? 1'h0 : _ctrlSignals_T_85; // @[Lookup.scala 34:39]
endmodule
module FU(
  input  [63:0] io_A,
  input  [63:0] io_B,
  input  [2:0]  io_fu_op,
  input  [1:0]  io_fu_type,
  input         io_signed,
  output [63:0] io_out
);
  wire  _T_1 = io_fu_type == 2'h0; // @[FU.scala 45:21]
  wire [126:0] _GEN_15 = {{63'd0}, io_A}; // @[FU.scala 47:22]
  wire [126:0] _output_T_1 = _GEN_15 << io_B[5:0]; // @[FU.scala 47:22]
  wire  _T_2 = io_fu_type == 2'h1; // @[FU.scala 48:27]
  wire [63:0] _output_T_3 = io_A >> io_B[5:0]; // @[FU.scala 50:22]
  wire [63:0] _output_T_7 = $signed(io_A) >>> io_B[5:0]; // @[FU.scala 53:43]
  wire [63:0] _output_T_9 = {io_A[63],_output_T_7[62:0]}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_0 = io_fu_type == 2'h1 ? _output_T_3 : _output_T_9; // @[FU.scala 48:41 50:14 53:14]
  wire [126:0] _GEN_1 = io_fu_type == 2'h0 ? _output_T_1 : {{63'd0}, _GEN_0}; // @[FU.scala 45:35 47:14]
  wire [127:0] _output_T_13 = $signed(io_A) * $signed(io_B); // @[FU.scala 58:47]
  wire [63:0] _output_T_15 = io_A + io_B; // @[FU.scala 62:24]
  wire [63:0] _output_T_17 = io_A - io_B; // @[FU.scala 65:24]
  wire [127:0] _output_T_18 = io_A * io_B; // @[FU.scala 68:24]
  wire [127:0] _GEN_2 = _T_2 ? {{64'd0}, _output_T_17} : _output_T_18; // @[FU.scala 63:43 65:16 68:16]
  wire [127:0] _GEN_3 = _T_1 ? {{64'd0}, _output_T_15} : _GEN_2; // @[FU.scala 60:37 62:16]
  wire [127:0] _GEN_4 = io_signed ? _output_T_13 : _GEN_3; // @[FU.scala 56:20 58:16]
  wire [63:0] _output_T_19 = io_A ^ io_B; // @[FU.scala 74:24]
  wire [63:0] _output_T_20 = io_A | io_B; // @[FU.scala 77:24]
  wire [63:0] _output_T_21 = io_A & io_B; // @[FU.scala 80:24]
  wire [63:0] _GEN_5 = _T_2 ? _output_T_20 : _output_T_21; // @[FU.scala 75:44 77:16 80:16]
  wire [63:0] _GEN_6 = _T_1 ? _output_T_19 : _GEN_5; // @[FU.scala 72:39 74:16]
  wire  _GEN_7 = io_signed ? $signed(io_A) < $signed(io_B) : io_A < io_B; // @[FU.scala 83:20 85:14 88:14]
  wire [2:0] _GEN_14 = {{1'd0}, io_fu_type}; // @[FU.scala 90:25]
  wire [63:0] _GEN_8 = io_A != 64'h0 ? io_B : 64'h0; // @[FU.scala 91:23 93:14 96:14]
  wire [63:0] _GEN_9 = _GEN_14 == 3'h3 ? _GEN_8 : io_A; // @[FU.scala 100:14 90:37]
  wire [63:0] _GEN_10 = io_fu_op == 3'h2 ? {{63'd0}, _GEN_7} : _GEN_9; // @[FU.scala 82:35]
  wire [63:0] _GEN_11 = io_fu_op == 3'h4 ? _GEN_6 : _GEN_10; // @[FU.scala 71:38]
  wire [127:0] _GEN_12 = io_fu_op == 3'h1 ? _GEN_4 : {{64'd0}, _GEN_11}; // @[FU.scala 55:36]
  wire [127:0] _GEN_13 = io_fu_op == 3'h0 ? {{1'd0}, _GEN_1} : _GEN_12; // @[FU.scala 44:30]
  assign io_out = _GEN_13[63:0]; // @[FU.scala 42:20]
endmodule
module SEOperation(
  input  [7:0]  io_inst,
  input         io_in_valid,
  input  [63:0] io_op1_input,
  input  [63:0] io_op2_input,
  output [63:0] io_result,
  output        io_out_valid
);
  wire [7:0] decode_io_inst_in; // @[SEOperation.scala 31:28]
  wire [2:0] decode_io_fu_op; // @[SEOperation.scala 31:28]
  wire [1:0] decode_io_fu_type; // @[SEOperation.scala 31:28]
  wire  decode_io_signed; // @[SEOperation.scala 31:28]
  wire [63:0] fu_io_A; // @[SEOperation.scala 32:24]
  wire [63:0] fu_io_B; // @[SEOperation.scala 32:24]
  wire [2:0] fu_io_fu_op; // @[SEOperation.scala 32:24]
  wire [1:0] fu_io_fu_type; // @[SEOperation.scala 32:24]
  wire  fu_io_signed; // @[SEOperation.scala 32:24]
  wire [63:0] fu_io_out; // @[SEOperation.scala 32:24]
  SEControl decode ( // @[SEOperation.scala 31:28]
    .io_inst_in(decode_io_inst_in),
    .io_fu_op(decode_io_fu_op),
    .io_fu_type(decode_io_fu_type),
    .io_signed(decode_io_signed)
  );
  FU fu ( // @[SEOperation.scala 32:24]
    .io_A(fu_io_A),
    .io_B(fu_io_B),
    .io_fu_op(fu_io_fu_op),
    .io_fu_type(fu_io_fu_type),
    .io_signed(fu_io_signed),
    .io_out(fu_io_out)
  );
  assign io_result = fu_io_out; // @[SEOperation.scala 45:19]
  assign io_out_valid = io_in_valid; // @[SEOperation.scala 46:22]
  assign decode_io_inst_in = io_inst; // @[SEOperation.scala 37:27]
  assign fu_io_A = io_op1_input; // @[SEOperation.scala 40:11]
  assign fu_io_B = io_op2_input; // @[SEOperation.scala 41:11]
  assign fu_io_fu_op = decode_io_fu_op; // @[SEOperation.scala 42:15]
  assign fu_io_fu_type = decode_io_fu_type; // @[SEOperation.scala 43:23]
  assign fu_io_signed = decode_io_signed; // @[SEOperation.scala 44:22]
endmodule
module AddRoundKey(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  input  [7:0] io_roundKey_0,
  input  [7:0] io_roundKey_1,
  input  [7:0] io_roundKey_2,
  input  [7:0] io_roundKey_3,
  input  [7:0] io_roundKey_4,
  input  [7:0] io_roundKey_5,
  input  [7:0] io_roundKey_6,
  input  [7:0] io_roundKey_7,
  input  [7:0] io_roundKey_8,
  input  [7:0] io_roundKey_9,
  input  [7:0] io_roundKey_10,
  input  [7:0] io_roundKey_11,
  input  [7:0] io_roundKey_12,
  input  [7:0] io_roundKey_13,
  input  [7:0] io_roundKey_14,
  input  [7:0] io_roundKey_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  assign io_state_out_0 = io_state_in_0 ^ io_roundKey_0; // @[AddRoundKey.scala 19:41]
  assign io_state_out_1 = io_state_in_1 ^ io_roundKey_1; // @[AddRoundKey.scala 19:41]
  assign io_state_out_2 = io_state_in_2 ^ io_roundKey_2; // @[AddRoundKey.scala 19:41]
  assign io_state_out_3 = io_state_in_3 ^ io_roundKey_3; // @[AddRoundKey.scala 19:41]
  assign io_state_out_4 = io_state_in_4 ^ io_roundKey_4; // @[AddRoundKey.scala 19:41]
  assign io_state_out_5 = io_state_in_5 ^ io_roundKey_5; // @[AddRoundKey.scala 19:41]
  assign io_state_out_6 = io_state_in_6 ^ io_roundKey_6; // @[AddRoundKey.scala 19:41]
  assign io_state_out_7 = io_state_in_7 ^ io_roundKey_7; // @[AddRoundKey.scala 19:41]
  assign io_state_out_8 = io_state_in_8 ^ io_roundKey_8; // @[AddRoundKey.scala 19:41]
  assign io_state_out_9 = io_state_in_9 ^ io_roundKey_9; // @[AddRoundKey.scala 19:41]
  assign io_state_out_10 = io_state_in_10 ^ io_roundKey_10; // @[AddRoundKey.scala 19:41]
  assign io_state_out_11 = io_state_in_11 ^ io_roundKey_11; // @[AddRoundKey.scala 19:41]
  assign io_state_out_12 = io_state_in_12 ^ io_roundKey_12; // @[AddRoundKey.scala 19:41]
  assign io_state_out_13 = io_state_in_13 ^ io_roundKey_13; // @[AddRoundKey.scala 19:41]
  assign io_state_out_14 = io_state_in_14 ^ io_roundKey_14; // @[AddRoundKey.scala 19:41]
  assign io_state_out_15 = io_state_in_15 ^ io_roundKey_15; // @[AddRoundKey.scala 19:41]
endmodule
module InvSubBytes(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  wire [7:0] _GEN_1 = 8'h1 == io_state_in_0 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2 = 8'h2 == io_state_in_0 ? 8'h6a : _GEN_1; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3 = 8'h3 == io_state_in_0 ? 8'hd5 : _GEN_2; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4 = 8'h4 == io_state_in_0 ? 8'h30 : _GEN_3; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_5 = 8'h5 == io_state_in_0 ? 8'h36 : _GEN_4; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_6 = 8'h6 == io_state_in_0 ? 8'ha5 : _GEN_5; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_7 = 8'h7 == io_state_in_0 ? 8'h38 : _GEN_6; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_8 = 8'h8 == io_state_in_0 ? 8'hbf : _GEN_7; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_9 = 8'h9 == io_state_in_0 ? 8'h40 : _GEN_8; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_10 = 8'ha == io_state_in_0 ? 8'ha3 : _GEN_9; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_11 = 8'hb == io_state_in_0 ? 8'h9e : _GEN_10; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_12 = 8'hc == io_state_in_0 ? 8'h81 : _GEN_11; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_13 = 8'hd == io_state_in_0 ? 8'hf3 : _GEN_12; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_14 = 8'he == io_state_in_0 ? 8'hd7 : _GEN_13; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_15 = 8'hf == io_state_in_0 ? 8'hfb : _GEN_14; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_16 = 8'h10 == io_state_in_0 ? 8'h7c : _GEN_15; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_17 = 8'h11 == io_state_in_0 ? 8'he3 : _GEN_16; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_18 = 8'h12 == io_state_in_0 ? 8'h39 : _GEN_17; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_19 = 8'h13 == io_state_in_0 ? 8'h82 : _GEN_18; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_20 = 8'h14 == io_state_in_0 ? 8'h9b : _GEN_19; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_21 = 8'h15 == io_state_in_0 ? 8'h2f : _GEN_20; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_22 = 8'h16 == io_state_in_0 ? 8'hff : _GEN_21; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_23 = 8'h17 == io_state_in_0 ? 8'h87 : _GEN_22; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_24 = 8'h18 == io_state_in_0 ? 8'h34 : _GEN_23; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_25 = 8'h19 == io_state_in_0 ? 8'h8e : _GEN_24; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_26 = 8'h1a == io_state_in_0 ? 8'h43 : _GEN_25; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_27 = 8'h1b == io_state_in_0 ? 8'h44 : _GEN_26; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_28 = 8'h1c == io_state_in_0 ? 8'hc4 : _GEN_27; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_29 = 8'h1d == io_state_in_0 ? 8'hde : _GEN_28; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_30 = 8'h1e == io_state_in_0 ? 8'he9 : _GEN_29; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_31 = 8'h1f == io_state_in_0 ? 8'hcb : _GEN_30; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_32 = 8'h20 == io_state_in_0 ? 8'h54 : _GEN_31; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_33 = 8'h21 == io_state_in_0 ? 8'h7b : _GEN_32; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_34 = 8'h22 == io_state_in_0 ? 8'h94 : _GEN_33; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_35 = 8'h23 == io_state_in_0 ? 8'h32 : _GEN_34; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_36 = 8'h24 == io_state_in_0 ? 8'ha6 : _GEN_35; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_37 = 8'h25 == io_state_in_0 ? 8'hc2 : _GEN_36; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_38 = 8'h26 == io_state_in_0 ? 8'h23 : _GEN_37; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_39 = 8'h27 == io_state_in_0 ? 8'h3d : _GEN_38; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_40 = 8'h28 == io_state_in_0 ? 8'hee : _GEN_39; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_41 = 8'h29 == io_state_in_0 ? 8'h4c : _GEN_40; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_42 = 8'h2a == io_state_in_0 ? 8'h95 : _GEN_41; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_43 = 8'h2b == io_state_in_0 ? 8'hb : _GEN_42; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_44 = 8'h2c == io_state_in_0 ? 8'h42 : _GEN_43; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_45 = 8'h2d == io_state_in_0 ? 8'hfa : _GEN_44; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_46 = 8'h2e == io_state_in_0 ? 8'hc3 : _GEN_45; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_47 = 8'h2f == io_state_in_0 ? 8'h4e : _GEN_46; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_48 = 8'h30 == io_state_in_0 ? 8'h8 : _GEN_47; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_49 = 8'h31 == io_state_in_0 ? 8'h2e : _GEN_48; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_50 = 8'h32 == io_state_in_0 ? 8'ha1 : _GEN_49; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_51 = 8'h33 == io_state_in_0 ? 8'h66 : _GEN_50; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_52 = 8'h34 == io_state_in_0 ? 8'h28 : _GEN_51; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_53 = 8'h35 == io_state_in_0 ? 8'hd9 : _GEN_52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_54 = 8'h36 == io_state_in_0 ? 8'h24 : _GEN_53; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_55 = 8'h37 == io_state_in_0 ? 8'hb2 : _GEN_54; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_56 = 8'h38 == io_state_in_0 ? 8'h76 : _GEN_55; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_57 = 8'h39 == io_state_in_0 ? 8'h5b : _GEN_56; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_58 = 8'h3a == io_state_in_0 ? 8'ha2 : _GEN_57; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_59 = 8'h3b == io_state_in_0 ? 8'h49 : _GEN_58; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_60 = 8'h3c == io_state_in_0 ? 8'h6d : _GEN_59; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_61 = 8'h3d == io_state_in_0 ? 8'h8b : _GEN_60; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_62 = 8'h3e == io_state_in_0 ? 8'hd1 : _GEN_61; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_63 = 8'h3f == io_state_in_0 ? 8'h25 : _GEN_62; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_64 = 8'h40 == io_state_in_0 ? 8'h72 : _GEN_63; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_65 = 8'h41 == io_state_in_0 ? 8'hf8 : _GEN_64; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_66 = 8'h42 == io_state_in_0 ? 8'hf6 : _GEN_65; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_67 = 8'h43 == io_state_in_0 ? 8'h64 : _GEN_66; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_68 = 8'h44 == io_state_in_0 ? 8'h86 : _GEN_67; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_69 = 8'h45 == io_state_in_0 ? 8'h68 : _GEN_68; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_70 = 8'h46 == io_state_in_0 ? 8'h98 : _GEN_69; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_71 = 8'h47 == io_state_in_0 ? 8'h16 : _GEN_70; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_72 = 8'h48 == io_state_in_0 ? 8'hd4 : _GEN_71; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_73 = 8'h49 == io_state_in_0 ? 8'ha4 : _GEN_72; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_74 = 8'h4a == io_state_in_0 ? 8'h5c : _GEN_73; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_75 = 8'h4b == io_state_in_0 ? 8'hcc : _GEN_74; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_76 = 8'h4c == io_state_in_0 ? 8'h5d : _GEN_75; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_77 = 8'h4d == io_state_in_0 ? 8'h65 : _GEN_76; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_78 = 8'h4e == io_state_in_0 ? 8'hb6 : _GEN_77; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_79 = 8'h4f == io_state_in_0 ? 8'h92 : _GEN_78; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_80 = 8'h50 == io_state_in_0 ? 8'h6c : _GEN_79; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_81 = 8'h51 == io_state_in_0 ? 8'h70 : _GEN_80; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_82 = 8'h52 == io_state_in_0 ? 8'h48 : _GEN_81; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_83 = 8'h53 == io_state_in_0 ? 8'h50 : _GEN_82; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_84 = 8'h54 == io_state_in_0 ? 8'hfd : _GEN_83; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_85 = 8'h55 == io_state_in_0 ? 8'hed : _GEN_84; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_86 = 8'h56 == io_state_in_0 ? 8'hb9 : _GEN_85; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_87 = 8'h57 == io_state_in_0 ? 8'hda : _GEN_86; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_88 = 8'h58 == io_state_in_0 ? 8'h5e : _GEN_87; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_89 = 8'h59 == io_state_in_0 ? 8'h15 : _GEN_88; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_90 = 8'h5a == io_state_in_0 ? 8'h46 : _GEN_89; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_91 = 8'h5b == io_state_in_0 ? 8'h57 : _GEN_90; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_92 = 8'h5c == io_state_in_0 ? 8'ha7 : _GEN_91; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_93 = 8'h5d == io_state_in_0 ? 8'h8d : _GEN_92; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_94 = 8'h5e == io_state_in_0 ? 8'h9d : _GEN_93; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_95 = 8'h5f == io_state_in_0 ? 8'h84 : _GEN_94; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_96 = 8'h60 == io_state_in_0 ? 8'h90 : _GEN_95; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_97 = 8'h61 == io_state_in_0 ? 8'hd8 : _GEN_96; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_98 = 8'h62 == io_state_in_0 ? 8'hab : _GEN_97; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_99 = 8'h63 == io_state_in_0 ? 8'h0 : _GEN_98; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_100 = 8'h64 == io_state_in_0 ? 8'h8c : _GEN_99; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_101 = 8'h65 == io_state_in_0 ? 8'hbc : _GEN_100; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_102 = 8'h66 == io_state_in_0 ? 8'hd3 : _GEN_101; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_103 = 8'h67 == io_state_in_0 ? 8'ha : _GEN_102; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_104 = 8'h68 == io_state_in_0 ? 8'hf7 : _GEN_103; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_105 = 8'h69 == io_state_in_0 ? 8'he4 : _GEN_104; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_106 = 8'h6a == io_state_in_0 ? 8'h58 : _GEN_105; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_107 = 8'h6b == io_state_in_0 ? 8'h5 : _GEN_106; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_108 = 8'h6c == io_state_in_0 ? 8'hb8 : _GEN_107; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_109 = 8'h6d == io_state_in_0 ? 8'hb3 : _GEN_108; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_110 = 8'h6e == io_state_in_0 ? 8'h45 : _GEN_109; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_111 = 8'h6f == io_state_in_0 ? 8'h6 : _GEN_110; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_112 = 8'h70 == io_state_in_0 ? 8'hd0 : _GEN_111; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_113 = 8'h71 == io_state_in_0 ? 8'h2c : _GEN_112; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_114 = 8'h72 == io_state_in_0 ? 8'h1e : _GEN_113; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_115 = 8'h73 == io_state_in_0 ? 8'h8f : _GEN_114; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_116 = 8'h74 == io_state_in_0 ? 8'hca : _GEN_115; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_117 = 8'h75 == io_state_in_0 ? 8'h3f : _GEN_116; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_118 = 8'h76 == io_state_in_0 ? 8'hf : _GEN_117; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_119 = 8'h77 == io_state_in_0 ? 8'h2 : _GEN_118; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_120 = 8'h78 == io_state_in_0 ? 8'hc1 : _GEN_119; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_121 = 8'h79 == io_state_in_0 ? 8'haf : _GEN_120; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_122 = 8'h7a == io_state_in_0 ? 8'hbd : _GEN_121; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_123 = 8'h7b == io_state_in_0 ? 8'h3 : _GEN_122; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_124 = 8'h7c == io_state_in_0 ? 8'h1 : _GEN_123; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_125 = 8'h7d == io_state_in_0 ? 8'h13 : _GEN_124; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_126 = 8'h7e == io_state_in_0 ? 8'h8a : _GEN_125; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_127 = 8'h7f == io_state_in_0 ? 8'h6b : _GEN_126; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_128 = 8'h80 == io_state_in_0 ? 8'h3a : _GEN_127; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_129 = 8'h81 == io_state_in_0 ? 8'h91 : _GEN_128; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_130 = 8'h82 == io_state_in_0 ? 8'h11 : _GEN_129; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_131 = 8'h83 == io_state_in_0 ? 8'h41 : _GEN_130; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_132 = 8'h84 == io_state_in_0 ? 8'h4f : _GEN_131; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_133 = 8'h85 == io_state_in_0 ? 8'h67 : _GEN_132; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_134 = 8'h86 == io_state_in_0 ? 8'hdc : _GEN_133; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_135 = 8'h87 == io_state_in_0 ? 8'hea : _GEN_134; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_136 = 8'h88 == io_state_in_0 ? 8'h97 : _GEN_135; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_137 = 8'h89 == io_state_in_0 ? 8'hf2 : _GEN_136; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_138 = 8'h8a == io_state_in_0 ? 8'hcf : _GEN_137; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_139 = 8'h8b == io_state_in_0 ? 8'hce : _GEN_138; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_140 = 8'h8c == io_state_in_0 ? 8'hf0 : _GEN_139; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_141 = 8'h8d == io_state_in_0 ? 8'hb4 : _GEN_140; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_142 = 8'h8e == io_state_in_0 ? 8'he6 : _GEN_141; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_143 = 8'h8f == io_state_in_0 ? 8'h73 : _GEN_142; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_144 = 8'h90 == io_state_in_0 ? 8'h96 : _GEN_143; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_145 = 8'h91 == io_state_in_0 ? 8'hac : _GEN_144; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_146 = 8'h92 == io_state_in_0 ? 8'h74 : _GEN_145; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_147 = 8'h93 == io_state_in_0 ? 8'h22 : _GEN_146; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_148 = 8'h94 == io_state_in_0 ? 8'he7 : _GEN_147; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_149 = 8'h95 == io_state_in_0 ? 8'had : _GEN_148; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_150 = 8'h96 == io_state_in_0 ? 8'h35 : _GEN_149; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_151 = 8'h97 == io_state_in_0 ? 8'h85 : _GEN_150; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_152 = 8'h98 == io_state_in_0 ? 8'he2 : _GEN_151; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_153 = 8'h99 == io_state_in_0 ? 8'hf9 : _GEN_152; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_154 = 8'h9a == io_state_in_0 ? 8'h37 : _GEN_153; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_155 = 8'h9b == io_state_in_0 ? 8'he8 : _GEN_154; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_156 = 8'h9c == io_state_in_0 ? 8'h1c : _GEN_155; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_157 = 8'h9d == io_state_in_0 ? 8'h75 : _GEN_156; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_158 = 8'h9e == io_state_in_0 ? 8'hdf : _GEN_157; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_159 = 8'h9f == io_state_in_0 ? 8'h6e : _GEN_158; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_160 = 8'ha0 == io_state_in_0 ? 8'h47 : _GEN_159; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_161 = 8'ha1 == io_state_in_0 ? 8'hf1 : _GEN_160; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_162 = 8'ha2 == io_state_in_0 ? 8'h1a : _GEN_161; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_163 = 8'ha3 == io_state_in_0 ? 8'h71 : _GEN_162; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_164 = 8'ha4 == io_state_in_0 ? 8'h1d : _GEN_163; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_165 = 8'ha5 == io_state_in_0 ? 8'h29 : _GEN_164; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_166 = 8'ha6 == io_state_in_0 ? 8'hc5 : _GEN_165; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_167 = 8'ha7 == io_state_in_0 ? 8'h89 : _GEN_166; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_168 = 8'ha8 == io_state_in_0 ? 8'h6f : _GEN_167; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_169 = 8'ha9 == io_state_in_0 ? 8'hb7 : _GEN_168; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_170 = 8'haa == io_state_in_0 ? 8'h62 : _GEN_169; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_171 = 8'hab == io_state_in_0 ? 8'he : _GEN_170; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_172 = 8'hac == io_state_in_0 ? 8'haa : _GEN_171; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_173 = 8'had == io_state_in_0 ? 8'h18 : _GEN_172; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_174 = 8'hae == io_state_in_0 ? 8'hbe : _GEN_173; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_175 = 8'haf == io_state_in_0 ? 8'h1b : _GEN_174; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_176 = 8'hb0 == io_state_in_0 ? 8'hfc : _GEN_175; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_177 = 8'hb1 == io_state_in_0 ? 8'h56 : _GEN_176; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_178 = 8'hb2 == io_state_in_0 ? 8'h3e : _GEN_177; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_179 = 8'hb3 == io_state_in_0 ? 8'h4b : _GEN_178; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_180 = 8'hb4 == io_state_in_0 ? 8'hc6 : _GEN_179; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_181 = 8'hb5 == io_state_in_0 ? 8'hd2 : _GEN_180; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_182 = 8'hb6 == io_state_in_0 ? 8'h79 : _GEN_181; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_183 = 8'hb7 == io_state_in_0 ? 8'h20 : _GEN_182; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_184 = 8'hb8 == io_state_in_0 ? 8'h9a : _GEN_183; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_185 = 8'hb9 == io_state_in_0 ? 8'hdb : _GEN_184; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_186 = 8'hba == io_state_in_0 ? 8'hc0 : _GEN_185; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_187 = 8'hbb == io_state_in_0 ? 8'hfe : _GEN_186; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_188 = 8'hbc == io_state_in_0 ? 8'h78 : _GEN_187; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_189 = 8'hbd == io_state_in_0 ? 8'hcd : _GEN_188; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_190 = 8'hbe == io_state_in_0 ? 8'h5a : _GEN_189; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_191 = 8'hbf == io_state_in_0 ? 8'hf4 : _GEN_190; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_192 = 8'hc0 == io_state_in_0 ? 8'h1f : _GEN_191; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_193 = 8'hc1 == io_state_in_0 ? 8'hdd : _GEN_192; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_194 = 8'hc2 == io_state_in_0 ? 8'ha8 : _GEN_193; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_195 = 8'hc3 == io_state_in_0 ? 8'h33 : _GEN_194; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_196 = 8'hc4 == io_state_in_0 ? 8'h88 : _GEN_195; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_197 = 8'hc5 == io_state_in_0 ? 8'h7 : _GEN_196; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_198 = 8'hc6 == io_state_in_0 ? 8'hc7 : _GEN_197; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_199 = 8'hc7 == io_state_in_0 ? 8'h31 : _GEN_198; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_200 = 8'hc8 == io_state_in_0 ? 8'hb1 : _GEN_199; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_201 = 8'hc9 == io_state_in_0 ? 8'h12 : _GEN_200; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_202 = 8'hca == io_state_in_0 ? 8'h10 : _GEN_201; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_203 = 8'hcb == io_state_in_0 ? 8'h59 : _GEN_202; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_204 = 8'hcc == io_state_in_0 ? 8'h27 : _GEN_203; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_205 = 8'hcd == io_state_in_0 ? 8'h80 : _GEN_204; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_206 = 8'hce == io_state_in_0 ? 8'hec : _GEN_205; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_207 = 8'hcf == io_state_in_0 ? 8'h5f : _GEN_206; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_208 = 8'hd0 == io_state_in_0 ? 8'h60 : _GEN_207; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_209 = 8'hd1 == io_state_in_0 ? 8'h51 : _GEN_208; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_210 = 8'hd2 == io_state_in_0 ? 8'h7f : _GEN_209; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_211 = 8'hd3 == io_state_in_0 ? 8'ha9 : _GEN_210; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_212 = 8'hd4 == io_state_in_0 ? 8'h19 : _GEN_211; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_213 = 8'hd5 == io_state_in_0 ? 8'hb5 : _GEN_212; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_214 = 8'hd6 == io_state_in_0 ? 8'h4a : _GEN_213; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_215 = 8'hd7 == io_state_in_0 ? 8'hd : _GEN_214; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_216 = 8'hd8 == io_state_in_0 ? 8'h2d : _GEN_215; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_217 = 8'hd9 == io_state_in_0 ? 8'he5 : _GEN_216; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_218 = 8'hda == io_state_in_0 ? 8'h7a : _GEN_217; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_219 = 8'hdb == io_state_in_0 ? 8'h9f : _GEN_218; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_220 = 8'hdc == io_state_in_0 ? 8'h93 : _GEN_219; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_221 = 8'hdd == io_state_in_0 ? 8'hc9 : _GEN_220; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_222 = 8'hde == io_state_in_0 ? 8'h9c : _GEN_221; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_223 = 8'hdf == io_state_in_0 ? 8'hef : _GEN_222; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_224 = 8'he0 == io_state_in_0 ? 8'ha0 : _GEN_223; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_225 = 8'he1 == io_state_in_0 ? 8'he0 : _GEN_224; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_226 = 8'he2 == io_state_in_0 ? 8'h3b : _GEN_225; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_227 = 8'he3 == io_state_in_0 ? 8'h4d : _GEN_226; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_228 = 8'he4 == io_state_in_0 ? 8'hae : _GEN_227; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_229 = 8'he5 == io_state_in_0 ? 8'h2a : _GEN_228; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_230 = 8'he6 == io_state_in_0 ? 8'hf5 : _GEN_229; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_231 = 8'he7 == io_state_in_0 ? 8'hb0 : _GEN_230; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_232 = 8'he8 == io_state_in_0 ? 8'hc8 : _GEN_231; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_233 = 8'he9 == io_state_in_0 ? 8'heb : _GEN_232; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_234 = 8'hea == io_state_in_0 ? 8'hbb : _GEN_233; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_235 = 8'heb == io_state_in_0 ? 8'h3c : _GEN_234; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_236 = 8'hec == io_state_in_0 ? 8'h83 : _GEN_235; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_237 = 8'hed == io_state_in_0 ? 8'h53 : _GEN_236; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_238 = 8'hee == io_state_in_0 ? 8'h99 : _GEN_237; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_239 = 8'hef == io_state_in_0 ? 8'h61 : _GEN_238; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_240 = 8'hf0 == io_state_in_0 ? 8'h17 : _GEN_239; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_241 = 8'hf1 == io_state_in_0 ? 8'h2b : _GEN_240; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_242 = 8'hf2 == io_state_in_0 ? 8'h4 : _GEN_241; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_243 = 8'hf3 == io_state_in_0 ? 8'h7e : _GEN_242; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_244 = 8'hf4 == io_state_in_0 ? 8'hba : _GEN_243; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_245 = 8'hf5 == io_state_in_0 ? 8'h77 : _GEN_244; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_246 = 8'hf6 == io_state_in_0 ? 8'hd6 : _GEN_245; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_247 = 8'hf7 == io_state_in_0 ? 8'h26 : _GEN_246; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_248 = 8'hf8 == io_state_in_0 ? 8'he1 : _GEN_247; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_249 = 8'hf9 == io_state_in_0 ? 8'h69 : _GEN_248; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_250 = 8'hfa == io_state_in_0 ? 8'h14 : _GEN_249; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_251 = 8'hfb == io_state_in_0 ? 8'h63 : _GEN_250; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_252 = 8'hfc == io_state_in_0 ? 8'h55 : _GEN_251; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_253 = 8'hfd == io_state_in_0 ? 8'h21 : _GEN_252; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_254 = 8'hfe == io_state_in_0 ? 8'hc : _GEN_253; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_257 = 8'h1 == io_state_in_1 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_258 = 8'h2 == io_state_in_1 ? 8'h6a : _GEN_257; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_259 = 8'h3 == io_state_in_1 ? 8'hd5 : _GEN_258; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_260 = 8'h4 == io_state_in_1 ? 8'h30 : _GEN_259; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_261 = 8'h5 == io_state_in_1 ? 8'h36 : _GEN_260; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_262 = 8'h6 == io_state_in_1 ? 8'ha5 : _GEN_261; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_263 = 8'h7 == io_state_in_1 ? 8'h38 : _GEN_262; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_264 = 8'h8 == io_state_in_1 ? 8'hbf : _GEN_263; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_265 = 8'h9 == io_state_in_1 ? 8'h40 : _GEN_264; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_266 = 8'ha == io_state_in_1 ? 8'ha3 : _GEN_265; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_267 = 8'hb == io_state_in_1 ? 8'h9e : _GEN_266; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_268 = 8'hc == io_state_in_1 ? 8'h81 : _GEN_267; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_269 = 8'hd == io_state_in_1 ? 8'hf3 : _GEN_268; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_270 = 8'he == io_state_in_1 ? 8'hd7 : _GEN_269; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_271 = 8'hf == io_state_in_1 ? 8'hfb : _GEN_270; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_272 = 8'h10 == io_state_in_1 ? 8'h7c : _GEN_271; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_273 = 8'h11 == io_state_in_1 ? 8'he3 : _GEN_272; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_274 = 8'h12 == io_state_in_1 ? 8'h39 : _GEN_273; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_275 = 8'h13 == io_state_in_1 ? 8'h82 : _GEN_274; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_276 = 8'h14 == io_state_in_1 ? 8'h9b : _GEN_275; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_277 = 8'h15 == io_state_in_1 ? 8'h2f : _GEN_276; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_278 = 8'h16 == io_state_in_1 ? 8'hff : _GEN_277; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_279 = 8'h17 == io_state_in_1 ? 8'h87 : _GEN_278; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_280 = 8'h18 == io_state_in_1 ? 8'h34 : _GEN_279; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_281 = 8'h19 == io_state_in_1 ? 8'h8e : _GEN_280; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_282 = 8'h1a == io_state_in_1 ? 8'h43 : _GEN_281; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_283 = 8'h1b == io_state_in_1 ? 8'h44 : _GEN_282; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_284 = 8'h1c == io_state_in_1 ? 8'hc4 : _GEN_283; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_285 = 8'h1d == io_state_in_1 ? 8'hde : _GEN_284; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_286 = 8'h1e == io_state_in_1 ? 8'he9 : _GEN_285; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_287 = 8'h1f == io_state_in_1 ? 8'hcb : _GEN_286; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_288 = 8'h20 == io_state_in_1 ? 8'h54 : _GEN_287; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_289 = 8'h21 == io_state_in_1 ? 8'h7b : _GEN_288; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_290 = 8'h22 == io_state_in_1 ? 8'h94 : _GEN_289; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_291 = 8'h23 == io_state_in_1 ? 8'h32 : _GEN_290; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_292 = 8'h24 == io_state_in_1 ? 8'ha6 : _GEN_291; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_293 = 8'h25 == io_state_in_1 ? 8'hc2 : _GEN_292; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_294 = 8'h26 == io_state_in_1 ? 8'h23 : _GEN_293; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_295 = 8'h27 == io_state_in_1 ? 8'h3d : _GEN_294; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_296 = 8'h28 == io_state_in_1 ? 8'hee : _GEN_295; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_297 = 8'h29 == io_state_in_1 ? 8'h4c : _GEN_296; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_298 = 8'h2a == io_state_in_1 ? 8'h95 : _GEN_297; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_299 = 8'h2b == io_state_in_1 ? 8'hb : _GEN_298; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_300 = 8'h2c == io_state_in_1 ? 8'h42 : _GEN_299; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_301 = 8'h2d == io_state_in_1 ? 8'hfa : _GEN_300; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_302 = 8'h2e == io_state_in_1 ? 8'hc3 : _GEN_301; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_303 = 8'h2f == io_state_in_1 ? 8'h4e : _GEN_302; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_304 = 8'h30 == io_state_in_1 ? 8'h8 : _GEN_303; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_305 = 8'h31 == io_state_in_1 ? 8'h2e : _GEN_304; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_306 = 8'h32 == io_state_in_1 ? 8'ha1 : _GEN_305; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_307 = 8'h33 == io_state_in_1 ? 8'h66 : _GEN_306; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_308 = 8'h34 == io_state_in_1 ? 8'h28 : _GEN_307; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_309 = 8'h35 == io_state_in_1 ? 8'hd9 : _GEN_308; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_310 = 8'h36 == io_state_in_1 ? 8'h24 : _GEN_309; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_311 = 8'h37 == io_state_in_1 ? 8'hb2 : _GEN_310; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_312 = 8'h38 == io_state_in_1 ? 8'h76 : _GEN_311; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_313 = 8'h39 == io_state_in_1 ? 8'h5b : _GEN_312; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_314 = 8'h3a == io_state_in_1 ? 8'ha2 : _GEN_313; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_315 = 8'h3b == io_state_in_1 ? 8'h49 : _GEN_314; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_316 = 8'h3c == io_state_in_1 ? 8'h6d : _GEN_315; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_317 = 8'h3d == io_state_in_1 ? 8'h8b : _GEN_316; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_318 = 8'h3e == io_state_in_1 ? 8'hd1 : _GEN_317; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_319 = 8'h3f == io_state_in_1 ? 8'h25 : _GEN_318; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_320 = 8'h40 == io_state_in_1 ? 8'h72 : _GEN_319; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_321 = 8'h41 == io_state_in_1 ? 8'hf8 : _GEN_320; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_322 = 8'h42 == io_state_in_1 ? 8'hf6 : _GEN_321; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_323 = 8'h43 == io_state_in_1 ? 8'h64 : _GEN_322; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_324 = 8'h44 == io_state_in_1 ? 8'h86 : _GEN_323; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_325 = 8'h45 == io_state_in_1 ? 8'h68 : _GEN_324; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_326 = 8'h46 == io_state_in_1 ? 8'h98 : _GEN_325; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_327 = 8'h47 == io_state_in_1 ? 8'h16 : _GEN_326; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_328 = 8'h48 == io_state_in_1 ? 8'hd4 : _GEN_327; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_329 = 8'h49 == io_state_in_1 ? 8'ha4 : _GEN_328; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_330 = 8'h4a == io_state_in_1 ? 8'h5c : _GEN_329; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_331 = 8'h4b == io_state_in_1 ? 8'hcc : _GEN_330; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_332 = 8'h4c == io_state_in_1 ? 8'h5d : _GEN_331; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_333 = 8'h4d == io_state_in_1 ? 8'h65 : _GEN_332; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_334 = 8'h4e == io_state_in_1 ? 8'hb6 : _GEN_333; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_335 = 8'h4f == io_state_in_1 ? 8'h92 : _GEN_334; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_336 = 8'h50 == io_state_in_1 ? 8'h6c : _GEN_335; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_337 = 8'h51 == io_state_in_1 ? 8'h70 : _GEN_336; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_338 = 8'h52 == io_state_in_1 ? 8'h48 : _GEN_337; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_339 = 8'h53 == io_state_in_1 ? 8'h50 : _GEN_338; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_340 = 8'h54 == io_state_in_1 ? 8'hfd : _GEN_339; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_341 = 8'h55 == io_state_in_1 ? 8'hed : _GEN_340; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_342 = 8'h56 == io_state_in_1 ? 8'hb9 : _GEN_341; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_343 = 8'h57 == io_state_in_1 ? 8'hda : _GEN_342; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_344 = 8'h58 == io_state_in_1 ? 8'h5e : _GEN_343; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_345 = 8'h59 == io_state_in_1 ? 8'h15 : _GEN_344; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_346 = 8'h5a == io_state_in_1 ? 8'h46 : _GEN_345; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_347 = 8'h5b == io_state_in_1 ? 8'h57 : _GEN_346; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_348 = 8'h5c == io_state_in_1 ? 8'ha7 : _GEN_347; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_349 = 8'h5d == io_state_in_1 ? 8'h8d : _GEN_348; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_350 = 8'h5e == io_state_in_1 ? 8'h9d : _GEN_349; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_351 = 8'h5f == io_state_in_1 ? 8'h84 : _GEN_350; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_352 = 8'h60 == io_state_in_1 ? 8'h90 : _GEN_351; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_353 = 8'h61 == io_state_in_1 ? 8'hd8 : _GEN_352; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_354 = 8'h62 == io_state_in_1 ? 8'hab : _GEN_353; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_355 = 8'h63 == io_state_in_1 ? 8'h0 : _GEN_354; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_356 = 8'h64 == io_state_in_1 ? 8'h8c : _GEN_355; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_357 = 8'h65 == io_state_in_1 ? 8'hbc : _GEN_356; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_358 = 8'h66 == io_state_in_1 ? 8'hd3 : _GEN_357; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_359 = 8'h67 == io_state_in_1 ? 8'ha : _GEN_358; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_360 = 8'h68 == io_state_in_1 ? 8'hf7 : _GEN_359; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_361 = 8'h69 == io_state_in_1 ? 8'he4 : _GEN_360; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_362 = 8'h6a == io_state_in_1 ? 8'h58 : _GEN_361; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_363 = 8'h6b == io_state_in_1 ? 8'h5 : _GEN_362; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_364 = 8'h6c == io_state_in_1 ? 8'hb8 : _GEN_363; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_365 = 8'h6d == io_state_in_1 ? 8'hb3 : _GEN_364; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_366 = 8'h6e == io_state_in_1 ? 8'h45 : _GEN_365; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_367 = 8'h6f == io_state_in_1 ? 8'h6 : _GEN_366; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_368 = 8'h70 == io_state_in_1 ? 8'hd0 : _GEN_367; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_369 = 8'h71 == io_state_in_1 ? 8'h2c : _GEN_368; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_370 = 8'h72 == io_state_in_1 ? 8'h1e : _GEN_369; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_371 = 8'h73 == io_state_in_1 ? 8'h8f : _GEN_370; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_372 = 8'h74 == io_state_in_1 ? 8'hca : _GEN_371; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_373 = 8'h75 == io_state_in_1 ? 8'h3f : _GEN_372; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_374 = 8'h76 == io_state_in_1 ? 8'hf : _GEN_373; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_375 = 8'h77 == io_state_in_1 ? 8'h2 : _GEN_374; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_376 = 8'h78 == io_state_in_1 ? 8'hc1 : _GEN_375; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_377 = 8'h79 == io_state_in_1 ? 8'haf : _GEN_376; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_378 = 8'h7a == io_state_in_1 ? 8'hbd : _GEN_377; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_379 = 8'h7b == io_state_in_1 ? 8'h3 : _GEN_378; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_380 = 8'h7c == io_state_in_1 ? 8'h1 : _GEN_379; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_381 = 8'h7d == io_state_in_1 ? 8'h13 : _GEN_380; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_382 = 8'h7e == io_state_in_1 ? 8'h8a : _GEN_381; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_383 = 8'h7f == io_state_in_1 ? 8'h6b : _GEN_382; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_384 = 8'h80 == io_state_in_1 ? 8'h3a : _GEN_383; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_385 = 8'h81 == io_state_in_1 ? 8'h91 : _GEN_384; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_386 = 8'h82 == io_state_in_1 ? 8'h11 : _GEN_385; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_387 = 8'h83 == io_state_in_1 ? 8'h41 : _GEN_386; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_388 = 8'h84 == io_state_in_1 ? 8'h4f : _GEN_387; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_389 = 8'h85 == io_state_in_1 ? 8'h67 : _GEN_388; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_390 = 8'h86 == io_state_in_1 ? 8'hdc : _GEN_389; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_391 = 8'h87 == io_state_in_1 ? 8'hea : _GEN_390; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_392 = 8'h88 == io_state_in_1 ? 8'h97 : _GEN_391; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_393 = 8'h89 == io_state_in_1 ? 8'hf2 : _GEN_392; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_394 = 8'h8a == io_state_in_1 ? 8'hcf : _GEN_393; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_395 = 8'h8b == io_state_in_1 ? 8'hce : _GEN_394; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_396 = 8'h8c == io_state_in_1 ? 8'hf0 : _GEN_395; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_397 = 8'h8d == io_state_in_1 ? 8'hb4 : _GEN_396; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_398 = 8'h8e == io_state_in_1 ? 8'he6 : _GEN_397; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_399 = 8'h8f == io_state_in_1 ? 8'h73 : _GEN_398; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_400 = 8'h90 == io_state_in_1 ? 8'h96 : _GEN_399; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_401 = 8'h91 == io_state_in_1 ? 8'hac : _GEN_400; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_402 = 8'h92 == io_state_in_1 ? 8'h74 : _GEN_401; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_403 = 8'h93 == io_state_in_1 ? 8'h22 : _GEN_402; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_404 = 8'h94 == io_state_in_1 ? 8'he7 : _GEN_403; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_405 = 8'h95 == io_state_in_1 ? 8'had : _GEN_404; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_406 = 8'h96 == io_state_in_1 ? 8'h35 : _GEN_405; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_407 = 8'h97 == io_state_in_1 ? 8'h85 : _GEN_406; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_408 = 8'h98 == io_state_in_1 ? 8'he2 : _GEN_407; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_409 = 8'h99 == io_state_in_1 ? 8'hf9 : _GEN_408; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_410 = 8'h9a == io_state_in_1 ? 8'h37 : _GEN_409; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_411 = 8'h9b == io_state_in_1 ? 8'he8 : _GEN_410; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_412 = 8'h9c == io_state_in_1 ? 8'h1c : _GEN_411; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_413 = 8'h9d == io_state_in_1 ? 8'h75 : _GEN_412; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_414 = 8'h9e == io_state_in_1 ? 8'hdf : _GEN_413; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_415 = 8'h9f == io_state_in_1 ? 8'h6e : _GEN_414; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_416 = 8'ha0 == io_state_in_1 ? 8'h47 : _GEN_415; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_417 = 8'ha1 == io_state_in_1 ? 8'hf1 : _GEN_416; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_418 = 8'ha2 == io_state_in_1 ? 8'h1a : _GEN_417; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_419 = 8'ha3 == io_state_in_1 ? 8'h71 : _GEN_418; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_420 = 8'ha4 == io_state_in_1 ? 8'h1d : _GEN_419; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_421 = 8'ha5 == io_state_in_1 ? 8'h29 : _GEN_420; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_422 = 8'ha6 == io_state_in_1 ? 8'hc5 : _GEN_421; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_423 = 8'ha7 == io_state_in_1 ? 8'h89 : _GEN_422; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_424 = 8'ha8 == io_state_in_1 ? 8'h6f : _GEN_423; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_425 = 8'ha9 == io_state_in_1 ? 8'hb7 : _GEN_424; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_426 = 8'haa == io_state_in_1 ? 8'h62 : _GEN_425; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_427 = 8'hab == io_state_in_1 ? 8'he : _GEN_426; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_428 = 8'hac == io_state_in_1 ? 8'haa : _GEN_427; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_429 = 8'had == io_state_in_1 ? 8'h18 : _GEN_428; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_430 = 8'hae == io_state_in_1 ? 8'hbe : _GEN_429; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_431 = 8'haf == io_state_in_1 ? 8'h1b : _GEN_430; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_432 = 8'hb0 == io_state_in_1 ? 8'hfc : _GEN_431; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_433 = 8'hb1 == io_state_in_1 ? 8'h56 : _GEN_432; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_434 = 8'hb2 == io_state_in_1 ? 8'h3e : _GEN_433; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_435 = 8'hb3 == io_state_in_1 ? 8'h4b : _GEN_434; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_436 = 8'hb4 == io_state_in_1 ? 8'hc6 : _GEN_435; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_437 = 8'hb5 == io_state_in_1 ? 8'hd2 : _GEN_436; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_438 = 8'hb6 == io_state_in_1 ? 8'h79 : _GEN_437; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_439 = 8'hb7 == io_state_in_1 ? 8'h20 : _GEN_438; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_440 = 8'hb8 == io_state_in_1 ? 8'h9a : _GEN_439; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_441 = 8'hb9 == io_state_in_1 ? 8'hdb : _GEN_440; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_442 = 8'hba == io_state_in_1 ? 8'hc0 : _GEN_441; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_443 = 8'hbb == io_state_in_1 ? 8'hfe : _GEN_442; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_444 = 8'hbc == io_state_in_1 ? 8'h78 : _GEN_443; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_445 = 8'hbd == io_state_in_1 ? 8'hcd : _GEN_444; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_446 = 8'hbe == io_state_in_1 ? 8'h5a : _GEN_445; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_447 = 8'hbf == io_state_in_1 ? 8'hf4 : _GEN_446; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_448 = 8'hc0 == io_state_in_1 ? 8'h1f : _GEN_447; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_449 = 8'hc1 == io_state_in_1 ? 8'hdd : _GEN_448; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_450 = 8'hc2 == io_state_in_1 ? 8'ha8 : _GEN_449; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_451 = 8'hc3 == io_state_in_1 ? 8'h33 : _GEN_450; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_452 = 8'hc4 == io_state_in_1 ? 8'h88 : _GEN_451; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_453 = 8'hc5 == io_state_in_1 ? 8'h7 : _GEN_452; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_454 = 8'hc6 == io_state_in_1 ? 8'hc7 : _GEN_453; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_455 = 8'hc7 == io_state_in_1 ? 8'h31 : _GEN_454; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_456 = 8'hc8 == io_state_in_1 ? 8'hb1 : _GEN_455; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_457 = 8'hc9 == io_state_in_1 ? 8'h12 : _GEN_456; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_458 = 8'hca == io_state_in_1 ? 8'h10 : _GEN_457; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_459 = 8'hcb == io_state_in_1 ? 8'h59 : _GEN_458; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_460 = 8'hcc == io_state_in_1 ? 8'h27 : _GEN_459; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_461 = 8'hcd == io_state_in_1 ? 8'h80 : _GEN_460; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_462 = 8'hce == io_state_in_1 ? 8'hec : _GEN_461; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_463 = 8'hcf == io_state_in_1 ? 8'h5f : _GEN_462; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_464 = 8'hd0 == io_state_in_1 ? 8'h60 : _GEN_463; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_465 = 8'hd1 == io_state_in_1 ? 8'h51 : _GEN_464; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_466 = 8'hd2 == io_state_in_1 ? 8'h7f : _GEN_465; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_467 = 8'hd3 == io_state_in_1 ? 8'ha9 : _GEN_466; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_468 = 8'hd4 == io_state_in_1 ? 8'h19 : _GEN_467; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_469 = 8'hd5 == io_state_in_1 ? 8'hb5 : _GEN_468; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_470 = 8'hd6 == io_state_in_1 ? 8'h4a : _GEN_469; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_471 = 8'hd7 == io_state_in_1 ? 8'hd : _GEN_470; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_472 = 8'hd8 == io_state_in_1 ? 8'h2d : _GEN_471; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_473 = 8'hd9 == io_state_in_1 ? 8'he5 : _GEN_472; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_474 = 8'hda == io_state_in_1 ? 8'h7a : _GEN_473; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_475 = 8'hdb == io_state_in_1 ? 8'h9f : _GEN_474; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_476 = 8'hdc == io_state_in_1 ? 8'h93 : _GEN_475; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_477 = 8'hdd == io_state_in_1 ? 8'hc9 : _GEN_476; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_478 = 8'hde == io_state_in_1 ? 8'h9c : _GEN_477; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_479 = 8'hdf == io_state_in_1 ? 8'hef : _GEN_478; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_480 = 8'he0 == io_state_in_1 ? 8'ha0 : _GEN_479; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_481 = 8'he1 == io_state_in_1 ? 8'he0 : _GEN_480; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_482 = 8'he2 == io_state_in_1 ? 8'h3b : _GEN_481; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_483 = 8'he3 == io_state_in_1 ? 8'h4d : _GEN_482; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_484 = 8'he4 == io_state_in_1 ? 8'hae : _GEN_483; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_485 = 8'he5 == io_state_in_1 ? 8'h2a : _GEN_484; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_486 = 8'he6 == io_state_in_1 ? 8'hf5 : _GEN_485; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_487 = 8'he7 == io_state_in_1 ? 8'hb0 : _GEN_486; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_488 = 8'he8 == io_state_in_1 ? 8'hc8 : _GEN_487; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_489 = 8'he9 == io_state_in_1 ? 8'heb : _GEN_488; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_490 = 8'hea == io_state_in_1 ? 8'hbb : _GEN_489; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_491 = 8'heb == io_state_in_1 ? 8'h3c : _GEN_490; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_492 = 8'hec == io_state_in_1 ? 8'h83 : _GEN_491; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_493 = 8'hed == io_state_in_1 ? 8'h53 : _GEN_492; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_494 = 8'hee == io_state_in_1 ? 8'h99 : _GEN_493; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_495 = 8'hef == io_state_in_1 ? 8'h61 : _GEN_494; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_496 = 8'hf0 == io_state_in_1 ? 8'h17 : _GEN_495; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_497 = 8'hf1 == io_state_in_1 ? 8'h2b : _GEN_496; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_498 = 8'hf2 == io_state_in_1 ? 8'h4 : _GEN_497; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_499 = 8'hf3 == io_state_in_1 ? 8'h7e : _GEN_498; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_500 = 8'hf4 == io_state_in_1 ? 8'hba : _GEN_499; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_501 = 8'hf5 == io_state_in_1 ? 8'h77 : _GEN_500; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_502 = 8'hf6 == io_state_in_1 ? 8'hd6 : _GEN_501; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_503 = 8'hf7 == io_state_in_1 ? 8'h26 : _GEN_502; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_504 = 8'hf8 == io_state_in_1 ? 8'he1 : _GEN_503; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_505 = 8'hf9 == io_state_in_1 ? 8'h69 : _GEN_504; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_506 = 8'hfa == io_state_in_1 ? 8'h14 : _GEN_505; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_507 = 8'hfb == io_state_in_1 ? 8'h63 : _GEN_506; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_508 = 8'hfc == io_state_in_1 ? 8'h55 : _GEN_507; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_509 = 8'hfd == io_state_in_1 ? 8'h21 : _GEN_508; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_510 = 8'hfe == io_state_in_1 ? 8'hc : _GEN_509; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_513 = 8'h1 == io_state_in_2 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_514 = 8'h2 == io_state_in_2 ? 8'h6a : _GEN_513; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_515 = 8'h3 == io_state_in_2 ? 8'hd5 : _GEN_514; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_516 = 8'h4 == io_state_in_2 ? 8'h30 : _GEN_515; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_517 = 8'h5 == io_state_in_2 ? 8'h36 : _GEN_516; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_518 = 8'h6 == io_state_in_2 ? 8'ha5 : _GEN_517; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_519 = 8'h7 == io_state_in_2 ? 8'h38 : _GEN_518; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_520 = 8'h8 == io_state_in_2 ? 8'hbf : _GEN_519; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_521 = 8'h9 == io_state_in_2 ? 8'h40 : _GEN_520; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_522 = 8'ha == io_state_in_2 ? 8'ha3 : _GEN_521; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_523 = 8'hb == io_state_in_2 ? 8'h9e : _GEN_522; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_524 = 8'hc == io_state_in_2 ? 8'h81 : _GEN_523; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_525 = 8'hd == io_state_in_2 ? 8'hf3 : _GEN_524; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_526 = 8'he == io_state_in_2 ? 8'hd7 : _GEN_525; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_527 = 8'hf == io_state_in_2 ? 8'hfb : _GEN_526; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_528 = 8'h10 == io_state_in_2 ? 8'h7c : _GEN_527; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_529 = 8'h11 == io_state_in_2 ? 8'he3 : _GEN_528; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_530 = 8'h12 == io_state_in_2 ? 8'h39 : _GEN_529; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_531 = 8'h13 == io_state_in_2 ? 8'h82 : _GEN_530; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_532 = 8'h14 == io_state_in_2 ? 8'h9b : _GEN_531; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_533 = 8'h15 == io_state_in_2 ? 8'h2f : _GEN_532; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_534 = 8'h16 == io_state_in_2 ? 8'hff : _GEN_533; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_535 = 8'h17 == io_state_in_2 ? 8'h87 : _GEN_534; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_536 = 8'h18 == io_state_in_2 ? 8'h34 : _GEN_535; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_537 = 8'h19 == io_state_in_2 ? 8'h8e : _GEN_536; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_538 = 8'h1a == io_state_in_2 ? 8'h43 : _GEN_537; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_539 = 8'h1b == io_state_in_2 ? 8'h44 : _GEN_538; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_540 = 8'h1c == io_state_in_2 ? 8'hc4 : _GEN_539; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_541 = 8'h1d == io_state_in_2 ? 8'hde : _GEN_540; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_542 = 8'h1e == io_state_in_2 ? 8'he9 : _GEN_541; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_543 = 8'h1f == io_state_in_2 ? 8'hcb : _GEN_542; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_544 = 8'h20 == io_state_in_2 ? 8'h54 : _GEN_543; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_545 = 8'h21 == io_state_in_2 ? 8'h7b : _GEN_544; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_546 = 8'h22 == io_state_in_2 ? 8'h94 : _GEN_545; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_547 = 8'h23 == io_state_in_2 ? 8'h32 : _GEN_546; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_548 = 8'h24 == io_state_in_2 ? 8'ha6 : _GEN_547; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_549 = 8'h25 == io_state_in_2 ? 8'hc2 : _GEN_548; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_550 = 8'h26 == io_state_in_2 ? 8'h23 : _GEN_549; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_551 = 8'h27 == io_state_in_2 ? 8'h3d : _GEN_550; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_552 = 8'h28 == io_state_in_2 ? 8'hee : _GEN_551; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_553 = 8'h29 == io_state_in_2 ? 8'h4c : _GEN_552; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_554 = 8'h2a == io_state_in_2 ? 8'h95 : _GEN_553; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_555 = 8'h2b == io_state_in_2 ? 8'hb : _GEN_554; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_556 = 8'h2c == io_state_in_2 ? 8'h42 : _GEN_555; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_557 = 8'h2d == io_state_in_2 ? 8'hfa : _GEN_556; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_558 = 8'h2e == io_state_in_2 ? 8'hc3 : _GEN_557; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_559 = 8'h2f == io_state_in_2 ? 8'h4e : _GEN_558; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_560 = 8'h30 == io_state_in_2 ? 8'h8 : _GEN_559; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_561 = 8'h31 == io_state_in_2 ? 8'h2e : _GEN_560; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_562 = 8'h32 == io_state_in_2 ? 8'ha1 : _GEN_561; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_563 = 8'h33 == io_state_in_2 ? 8'h66 : _GEN_562; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_564 = 8'h34 == io_state_in_2 ? 8'h28 : _GEN_563; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_565 = 8'h35 == io_state_in_2 ? 8'hd9 : _GEN_564; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_566 = 8'h36 == io_state_in_2 ? 8'h24 : _GEN_565; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_567 = 8'h37 == io_state_in_2 ? 8'hb2 : _GEN_566; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_568 = 8'h38 == io_state_in_2 ? 8'h76 : _GEN_567; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_569 = 8'h39 == io_state_in_2 ? 8'h5b : _GEN_568; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_570 = 8'h3a == io_state_in_2 ? 8'ha2 : _GEN_569; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_571 = 8'h3b == io_state_in_2 ? 8'h49 : _GEN_570; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_572 = 8'h3c == io_state_in_2 ? 8'h6d : _GEN_571; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_573 = 8'h3d == io_state_in_2 ? 8'h8b : _GEN_572; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_574 = 8'h3e == io_state_in_2 ? 8'hd1 : _GEN_573; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_575 = 8'h3f == io_state_in_2 ? 8'h25 : _GEN_574; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_576 = 8'h40 == io_state_in_2 ? 8'h72 : _GEN_575; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_577 = 8'h41 == io_state_in_2 ? 8'hf8 : _GEN_576; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_578 = 8'h42 == io_state_in_2 ? 8'hf6 : _GEN_577; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_579 = 8'h43 == io_state_in_2 ? 8'h64 : _GEN_578; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_580 = 8'h44 == io_state_in_2 ? 8'h86 : _GEN_579; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_581 = 8'h45 == io_state_in_2 ? 8'h68 : _GEN_580; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_582 = 8'h46 == io_state_in_2 ? 8'h98 : _GEN_581; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_583 = 8'h47 == io_state_in_2 ? 8'h16 : _GEN_582; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_584 = 8'h48 == io_state_in_2 ? 8'hd4 : _GEN_583; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_585 = 8'h49 == io_state_in_2 ? 8'ha4 : _GEN_584; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_586 = 8'h4a == io_state_in_2 ? 8'h5c : _GEN_585; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_587 = 8'h4b == io_state_in_2 ? 8'hcc : _GEN_586; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_588 = 8'h4c == io_state_in_2 ? 8'h5d : _GEN_587; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_589 = 8'h4d == io_state_in_2 ? 8'h65 : _GEN_588; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_590 = 8'h4e == io_state_in_2 ? 8'hb6 : _GEN_589; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_591 = 8'h4f == io_state_in_2 ? 8'h92 : _GEN_590; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_592 = 8'h50 == io_state_in_2 ? 8'h6c : _GEN_591; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_593 = 8'h51 == io_state_in_2 ? 8'h70 : _GEN_592; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_594 = 8'h52 == io_state_in_2 ? 8'h48 : _GEN_593; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_595 = 8'h53 == io_state_in_2 ? 8'h50 : _GEN_594; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_596 = 8'h54 == io_state_in_2 ? 8'hfd : _GEN_595; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_597 = 8'h55 == io_state_in_2 ? 8'hed : _GEN_596; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_598 = 8'h56 == io_state_in_2 ? 8'hb9 : _GEN_597; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_599 = 8'h57 == io_state_in_2 ? 8'hda : _GEN_598; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_600 = 8'h58 == io_state_in_2 ? 8'h5e : _GEN_599; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_601 = 8'h59 == io_state_in_2 ? 8'h15 : _GEN_600; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_602 = 8'h5a == io_state_in_2 ? 8'h46 : _GEN_601; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_603 = 8'h5b == io_state_in_2 ? 8'h57 : _GEN_602; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_604 = 8'h5c == io_state_in_2 ? 8'ha7 : _GEN_603; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_605 = 8'h5d == io_state_in_2 ? 8'h8d : _GEN_604; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_606 = 8'h5e == io_state_in_2 ? 8'h9d : _GEN_605; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_607 = 8'h5f == io_state_in_2 ? 8'h84 : _GEN_606; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_608 = 8'h60 == io_state_in_2 ? 8'h90 : _GEN_607; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_609 = 8'h61 == io_state_in_2 ? 8'hd8 : _GEN_608; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_610 = 8'h62 == io_state_in_2 ? 8'hab : _GEN_609; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_611 = 8'h63 == io_state_in_2 ? 8'h0 : _GEN_610; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_612 = 8'h64 == io_state_in_2 ? 8'h8c : _GEN_611; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_613 = 8'h65 == io_state_in_2 ? 8'hbc : _GEN_612; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_614 = 8'h66 == io_state_in_2 ? 8'hd3 : _GEN_613; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_615 = 8'h67 == io_state_in_2 ? 8'ha : _GEN_614; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_616 = 8'h68 == io_state_in_2 ? 8'hf7 : _GEN_615; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_617 = 8'h69 == io_state_in_2 ? 8'he4 : _GEN_616; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_618 = 8'h6a == io_state_in_2 ? 8'h58 : _GEN_617; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_619 = 8'h6b == io_state_in_2 ? 8'h5 : _GEN_618; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_620 = 8'h6c == io_state_in_2 ? 8'hb8 : _GEN_619; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_621 = 8'h6d == io_state_in_2 ? 8'hb3 : _GEN_620; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_622 = 8'h6e == io_state_in_2 ? 8'h45 : _GEN_621; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_623 = 8'h6f == io_state_in_2 ? 8'h6 : _GEN_622; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_624 = 8'h70 == io_state_in_2 ? 8'hd0 : _GEN_623; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_625 = 8'h71 == io_state_in_2 ? 8'h2c : _GEN_624; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_626 = 8'h72 == io_state_in_2 ? 8'h1e : _GEN_625; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_627 = 8'h73 == io_state_in_2 ? 8'h8f : _GEN_626; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_628 = 8'h74 == io_state_in_2 ? 8'hca : _GEN_627; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_629 = 8'h75 == io_state_in_2 ? 8'h3f : _GEN_628; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_630 = 8'h76 == io_state_in_2 ? 8'hf : _GEN_629; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_631 = 8'h77 == io_state_in_2 ? 8'h2 : _GEN_630; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_632 = 8'h78 == io_state_in_2 ? 8'hc1 : _GEN_631; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_633 = 8'h79 == io_state_in_2 ? 8'haf : _GEN_632; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_634 = 8'h7a == io_state_in_2 ? 8'hbd : _GEN_633; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_635 = 8'h7b == io_state_in_2 ? 8'h3 : _GEN_634; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_636 = 8'h7c == io_state_in_2 ? 8'h1 : _GEN_635; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_637 = 8'h7d == io_state_in_2 ? 8'h13 : _GEN_636; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_638 = 8'h7e == io_state_in_2 ? 8'h8a : _GEN_637; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_639 = 8'h7f == io_state_in_2 ? 8'h6b : _GEN_638; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_640 = 8'h80 == io_state_in_2 ? 8'h3a : _GEN_639; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_641 = 8'h81 == io_state_in_2 ? 8'h91 : _GEN_640; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_642 = 8'h82 == io_state_in_2 ? 8'h11 : _GEN_641; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_643 = 8'h83 == io_state_in_2 ? 8'h41 : _GEN_642; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_644 = 8'h84 == io_state_in_2 ? 8'h4f : _GEN_643; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_645 = 8'h85 == io_state_in_2 ? 8'h67 : _GEN_644; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_646 = 8'h86 == io_state_in_2 ? 8'hdc : _GEN_645; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_647 = 8'h87 == io_state_in_2 ? 8'hea : _GEN_646; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_648 = 8'h88 == io_state_in_2 ? 8'h97 : _GEN_647; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_649 = 8'h89 == io_state_in_2 ? 8'hf2 : _GEN_648; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_650 = 8'h8a == io_state_in_2 ? 8'hcf : _GEN_649; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_651 = 8'h8b == io_state_in_2 ? 8'hce : _GEN_650; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_652 = 8'h8c == io_state_in_2 ? 8'hf0 : _GEN_651; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_653 = 8'h8d == io_state_in_2 ? 8'hb4 : _GEN_652; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_654 = 8'h8e == io_state_in_2 ? 8'he6 : _GEN_653; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_655 = 8'h8f == io_state_in_2 ? 8'h73 : _GEN_654; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_656 = 8'h90 == io_state_in_2 ? 8'h96 : _GEN_655; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_657 = 8'h91 == io_state_in_2 ? 8'hac : _GEN_656; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_658 = 8'h92 == io_state_in_2 ? 8'h74 : _GEN_657; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_659 = 8'h93 == io_state_in_2 ? 8'h22 : _GEN_658; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_660 = 8'h94 == io_state_in_2 ? 8'he7 : _GEN_659; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_661 = 8'h95 == io_state_in_2 ? 8'had : _GEN_660; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_662 = 8'h96 == io_state_in_2 ? 8'h35 : _GEN_661; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_663 = 8'h97 == io_state_in_2 ? 8'h85 : _GEN_662; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_664 = 8'h98 == io_state_in_2 ? 8'he2 : _GEN_663; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_665 = 8'h99 == io_state_in_2 ? 8'hf9 : _GEN_664; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_666 = 8'h9a == io_state_in_2 ? 8'h37 : _GEN_665; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_667 = 8'h9b == io_state_in_2 ? 8'he8 : _GEN_666; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_668 = 8'h9c == io_state_in_2 ? 8'h1c : _GEN_667; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_669 = 8'h9d == io_state_in_2 ? 8'h75 : _GEN_668; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_670 = 8'h9e == io_state_in_2 ? 8'hdf : _GEN_669; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_671 = 8'h9f == io_state_in_2 ? 8'h6e : _GEN_670; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_672 = 8'ha0 == io_state_in_2 ? 8'h47 : _GEN_671; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_673 = 8'ha1 == io_state_in_2 ? 8'hf1 : _GEN_672; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_674 = 8'ha2 == io_state_in_2 ? 8'h1a : _GEN_673; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_675 = 8'ha3 == io_state_in_2 ? 8'h71 : _GEN_674; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_676 = 8'ha4 == io_state_in_2 ? 8'h1d : _GEN_675; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_677 = 8'ha5 == io_state_in_2 ? 8'h29 : _GEN_676; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_678 = 8'ha6 == io_state_in_2 ? 8'hc5 : _GEN_677; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_679 = 8'ha7 == io_state_in_2 ? 8'h89 : _GEN_678; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_680 = 8'ha8 == io_state_in_2 ? 8'h6f : _GEN_679; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_681 = 8'ha9 == io_state_in_2 ? 8'hb7 : _GEN_680; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_682 = 8'haa == io_state_in_2 ? 8'h62 : _GEN_681; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_683 = 8'hab == io_state_in_2 ? 8'he : _GEN_682; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_684 = 8'hac == io_state_in_2 ? 8'haa : _GEN_683; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_685 = 8'had == io_state_in_2 ? 8'h18 : _GEN_684; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_686 = 8'hae == io_state_in_2 ? 8'hbe : _GEN_685; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_687 = 8'haf == io_state_in_2 ? 8'h1b : _GEN_686; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_688 = 8'hb0 == io_state_in_2 ? 8'hfc : _GEN_687; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_689 = 8'hb1 == io_state_in_2 ? 8'h56 : _GEN_688; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_690 = 8'hb2 == io_state_in_2 ? 8'h3e : _GEN_689; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_691 = 8'hb3 == io_state_in_2 ? 8'h4b : _GEN_690; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_692 = 8'hb4 == io_state_in_2 ? 8'hc6 : _GEN_691; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_693 = 8'hb5 == io_state_in_2 ? 8'hd2 : _GEN_692; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_694 = 8'hb6 == io_state_in_2 ? 8'h79 : _GEN_693; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_695 = 8'hb7 == io_state_in_2 ? 8'h20 : _GEN_694; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_696 = 8'hb8 == io_state_in_2 ? 8'h9a : _GEN_695; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_697 = 8'hb9 == io_state_in_2 ? 8'hdb : _GEN_696; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_698 = 8'hba == io_state_in_2 ? 8'hc0 : _GEN_697; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_699 = 8'hbb == io_state_in_2 ? 8'hfe : _GEN_698; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_700 = 8'hbc == io_state_in_2 ? 8'h78 : _GEN_699; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_701 = 8'hbd == io_state_in_2 ? 8'hcd : _GEN_700; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_702 = 8'hbe == io_state_in_2 ? 8'h5a : _GEN_701; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_703 = 8'hbf == io_state_in_2 ? 8'hf4 : _GEN_702; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_704 = 8'hc0 == io_state_in_2 ? 8'h1f : _GEN_703; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_705 = 8'hc1 == io_state_in_2 ? 8'hdd : _GEN_704; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_706 = 8'hc2 == io_state_in_2 ? 8'ha8 : _GEN_705; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_707 = 8'hc3 == io_state_in_2 ? 8'h33 : _GEN_706; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_708 = 8'hc4 == io_state_in_2 ? 8'h88 : _GEN_707; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_709 = 8'hc5 == io_state_in_2 ? 8'h7 : _GEN_708; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_710 = 8'hc6 == io_state_in_2 ? 8'hc7 : _GEN_709; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_711 = 8'hc7 == io_state_in_2 ? 8'h31 : _GEN_710; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_712 = 8'hc8 == io_state_in_2 ? 8'hb1 : _GEN_711; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_713 = 8'hc9 == io_state_in_2 ? 8'h12 : _GEN_712; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_714 = 8'hca == io_state_in_2 ? 8'h10 : _GEN_713; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_715 = 8'hcb == io_state_in_2 ? 8'h59 : _GEN_714; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_716 = 8'hcc == io_state_in_2 ? 8'h27 : _GEN_715; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_717 = 8'hcd == io_state_in_2 ? 8'h80 : _GEN_716; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_718 = 8'hce == io_state_in_2 ? 8'hec : _GEN_717; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_719 = 8'hcf == io_state_in_2 ? 8'h5f : _GEN_718; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_720 = 8'hd0 == io_state_in_2 ? 8'h60 : _GEN_719; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_721 = 8'hd1 == io_state_in_2 ? 8'h51 : _GEN_720; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_722 = 8'hd2 == io_state_in_2 ? 8'h7f : _GEN_721; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_723 = 8'hd3 == io_state_in_2 ? 8'ha9 : _GEN_722; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_724 = 8'hd4 == io_state_in_2 ? 8'h19 : _GEN_723; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_725 = 8'hd5 == io_state_in_2 ? 8'hb5 : _GEN_724; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_726 = 8'hd6 == io_state_in_2 ? 8'h4a : _GEN_725; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_727 = 8'hd7 == io_state_in_2 ? 8'hd : _GEN_726; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_728 = 8'hd8 == io_state_in_2 ? 8'h2d : _GEN_727; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_729 = 8'hd9 == io_state_in_2 ? 8'he5 : _GEN_728; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_730 = 8'hda == io_state_in_2 ? 8'h7a : _GEN_729; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_731 = 8'hdb == io_state_in_2 ? 8'h9f : _GEN_730; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_732 = 8'hdc == io_state_in_2 ? 8'h93 : _GEN_731; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_733 = 8'hdd == io_state_in_2 ? 8'hc9 : _GEN_732; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_734 = 8'hde == io_state_in_2 ? 8'h9c : _GEN_733; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_735 = 8'hdf == io_state_in_2 ? 8'hef : _GEN_734; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_736 = 8'he0 == io_state_in_2 ? 8'ha0 : _GEN_735; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_737 = 8'he1 == io_state_in_2 ? 8'he0 : _GEN_736; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_738 = 8'he2 == io_state_in_2 ? 8'h3b : _GEN_737; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_739 = 8'he3 == io_state_in_2 ? 8'h4d : _GEN_738; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_740 = 8'he4 == io_state_in_2 ? 8'hae : _GEN_739; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_741 = 8'he5 == io_state_in_2 ? 8'h2a : _GEN_740; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_742 = 8'he6 == io_state_in_2 ? 8'hf5 : _GEN_741; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_743 = 8'he7 == io_state_in_2 ? 8'hb0 : _GEN_742; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_744 = 8'he8 == io_state_in_2 ? 8'hc8 : _GEN_743; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_745 = 8'he9 == io_state_in_2 ? 8'heb : _GEN_744; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_746 = 8'hea == io_state_in_2 ? 8'hbb : _GEN_745; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_747 = 8'heb == io_state_in_2 ? 8'h3c : _GEN_746; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_748 = 8'hec == io_state_in_2 ? 8'h83 : _GEN_747; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_749 = 8'hed == io_state_in_2 ? 8'h53 : _GEN_748; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_750 = 8'hee == io_state_in_2 ? 8'h99 : _GEN_749; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_751 = 8'hef == io_state_in_2 ? 8'h61 : _GEN_750; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_752 = 8'hf0 == io_state_in_2 ? 8'h17 : _GEN_751; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_753 = 8'hf1 == io_state_in_2 ? 8'h2b : _GEN_752; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_754 = 8'hf2 == io_state_in_2 ? 8'h4 : _GEN_753; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_755 = 8'hf3 == io_state_in_2 ? 8'h7e : _GEN_754; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_756 = 8'hf4 == io_state_in_2 ? 8'hba : _GEN_755; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_757 = 8'hf5 == io_state_in_2 ? 8'h77 : _GEN_756; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_758 = 8'hf6 == io_state_in_2 ? 8'hd6 : _GEN_757; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_759 = 8'hf7 == io_state_in_2 ? 8'h26 : _GEN_758; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_760 = 8'hf8 == io_state_in_2 ? 8'he1 : _GEN_759; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_761 = 8'hf9 == io_state_in_2 ? 8'h69 : _GEN_760; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_762 = 8'hfa == io_state_in_2 ? 8'h14 : _GEN_761; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_763 = 8'hfb == io_state_in_2 ? 8'h63 : _GEN_762; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_764 = 8'hfc == io_state_in_2 ? 8'h55 : _GEN_763; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_765 = 8'hfd == io_state_in_2 ? 8'h21 : _GEN_764; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_766 = 8'hfe == io_state_in_2 ? 8'hc : _GEN_765; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_769 = 8'h1 == io_state_in_3 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_770 = 8'h2 == io_state_in_3 ? 8'h6a : _GEN_769; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_771 = 8'h3 == io_state_in_3 ? 8'hd5 : _GEN_770; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_772 = 8'h4 == io_state_in_3 ? 8'h30 : _GEN_771; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_773 = 8'h5 == io_state_in_3 ? 8'h36 : _GEN_772; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_774 = 8'h6 == io_state_in_3 ? 8'ha5 : _GEN_773; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_775 = 8'h7 == io_state_in_3 ? 8'h38 : _GEN_774; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_776 = 8'h8 == io_state_in_3 ? 8'hbf : _GEN_775; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_777 = 8'h9 == io_state_in_3 ? 8'h40 : _GEN_776; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_778 = 8'ha == io_state_in_3 ? 8'ha3 : _GEN_777; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_779 = 8'hb == io_state_in_3 ? 8'h9e : _GEN_778; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_780 = 8'hc == io_state_in_3 ? 8'h81 : _GEN_779; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_781 = 8'hd == io_state_in_3 ? 8'hf3 : _GEN_780; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_782 = 8'he == io_state_in_3 ? 8'hd7 : _GEN_781; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_783 = 8'hf == io_state_in_3 ? 8'hfb : _GEN_782; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_784 = 8'h10 == io_state_in_3 ? 8'h7c : _GEN_783; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_785 = 8'h11 == io_state_in_3 ? 8'he3 : _GEN_784; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_786 = 8'h12 == io_state_in_3 ? 8'h39 : _GEN_785; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_787 = 8'h13 == io_state_in_3 ? 8'h82 : _GEN_786; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_788 = 8'h14 == io_state_in_3 ? 8'h9b : _GEN_787; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_789 = 8'h15 == io_state_in_3 ? 8'h2f : _GEN_788; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_790 = 8'h16 == io_state_in_3 ? 8'hff : _GEN_789; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_791 = 8'h17 == io_state_in_3 ? 8'h87 : _GEN_790; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_792 = 8'h18 == io_state_in_3 ? 8'h34 : _GEN_791; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_793 = 8'h19 == io_state_in_3 ? 8'h8e : _GEN_792; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_794 = 8'h1a == io_state_in_3 ? 8'h43 : _GEN_793; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_795 = 8'h1b == io_state_in_3 ? 8'h44 : _GEN_794; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_796 = 8'h1c == io_state_in_3 ? 8'hc4 : _GEN_795; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_797 = 8'h1d == io_state_in_3 ? 8'hde : _GEN_796; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_798 = 8'h1e == io_state_in_3 ? 8'he9 : _GEN_797; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_799 = 8'h1f == io_state_in_3 ? 8'hcb : _GEN_798; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_800 = 8'h20 == io_state_in_3 ? 8'h54 : _GEN_799; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_801 = 8'h21 == io_state_in_3 ? 8'h7b : _GEN_800; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_802 = 8'h22 == io_state_in_3 ? 8'h94 : _GEN_801; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_803 = 8'h23 == io_state_in_3 ? 8'h32 : _GEN_802; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_804 = 8'h24 == io_state_in_3 ? 8'ha6 : _GEN_803; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_805 = 8'h25 == io_state_in_3 ? 8'hc2 : _GEN_804; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_806 = 8'h26 == io_state_in_3 ? 8'h23 : _GEN_805; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_807 = 8'h27 == io_state_in_3 ? 8'h3d : _GEN_806; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_808 = 8'h28 == io_state_in_3 ? 8'hee : _GEN_807; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_809 = 8'h29 == io_state_in_3 ? 8'h4c : _GEN_808; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_810 = 8'h2a == io_state_in_3 ? 8'h95 : _GEN_809; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_811 = 8'h2b == io_state_in_3 ? 8'hb : _GEN_810; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_812 = 8'h2c == io_state_in_3 ? 8'h42 : _GEN_811; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_813 = 8'h2d == io_state_in_3 ? 8'hfa : _GEN_812; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_814 = 8'h2e == io_state_in_3 ? 8'hc3 : _GEN_813; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_815 = 8'h2f == io_state_in_3 ? 8'h4e : _GEN_814; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_816 = 8'h30 == io_state_in_3 ? 8'h8 : _GEN_815; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_817 = 8'h31 == io_state_in_3 ? 8'h2e : _GEN_816; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_818 = 8'h32 == io_state_in_3 ? 8'ha1 : _GEN_817; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_819 = 8'h33 == io_state_in_3 ? 8'h66 : _GEN_818; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_820 = 8'h34 == io_state_in_3 ? 8'h28 : _GEN_819; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_821 = 8'h35 == io_state_in_3 ? 8'hd9 : _GEN_820; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_822 = 8'h36 == io_state_in_3 ? 8'h24 : _GEN_821; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_823 = 8'h37 == io_state_in_3 ? 8'hb2 : _GEN_822; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_824 = 8'h38 == io_state_in_3 ? 8'h76 : _GEN_823; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_825 = 8'h39 == io_state_in_3 ? 8'h5b : _GEN_824; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_826 = 8'h3a == io_state_in_3 ? 8'ha2 : _GEN_825; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_827 = 8'h3b == io_state_in_3 ? 8'h49 : _GEN_826; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_828 = 8'h3c == io_state_in_3 ? 8'h6d : _GEN_827; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_829 = 8'h3d == io_state_in_3 ? 8'h8b : _GEN_828; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_830 = 8'h3e == io_state_in_3 ? 8'hd1 : _GEN_829; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_831 = 8'h3f == io_state_in_3 ? 8'h25 : _GEN_830; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_832 = 8'h40 == io_state_in_3 ? 8'h72 : _GEN_831; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_833 = 8'h41 == io_state_in_3 ? 8'hf8 : _GEN_832; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_834 = 8'h42 == io_state_in_3 ? 8'hf6 : _GEN_833; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_835 = 8'h43 == io_state_in_3 ? 8'h64 : _GEN_834; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_836 = 8'h44 == io_state_in_3 ? 8'h86 : _GEN_835; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_837 = 8'h45 == io_state_in_3 ? 8'h68 : _GEN_836; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_838 = 8'h46 == io_state_in_3 ? 8'h98 : _GEN_837; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_839 = 8'h47 == io_state_in_3 ? 8'h16 : _GEN_838; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_840 = 8'h48 == io_state_in_3 ? 8'hd4 : _GEN_839; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_841 = 8'h49 == io_state_in_3 ? 8'ha4 : _GEN_840; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_842 = 8'h4a == io_state_in_3 ? 8'h5c : _GEN_841; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_843 = 8'h4b == io_state_in_3 ? 8'hcc : _GEN_842; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_844 = 8'h4c == io_state_in_3 ? 8'h5d : _GEN_843; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_845 = 8'h4d == io_state_in_3 ? 8'h65 : _GEN_844; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_846 = 8'h4e == io_state_in_3 ? 8'hb6 : _GEN_845; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_847 = 8'h4f == io_state_in_3 ? 8'h92 : _GEN_846; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_848 = 8'h50 == io_state_in_3 ? 8'h6c : _GEN_847; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_849 = 8'h51 == io_state_in_3 ? 8'h70 : _GEN_848; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_850 = 8'h52 == io_state_in_3 ? 8'h48 : _GEN_849; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_851 = 8'h53 == io_state_in_3 ? 8'h50 : _GEN_850; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_852 = 8'h54 == io_state_in_3 ? 8'hfd : _GEN_851; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_853 = 8'h55 == io_state_in_3 ? 8'hed : _GEN_852; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_854 = 8'h56 == io_state_in_3 ? 8'hb9 : _GEN_853; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_855 = 8'h57 == io_state_in_3 ? 8'hda : _GEN_854; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_856 = 8'h58 == io_state_in_3 ? 8'h5e : _GEN_855; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_857 = 8'h59 == io_state_in_3 ? 8'h15 : _GEN_856; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_858 = 8'h5a == io_state_in_3 ? 8'h46 : _GEN_857; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_859 = 8'h5b == io_state_in_3 ? 8'h57 : _GEN_858; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_860 = 8'h5c == io_state_in_3 ? 8'ha7 : _GEN_859; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_861 = 8'h5d == io_state_in_3 ? 8'h8d : _GEN_860; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_862 = 8'h5e == io_state_in_3 ? 8'h9d : _GEN_861; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_863 = 8'h5f == io_state_in_3 ? 8'h84 : _GEN_862; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_864 = 8'h60 == io_state_in_3 ? 8'h90 : _GEN_863; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_865 = 8'h61 == io_state_in_3 ? 8'hd8 : _GEN_864; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_866 = 8'h62 == io_state_in_3 ? 8'hab : _GEN_865; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_867 = 8'h63 == io_state_in_3 ? 8'h0 : _GEN_866; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_868 = 8'h64 == io_state_in_3 ? 8'h8c : _GEN_867; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_869 = 8'h65 == io_state_in_3 ? 8'hbc : _GEN_868; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_870 = 8'h66 == io_state_in_3 ? 8'hd3 : _GEN_869; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_871 = 8'h67 == io_state_in_3 ? 8'ha : _GEN_870; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_872 = 8'h68 == io_state_in_3 ? 8'hf7 : _GEN_871; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_873 = 8'h69 == io_state_in_3 ? 8'he4 : _GEN_872; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_874 = 8'h6a == io_state_in_3 ? 8'h58 : _GEN_873; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_875 = 8'h6b == io_state_in_3 ? 8'h5 : _GEN_874; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_876 = 8'h6c == io_state_in_3 ? 8'hb8 : _GEN_875; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_877 = 8'h6d == io_state_in_3 ? 8'hb3 : _GEN_876; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_878 = 8'h6e == io_state_in_3 ? 8'h45 : _GEN_877; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_879 = 8'h6f == io_state_in_3 ? 8'h6 : _GEN_878; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_880 = 8'h70 == io_state_in_3 ? 8'hd0 : _GEN_879; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_881 = 8'h71 == io_state_in_3 ? 8'h2c : _GEN_880; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_882 = 8'h72 == io_state_in_3 ? 8'h1e : _GEN_881; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_883 = 8'h73 == io_state_in_3 ? 8'h8f : _GEN_882; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_884 = 8'h74 == io_state_in_3 ? 8'hca : _GEN_883; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_885 = 8'h75 == io_state_in_3 ? 8'h3f : _GEN_884; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_886 = 8'h76 == io_state_in_3 ? 8'hf : _GEN_885; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_887 = 8'h77 == io_state_in_3 ? 8'h2 : _GEN_886; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_888 = 8'h78 == io_state_in_3 ? 8'hc1 : _GEN_887; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_889 = 8'h79 == io_state_in_3 ? 8'haf : _GEN_888; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_890 = 8'h7a == io_state_in_3 ? 8'hbd : _GEN_889; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_891 = 8'h7b == io_state_in_3 ? 8'h3 : _GEN_890; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_892 = 8'h7c == io_state_in_3 ? 8'h1 : _GEN_891; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_893 = 8'h7d == io_state_in_3 ? 8'h13 : _GEN_892; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_894 = 8'h7e == io_state_in_3 ? 8'h8a : _GEN_893; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_895 = 8'h7f == io_state_in_3 ? 8'h6b : _GEN_894; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_896 = 8'h80 == io_state_in_3 ? 8'h3a : _GEN_895; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_897 = 8'h81 == io_state_in_3 ? 8'h91 : _GEN_896; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_898 = 8'h82 == io_state_in_3 ? 8'h11 : _GEN_897; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_899 = 8'h83 == io_state_in_3 ? 8'h41 : _GEN_898; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_900 = 8'h84 == io_state_in_3 ? 8'h4f : _GEN_899; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_901 = 8'h85 == io_state_in_3 ? 8'h67 : _GEN_900; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_902 = 8'h86 == io_state_in_3 ? 8'hdc : _GEN_901; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_903 = 8'h87 == io_state_in_3 ? 8'hea : _GEN_902; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_904 = 8'h88 == io_state_in_3 ? 8'h97 : _GEN_903; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_905 = 8'h89 == io_state_in_3 ? 8'hf2 : _GEN_904; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_906 = 8'h8a == io_state_in_3 ? 8'hcf : _GEN_905; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_907 = 8'h8b == io_state_in_3 ? 8'hce : _GEN_906; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_908 = 8'h8c == io_state_in_3 ? 8'hf0 : _GEN_907; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_909 = 8'h8d == io_state_in_3 ? 8'hb4 : _GEN_908; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_910 = 8'h8e == io_state_in_3 ? 8'he6 : _GEN_909; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_911 = 8'h8f == io_state_in_3 ? 8'h73 : _GEN_910; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_912 = 8'h90 == io_state_in_3 ? 8'h96 : _GEN_911; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_913 = 8'h91 == io_state_in_3 ? 8'hac : _GEN_912; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_914 = 8'h92 == io_state_in_3 ? 8'h74 : _GEN_913; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_915 = 8'h93 == io_state_in_3 ? 8'h22 : _GEN_914; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_916 = 8'h94 == io_state_in_3 ? 8'he7 : _GEN_915; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_917 = 8'h95 == io_state_in_3 ? 8'had : _GEN_916; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_918 = 8'h96 == io_state_in_3 ? 8'h35 : _GEN_917; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_919 = 8'h97 == io_state_in_3 ? 8'h85 : _GEN_918; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_920 = 8'h98 == io_state_in_3 ? 8'he2 : _GEN_919; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_921 = 8'h99 == io_state_in_3 ? 8'hf9 : _GEN_920; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_922 = 8'h9a == io_state_in_3 ? 8'h37 : _GEN_921; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_923 = 8'h9b == io_state_in_3 ? 8'he8 : _GEN_922; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_924 = 8'h9c == io_state_in_3 ? 8'h1c : _GEN_923; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_925 = 8'h9d == io_state_in_3 ? 8'h75 : _GEN_924; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_926 = 8'h9e == io_state_in_3 ? 8'hdf : _GEN_925; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_927 = 8'h9f == io_state_in_3 ? 8'h6e : _GEN_926; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_928 = 8'ha0 == io_state_in_3 ? 8'h47 : _GEN_927; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_929 = 8'ha1 == io_state_in_3 ? 8'hf1 : _GEN_928; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_930 = 8'ha2 == io_state_in_3 ? 8'h1a : _GEN_929; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_931 = 8'ha3 == io_state_in_3 ? 8'h71 : _GEN_930; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_932 = 8'ha4 == io_state_in_3 ? 8'h1d : _GEN_931; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_933 = 8'ha5 == io_state_in_3 ? 8'h29 : _GEN_932; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_934 = 8'ha6 == io_state_in_3 ? 8'hc5 : _GEN_933; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_935 = 8'ha7 == io_state_in_3 ? 8'h89 : _GEN_934; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_936 = 8'ha8 == io_state_in_3 ? 8'h6f : _GEN_935; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_937 = 8'ha9 == io_state_in_3 ? 8'hb7 : _GEN_936; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_938 = 8'haa == io_state_in_3 ? 8'h62 : _GEN_937; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_939 = 8'hab == io_state_in_3 ? 8'he : _GEN_938; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_940 = 8'hac == io_state_in_3 ? 8'haa : _GEN_939; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_941 = 8'had == io_state_in_3 ? 8'h18 : _GEN_940; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_942 = 8'hae == io_state_in_3 ? 8'hbe : _GEN_941; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_943 = 8'haf == io_state_in_3 ? 8'h1b : _GEN_942; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_944 = 8'hb0 == io_state_in_3 ? 8'hfc : _GEN_943; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_945 = 8'hb1 == io_state_in_3 ? 8'h56 : _GEN_944; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_946 = 8'hb2 == io_state_in_3 ? 8'h3e : _GEN_945; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_947 = 8'hb3 == io_state_in_3 ? 8'h4b : _GEN_946; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_948 = 8'hb4 == io_state_in_3 ? 8'hc6 : _GEN_947; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_949 = 8'hb5 == io_state_in_3 ? 8'hd2 : _GEN_948; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_950 = 8'hb6 == io_state_in_3 ? 8'h79 : _GEN_949; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_951 = 8'hb7 == io_state_in_3 ? 8'h20 : _GEN_950; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_952 = 8'hb8 == io_state_in_3 ? 8'h9a : _GEN_951; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_953 = 8'hb9 == io_state_in_3 ? 8'hdb : _GEN_952; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_954 = 8'hba == io_state_in_3 ? 8'hc0 : _GEN_953; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_955 = 8'hbb == io_state_in_3 ? 8'hfe : _GEN_954; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_956 = 8'hbc == io_state_in_3 ? 8'h78 : _GEN_955; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_957 = 8'hbd == io_state_in_3 ? 8'hcd : _GEN_956; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_958 = 8'hbe == io_state_in_3 ? 8'h5a : _GEN_957; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_959 = 8'hbf == io_state_in_3 ? 8'hf4 : _GEN_958; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_960 = 8'hc0 == io_state_in_3 ? 8'h1f : _GEN_959; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_961 = 8'hc1 == io_state_in_3 ? 8'hdd : _GEN_960; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_962 = 8'hc2 == io_state_in_3 ? 8'ha8 : _GEN_961; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_963 = 8'hc3 == io_state_in_3 ? 8'h33 : _GEN_962; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_964 = 8'hc4 == io_state_in_3 ? 8'h88 : _GEN_963; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_965 = 8'hc5 == io_state_in_3 ? 8'h7 : _GEN_964; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_966 = 8'hc6 == io_state_in_3 ? 8'hc7 : _GEN_965; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_967 = 8'hc7 == io_state_in_3 ? 8'h31 : _GEN_966; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_968 = 8'hc8 == io_state_in_3 ? 8'hb1 : _GEN_967; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_969 = 8'hc9 == io_state_in_3 ? 8'h12 : _GEN_968; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_970 = 8'hca == io_state_in_3 ? 8'h10 : _GEN_969; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_971 = 8'hcb == io_state_in_3 ? 8'h59 : _GEN_970; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_972 = 8'hcc == io_state_in_3 ? 8'h27 : _GEN_971; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_973 = 8'hcd == io_state_in_3 ? 8'h80 : _GEN_972; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_974 = 8'hce == io_state_in_3 ? 8'hec : _GEN_973; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_975 = 8'hcf == io_state_in_3 ? 8'h5f : _GEN_974; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_976 = 8'hd0 == io_state_in_3 ? 8'h60 : _GEN_975; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_977 = 8'hd1 == io_state_in_3 ? 8'h51 : _GEN_976; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_978 = 8'hd2 == io_state_in_3 ? 8'h7f : _GEN_977; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_979 = 8'hd3 == io_state_in_3 ? 8'ha9 : _GEN_978; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_980 = 8'hd4 == io_state_in_3 ? 8'h19 : _GEN_979; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_981 = 8'hd5 == io_state_in_3 ? 8'hb5 : _GEN_980; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_982 = 8'hd6 == io_state_in_3 ? 8'h4a : _GEN_981; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_983 = 8'hd7 == io_state_in_3 ? 8'hd : _GEN_982; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_984 = 8'hd8 == io_state_in_3 ? 8'h2d : _GEN_983; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_985 = 8'hd9 == io_state_in_3 ? 8'he5 : _GEN_984; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_986 = 8'hda == io_state_in_3 ? 8'h7a : _GEN_985; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_987 = 8'hdb == io_state_in_3 ? 8'h9f : _GEN_986; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_988 = 8'hdc == io_state_in_3 ? 8'h93 : _GEN_987; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_989 = 8'hdd == io_state_in_3 ? 8'hc9 : _GEN_988; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_990 = 8'hde == io_state_in_3 ? 8'h9c : _GEN_989; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_991 = 8'hdf == io_state_in_3 ? 8'hef : _GEN_990; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_992 = 8'he0 == io_state_in_3 ? 8'ha0 : _GEN_991; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_993 = 8'he1 == io_state_in_3 ? 8'he0 : _GEN_992; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_994 = 8'he2 == io_state_in_3 ? 8'h3b : _GEN_993; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_995 = 8'he3 == io_state_in_3 ? 8'h4d : _GEN_994; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_996 = 8'he4 == io_state_in_3 ? 8'hae : _GEN_995; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_997 = 8'he5 == io_state_in_3 ? 8'h2a : _GEN_996; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_998 = 8'he6 == io_state_in_3 ? 8'hf5 : _GEN_997; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_999 = 8'he7 == io_state_in_3 ? 8'hb0 : _GEN_998; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1000 = 8'he8 == io_state_in_3 ? 8'hc8 : _GEN_999; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1001 = 8'he9 == io_state_in_3 ? 8'heb : _GEN_1000; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1002 = 8'hea == io_state_in_3 ? 8'hbb : _GEN_1001; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1003 = 8'heb == io_state_in_3 ? 8'h3c : _GEN_1002; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1004 = 8'hec == io_state_in_3 ? 8'h83 : _GEN_1003; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1005 = 8'hed == io_state_in_3 ? 8'h53 : _GEN_1004; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1006 = 8'hee == io_state_in_3 ? 8'h99 : _GEN_1005; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1007 = 8'hef == io_state_in_3 ? 8'h61 : _GEN_1006; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1008 = 8'hf0 == io_state_in_3 ? 8'h17 : _GEN_1007; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1009 = 8'hf1 == io_state_in_3 ? 8'h2b : _GEN_1008; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1010 = 8'hf2 == io_state_in_3 ? 8'h4 : _GEN_1009; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1011 = 8'hf3 == io_state_in_3 ? 8'h7e : _GEN_1010; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1012 = 8'hf4 == io_state_in_3 ? 8'hba : _GEN_1011; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1013 = 8'hf5 == io_state_in_3 ? 8'h77 : _GEN_1012; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1014 = 8'hf6 == io_state_in_3 ? 8'hd6 : _GEN_1013; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1015 = 8'hf7 == io_state_in_3 ? 8'h26 : _GEN_1014; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1016 = 8'hf8 == io_state_in_3 ? 8'he1 : _GEN_1015; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1017 = 8'hf9 == io_state_in_3 ? 8'h69 : _GEN_1016; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1018 = 8'hfa == io_state_in_3 ? 8'h14 : _GEN_1017; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1019 = 8'hfb == io_state_in_3 ? 8'h63 : _GEN_1018; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1020 = 8'hfc == io_state_in_3 ? 8'h55 : _GEN_1019; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1021 = 8'hfd == io_state_in_3 ? 8'h21 : _GEN_1020; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1022 = 8'hfe == io_state_in_3 ? 8'hc : _GEN_1021; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1025 = 8'h1 == io_state_in_4 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1026 = 8'h2 == io_state_in_4 ? 8'h6a : _GEN_1025; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1027 = 8'h3 == io_state_in_4 ? 8'hd5 : _GEN_1026; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1028 = 8'h4 == io_state_in_4 ? 8'h30 : _GEN_1027; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1029 = 8'h5 == io_state_in_4 ? 8'h36 : _GEN_1028; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1030 = 8'h6 == io_state_in_4 ? 8'ha5 : _GEN_1029; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1031 = 8'h7 == io_state_in_4 ? 8'h38 : _GEN_1030; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1032 = 8'h8 == io_state_in_4 ? 8'hbf : _GEN_1031; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1033 = 8'h9 == io_state_in_4 ? 8'h40 : _GEN_1032; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1034 = 8'ha == io_state_in_4 ? 8'ha3 : _GEN_1033; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1035 = 8'hb == io_state_in_4 ? 8'h9e : _GEN_1034; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1036 = 8'hc == io_state_in_4 ? 8'h81 : _GEN_1035; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1037 = 8'hd == io_state_in_4 ? 8'hf3 : _GEN_1036; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1038 = 8'he == io_state_in_4 ? 8'hd7 : _GEN_1037; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1039 = 8'hf == io_state_in_4 ? 8'hfb : _GEN_1038; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1040 = 8'h10 == io_state_in_4 ? 8'h7c : _GEN_1039; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1041 = 8'h11 == io_state_in_4 ? 8'he3 : _GEN_1040; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1042 = 8'h12 == io_state_in_4 ? 8'h39 : _GEN_1041; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1043 = 8'h13 == io_state_in_4 ? 8'h82 : _GEN_1042; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1044 = 8'h14 == io_state_in_4 ? 8'h9b : _GEN_1043; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1045 = 8'h15 == io_state_in_4 ? 8'h2f : _GEN_1044; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1046 = 8'h16 == io_state_in_4 ? 8'hff : _GEN_1045; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1047 = 8'h17 == io_state_in_4 ? 8'h87 : _GEN_1046; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1048 = 8'h18 == io_state_in_4 ? 8'h34 : _GEN_1047; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1049 = 8'h19 == io_state_in_4 ? 8'h8e : _GEN_1048; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1050 = 8'h1a == io_state_in_4 ? 8'h43 : _GEN_1049; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1051 = 8'h1b == io_state_in_4 ? 8'h44 : _GEN_1050; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1052 = 8'h1c == io_state_in_4 ? 8'hc4 : _GEN_1051; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1053 = 8'h1d == io_state_in_4 ? 8'hde : _GEN_1052; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1054 = 8'h1e == io_state_in_4 ? 8'he9 : _GEN_1053; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1055 = 8'h1f == io_state_in_4 ? 8'hcb : _GEN_1054; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1056 = 8'h20 == io_state_in_4 ? 8'h54 : _GEN_1055; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1057 = 8'h21 == io_state_in_4 ? 8'h7b : _GEN_1056; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1058 = 8'h22 == io_state_in_4 ? 8'h94 : _GEN_1057; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1059 = 8'h23 == io_state_in_4 ? 8'h32 : _GEN_1058; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1060 = 8'h24 == io_state_in_4 ? 8'ha6 : _GEN_1059; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1061 = 8'h25 == io_state_in_4 ? 8'hc2 : _GEN_1060; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1062 = 8'h26 == io_state_in_4 ? 8'h23 : _GEN_1061; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1063 = 8'h27 == io_state_in_4 ? 8'h3d : _GEN_1062; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1064 = 8'h28 == io_state_in_4 ? 8'hee : _GEN_1063; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1065 = 8'h29 == io_state_in_4 ? 8'h4c : _GEN_1064; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1066 = 8'h2a == io_state_in_4 ? 8'h95 : _GEN_1065; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1067 = 8'h2b == io_state_in_4 ? 8'hb : _GEN_1066; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1068 = 8'h2c == io_state_in_4 ? 8'h42 : _GEN_1067; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1069 = 8'h2d == io_state_in_4 ? 8'hfa : _GEN_1068; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1070 = 8'h2e == io_state_in_4 ? 8'hc3 : _GEN_1069; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1071 = 8'h2f == io_state_in_4 ? 8'h4e : _GEN_1070; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1072 = 8'h30 == io_state_in_4 ? 8'h8 : _GEN_1071; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1073 = 8'h31 == io_state_in_4 ? 8'h2e : _GEN_1072; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1074 = 8'h32 == io_state_in_4 ? 8'ha1 : _GEN_1073; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1075 = 8'h33 == io_state_in_4 ? 8'h66 : _GEN_1074; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1076 = 8'h34 == io_state_in_4 ? 8'h28 : _GEN_1075; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1077 = 8'h35 == io_state_in_4 ? 8'hd9 : _GEN_1076; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1078 = 8'h36 == io_state_in_4 ? 8'h24 : _GEN_1077; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1079 = 8'h37 == io_state_in_4 ? 8'hb2 : _GEN_1078; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1080 = 8'h38 == io_state_in_4 ? 8'h76 : _GEN_1079; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1081 = 8'h39 == io_state_in_4 ? 8'h5b : _GEN_1080; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1082 = 8'h3a == io_state_in_4 ? 8'ha2 : _GEN_1081; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1083 = 8'h3b == io_state_in_4 ? 8'h49 : _GEN_1082; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1084 = 8'h3c == io_state_in_4 ? 8'h6d : _GEN_1083; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1085 = 8'h3d == io_state_in_4 ? 8'h8b : _GEN_1084; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1086 = 8'h3e == io_state_in_4 ? 8'hd1 : _GEN_1085; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1087 = 8'h3f == io_state_in_4 ? 8'h25 : _GEN_1086; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1088 = 8'h40 == io_state_in_4 ? 8'h72 : _GEN_1087; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1089 = 8'h41 == io_state_in_4 ? 8'hf8 : _GEN_1088; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1090 = 8'h42 == io_state_in_4 ? 8'hf6 : _GEN_1089; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1091 = 8'h43 == io_state_in_4 ? 8'h64 : _GEN_1090; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1092 = 8'h44 == io_state_in_4 ? 8'h86 : _GEN_1091; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1093 = 8'h45 == io_state_in_4 ? 8'h68 : _GEN_1092; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1094 = 8'h46 == io_state_in_4 ? 8'h98 : _GEN_1093; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1095 = 8'h47 == io_state_in_4 ? 8'h16 : _GEN_1094; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1096 = 8'h48 == io_state_in_4 ? 8'hd4 : _GEN_1095; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1097 = 8'h49 == io_state_in_4 ? 8'ha4 : _GEN_1096; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1098 = 8'h4a == io_state_in_4 ? 8'h5c : _GEN_1097; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1099 = 8'h4b == io_state_in_4 ? 8'hcc : _GEN_1098; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1100 = 8'h4c == io_state_in_4 ? 8'h5d : _GEN_1099; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1101 = 8'h4d == io_state_in_4 ? 8'h65 : _GEN_1100; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1102 = 8'h4e == io_state_in_4 ? 8'hb6 : _GEN_1101; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1103 = 8'h4f == io_state_in_4 ? 8'h92 : _GEN_1102; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1104 = 8'h50 == io_state_in_4 ? 8'h6c : _GEN_1103; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1105 = 8'h51 == io_state_in_4 ? 8'h70 : _GEN_1104; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1106 = 8'h52 == io_state_in_4 ? 8'h48 : _GEN_1105; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1107 = 8'h53 == io_state_in_4 ? 8'h50 : _GEN_1106; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1108 = 8'h54 == io_state_in_4 ? 8'hfd : _GEN_1107; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1109 = 8'h55 == io_state_in_4 ? 8'hed : _GEN_1108; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1110 = 8'h56 == io_state_in_4 ? 8'hb9 : _GEN_1109; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1111 = 8'h57 == io_state_in_4 ? 8'hda : _GEN_1110; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1112 = 8'h58 == io_state_in_4 ? 8'h5e : _GEN_1111; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1113 = 8'h59 == io_state_in_4 ? 8'h15 : _GEN_1112; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1114 = 8'h5a == io_state_in_4 ? 8'h46 : _GEN_1113; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1115 = 8'h5b == io_state_in_4 ? 8'h57 : _GEN_1114; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1116 = 8'h5c == io_state_in_4 ? 8'ha7 : _GEN_1115; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1117 = 8'h5d == io_state_in_4 ? 8'h8d : _GEN_1116; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1118 = 8'h5e == io_state_in_4 ? 8'h9d : _GEN_1117; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1119 = 8'h5f == io_state_in_4 ? 8'h84 : _GEN_1118; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1120 = 8'h60 == io_state_in_4 ? 8'h90 : _GEN_1119; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1121 = 8'h61 == io_state_in_4 ? 8'hd8 : _GEN_1120; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1122 = 8'h62 == io_state_in_4 ? 8'hab : _GEN_1121; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1123 = 8'h63 == io_state_in_4 ? 8'h0 : _GEN_1122; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1124 = 8'h64 == io_state_in_4 ? 8'h8c : _GEN_1123; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1125 = 8'h65 == io_state_in_4 ? 8'hbc : _GEN_1124; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1126 = 8'h66 == io_state_in_4 ? 8'hd3 : _GEN_1125; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1127 = 8'h67 == io_state_in_4 ? 8'ha : _GEN_1126; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1128 = 8'h68 == io_state_in_4 ? 8'hf7 : _GEN_1127; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1129 = 8'h69 == io_state_in_4 ? 8'he4 : _GEN_1128; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1130 = 8'h6a == io_state_in_4 ? 8'h58 : _GEN_1129; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1131 = 8'h6b == io_state_in_4 ? 8'h5 : _GEN_1130; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1132 = 8'h6c == io_state_in_4 ? 8'hb8 : _GEN_1131; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1133 = 8'h6d == io_state_in_4 ? 8'hb3 : _GEN_1132; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1134 = 8'h6e == io_state_in_4 ? 8'h45 : _GEN_1133; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1135 = 8'h6f == io_state_in_4 ? 8'h6 : _GEN_1134; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1136 = 8'h70 == io_state_in_4 ? 8'hd0 : _GEN_1135; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1137 = 8'h71 == io_state_in_4 ? 8'h2c : _GEN_1136; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1138 = 8'h72 == io_state_in_4 ? 8'h1e : _GEN_1137; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1139 = 8'h73 == io_state_in_4 ? 8'h8f : _GEN_1138; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1140 = 8'h74 == io_state_in_4 ? 8'hca : _GEN_1139; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1141 = 8'h75 == io_state_in_4 ? 8'h3f : _GEN_1140; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1142 = 8'h76 == io_state_in_4 ? 8'hf : _GEN_1141; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1143 = 8'h77 == io_state_in_4 ? 8'h2 : _GEN_1142; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1144 = 8'h78 == io_state_in_4 ? 8'hc1 : _GEN_1143; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1145 = 8'h79 == io_state_in_4 ? 8'haf : _GEN_1144; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1146 = 8'h7a == io_state_in_4 ? 8'hbd : _GEN_1145; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1147 = 8'h7b == io_state_in_4 ? 8'h3 : _GEN_1146; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1148 = 8'h7c == io_state_in_4 ? 8'h1 : _GEN_1147; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1149 = 8'h7d == io_state_in_4 ? 8'h13 : _GEN_1148; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1150 = 8'h7e == io_state_in_4 ? 8'h8a : _GEN_1149; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1151 = 8'h7f == io_state_in_4 ? 8'h6b : _GEN_1150; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1152 = 8'h80 == io_state_in_4 ? 8'h3a : _GEN_1151; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1153 = 8'h81 == io_state_in_4 ? 8'h91 : _GEN_1152; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1154 = 8'h82 == io_state_in_4 ? 8'h11 : _GEN_1153; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1155 = 8'h83 == io_state_in_4 ? 8'h41 : _GEN_1154; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1156 = 8'h84 == io_state_in_4 ? 8'h4f : _GEN_1155; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1157 = 8'h85 == io_state_in_4 ? 8'h67 : _GEN_1156; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1158 = 8'h86 == io_state_in_4 ? 8'hdc : _GEN_1157; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1159 = 8'h87 == io_state_in_4 ? 8'hea : _GEN_1158; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1160 = 8'h88 == io_state_in_4 ? 8'h97 : _GEN_1159; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1161 = 8'h89 == io_state_in_4 ? 8'hf2 : _GEN_1160; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1162 = 8'h8a == io_state_in_4 ? 8'hcf : _GEN_1161; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1163 = 8'h8b == io_state_in_4 ? 8'hce : _GEN_1162; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1164 = 8'h8c == io_state_in_4 ? 8'hf0 : _GEN_1163; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1165 = 8'h8d == io_state_in_4 ? 8'hb4 : _GEN_1164; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1166 = 8'h8e == io_state_in_4 ? 8'he6 : _GEN_1165; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1167 = 8'h8f == io_state_in_4 ? 8'h73 : _GEN_1166; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1168 = 8'h90 == io_state_in_4 ? 8'h96 : _GEN_1167; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1169 = 8'h91 == io_state_in_4 ? 8'hac : _GEN_1168; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1170 = 8'h92 == io_state_in_4 ? 8'h74 : _GEN_1169; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1171 = 8'h93 == io_state_in_4 ? 8'h22 : _GEN_1170; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1172 = 8'h94 == io_state_in_4 ? 8'he7 : _GEN_1171; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1173 = 8'h95 == io_state_in_4 ? 8'had : _GEN_1172; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1174 = 8'h96 == io_state_in_4 ? 8'h35 : _GEN_1173; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1175 = 8'h97 == io_state_in_4 ? 8'h85 : _GEN_1174; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1176 = 8'h98 == io_state_in_4 ? 8'he2 : _GEN_1175; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1177 = 8'h99 == io_state_in_4 ? 8'hf9 : _GEN_1176; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1178 = 8'h9a == io_state_in_4 ? 8'h37 : _GEN_1177; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1179 = 8'h9b == io_state_in_4 ? 8'he8 : _GEN_1178; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1180 = 8'h9c == io_state_in_4 ? 8'h1c : _GEN_1179; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1181 = 8'h9d == io_state_in_4 ? 8'h75 : _GEN_1180; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1182 = 8'h9e == io_state_in_4 ? 8'hdf : _GEN_1181; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1183 = 8'h9f == io_state_in_4 ? 8'h6e : _GEN_1182; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1184 = 8'ha0 == io_state_in_4 ? 8'h47 : _GEN_1183; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1185 = 8'ha1 == io_state_in_4 ? 8'hf1 : _GEN_1184; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1186 = 8'ha2 == io_state_in_4 ? 8'h1a : _GEN_1185; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1187 = 8'ha3 == io_state_in_4 ? 8'h71 : _GEN_1186; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1188 = 8'ha4 == io_state_in_4 ? 8'h1d : _GEN_1187; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1189 = 8'ha5 == io_state_in_4 ? 8'h29 : _GEN_1188; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1190 = 8'ha6 == io_state_in_4 ? 8'hc5 : _GEN_1189; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1191 = 8'ha7 == io_state_in_4 ? 8'h89 : _GEN_1190; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1192 = 8'ha8 == io_state_in_4 ? 8'h6f : _GEN_1191; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1193 = 8'ha9 == io_state_in_4 ? 8'hb7 : _GEN_1192; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1194 = 8'haa == io_state_in_4 ? 8'h62 : _GEN_1193; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1195 = 8'hab == io_state_in_4 ? 8'he : _GEN_1194; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1196 = 8'hac == io_state_in_4 ? 8'haa : _GEN_1195; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1197 = 8'had == io_state_in_4 ? 8'h18 : _GEN_1196; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1198 = 8'hae == io_state_in_4 ? 8'hbe : _GEN_1197; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1199 = 8'haf == io_state_in_4 ? 8'h1b : _GEN_1198; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1200 = 8'hb0 == io_state_in_4 ? 8'hfc : _GEN_1199; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1201 = 8'hb1 == io_state_in_4 ? 8'h56 : _GEN_1200; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1202 = 8'hb2 == io_state_in_4 ? 8'h3e : _GEN_1201; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1203 = 8'hb3 == io_state_in_4 ? 8'h4b : _GEN_1202; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1204 = 8'hb4 == io_state_in_4 ? 8'hc6 : _GEN_1203; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1205 = 8'hb5 == io_state_in_4 ? 8'hd2 : _GEN_1204; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1206 = 8'hb6 == io_state_in_4 ? 8'h79 : _GEN_1205; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1207 = 8'hb7 == io_state_in_4 ? 8'h20 : _GEN_1206; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1208 = 8'hb8 == io_state_in_4 ? 8'h9a : _GEN_1207; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1209 = 8'hb9 == io_state_in_4 ? 8'hdb : _GEN_1208; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1210 = 8'hba == io_state_in_4 ? 8'hc0 : _GEN_1209; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1211 = 8'hbb == io_state_in_4 ? 8'hfe : _GEN_1210; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1212 = 8'hbc == io_state_in_4 ? 8'h78 : _GEN_1211; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1213 = 8'hbd == io_state_in_4 ? 8'hcd : _GEN_1212; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1214 = 8'hbe == io_state_in_4 ? 8'h5a : _GEN_1213; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1215 = 8'hbf == io_state_in_4 ? 8'hf4 : _GEN_1214; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1216 = 8'hc0 == io_state_in_4 ? 8'h1f : _GEN_1215; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1217 = 8'hc1 == io_state_in_4 ? 8'hdd : _GEN_1216; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1218 = 8'hc2 == io_state_in_4 ? 8'ha8 : _GEN_1217; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1219 = 8'hc3 == io_state_in_4 ? 8'h33 : _GEN_1218; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1220 = 8'hc4 == io_state_in_4 ? 8'h88 : _GEN_1219; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1221 = 8'hc5 == io_state_in_4 ? 8'h7 : _GEN_1220; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1222 = 8'hc6 == io_state_in_4 ? 8'hc7 : _GEN_1221; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1223 = 8'hc7 == io_state_in_4 ? 8'h31 : _GEN_1222; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1224 = 8'hc8 == io_state_in_4 ? 8'hb1 : _GEN_1223; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1225 = 8'hc9 == io_state_in_4 ? 8'h12 : _GEN_1224; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1226 = 8'hca == io_state_in_4 ? 8'h10 : _GEN_1225; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1227 = 8'hcb == io_state_in_4 ? 8'h59 : _GEN_1226; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1228 = 8'hcc == io_state_in_4 ? 8'h27 : _GEN_1227; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1229 = 8'hcd == io_state_in_4 ? 8'h80 : _GEN_1228; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1230 = 8'hce == io_state_in_4 ? 8'hec : _GEN_1229; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1231 = 8'hcf == io_state_in_4 ? 8'h5f : _GEN_1230; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1232 = 8'hd0 == io_state_in_4 ? 8'h60 : _GEN_1231; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1233 = 8'hd1 == io_state_in_4 ? 8'h51 : _GEN_1232; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1234 = 8'hd2 == io_state_in_4 ? 8'h7f : _GEN_1233; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1235 = 8'hd3 == io_state_in_4 ? 8'ha9 : _GEN_1234; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1236 = 8'hd4 == io_state_in_4 ? 8'h19 : _GEN_1235; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1237 = 8'hd5 == io_state_in_4 ? 8'hb5 : _GEN_1236; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1238 = 8'hd6 == io_state_in_4 ? 8'h4a : _GEN_1237; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1239 = 8'hd7 == io_state_in_4 ? 8'hd : _GEN_1238; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1240 = 8'hd8 == io_state_in_4 ? 8'h2d : _GEN_1239; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1241 = 8'hd9 == io_state_in_4 ? 8'he5 : _GEN_1240; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1242 = 8'hda == io_state_in_4 ? 8'h7a : _GEN_1241; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1243 = 8'hdb == io_state_in_4 ? 8'h9f : _GEN_1242; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1244 = 8'hdc == io_state_in_4 ? 8'h93 : _GEN_1243; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1245 = 8'hdd == io_state_in_4 ? 8'hc9 : _GEN_1244; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1246 = 8'hde == io_state_in_4 ? 8'h9c : _GEN_1245; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1247 = 8'hdf == io_state_in_4 ? 8'hef : _GEN_1246; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1248 = 8'he0 == io_state_in_4 ? 8'ha0 : _GEN_1247; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1249 = 8'he1 == io_state_in_4 ? 8'he0 : _GEN_1248; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1250 = 8'he2 == io_state_in_4 ? 8'h3b : _GEN_1249; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1251 = 8'he3 == io_state_in_4 ? 8'h4d : _GEN_1250; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1252 = 8'he4 == io_state_in_4 ? 8'hae : _GEN_1251; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1253 = 8'he5 == io_state_in_4 ? 8'h2a : _GEN_1252; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1254 = 8'he6 == io_state_in_4 ? 8'hf5 : _GEN_1253; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1255 = 8'he7 == io_state_in_4 ? 8'hb0 : _GEN_1254; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1256 = 8'he8 == io_state_in_4 ? 8'hc8 : _GEN_1255; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1257 = 8'he9 == io_state_in_4 ? 8'heb : _GEN_1256; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1258 = 8'hea == io_state_in_4 ? 8'hbb : _GEN_1257; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1259 = 8'heb == io_state_in_4 ? 8'h3c : _GEN_1258; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1260 = 8'hec == io_state_in_4 ? 8'h83 : _GEN_1259; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1261 = 8'hed == io_state_in_4 ? 8'h53 : _GEN_1260; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1262 = 8'hee == io_state_in_4 ? 8'h99 : _GEN_1261; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1263 = 8'hef == io_state_in_4 ? 8'h61 : _GEN_1262; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1264 = 8'hf0 == io_state_in_4 ? 8'h17 : _GEN_1263; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1265 = 8'hf1 == io_state_in_4 ? 8'h2b : _GEN_1264; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1266 = 8'hf2 == io_state_in_4 ? 8'h4 : _GEN_1265; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1267 = 8'hf3 == io_state_in_4 ? 8'h7e : _GEN_1266; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1268 = 8'hf4 == io_state_in_4 ? 8'hba : _GEN_1267; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1269 = 8'hf5 == io_state_in_4 ? 8'h77 : _GEN_1268; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1270 = 8'hf6 == io_state_in_4 ? 8'hd6 : _GEN_1269; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1271 = 8'hf7 == io_state_in_4 ? 8'h26 : _GEN_1270; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1272 = 8'hf8 == io_state_in_4 ? 8'he1 : _GEN_1271; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1273 = 8'hf9 == io_state_in_4 ? 8'h69 : _GEN_1272; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1274 = 8'hfa == io_state_in_4 ? 8'h14 : _GEN_1273; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1275 = 8'hfb == io_state_in_4 ? 8'h63 : _GEN_1274; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1276 = 8'hfc == io_state_in_4 ? 8'h55 : _GEN_1275; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1277 = 8'hfd == io_state_in_4 ? 8'h21 : _GEN_1276; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1278 = 8'hfe == io_state_in_4 ? 8'hc : _GEN_1277; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1281 = 8'h1 == io_state_in_5 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1282 = 8'h2 == io_state_in_5 ? 8'h6a : _GEN_1281; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1283 = 8'h3 == io_state_in_5 ? 8'hd5 : _GEN_1282; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1284 = 8'h4 == io_state_in_5 ? 8'h30 : _GEN_1283; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1285 = 8'h5 == io_state_in_5 ? 8'h36 : _GEN_1284; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1286 = 8'h6 == io_state_in_5 ? 8'ha5 : _GEN_1285; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1287 = 8'h7 == io_state_in_5 ? 8'h38 : _GEN_1286; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1288 = 8'h8 == io_state_in_5 ? 8'hbf : _GEN_1287; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1289 = 8'h9 == io_state_in_5 ? 8'h40 : _GEN_1288; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1290 = 8'ha == io_state_in_5 ? 8'ha3 : _GEN_1289; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1291 = 8'hb == io_state_in_5 ? 8'h9e : _GEN_1290; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1292 = 8'hc == io_state_in_5 ? 8'h81 : _GEN_1291; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1293 = 8'hd == io_state_in_5 ? 8'hf3 : _GEN_1292; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1294 = 8'he == io_state_in_5 ? 8'hd7 : _GEN_1293; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1295 = 8'hf == io_state_in_5 ? 8'hfb : _GEN_1294; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1296 = 8'h10 == io_state_in_5 ? 8'h7c : _GEN_1295; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1297 = 8'h11 == io_state_in_5 ? 8'he3 : _GEN_1296; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1298 = 8'h12 == io_state_in_5 ? 8'h39 : _GEN_1297; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1299 = 8'h13 == io_state_in_5 ? 8'h82 : _GEN_1298; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1300 = 8'h14 == io_state_in_5 ? 8'h9b : _GEN_1299; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1301 = 8'h15 == io_state_in_5 ? 8'h2f : _GEN_1300; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1302 = 8'h16 == io_state_in_5 ? 8'hff : _GEN_1301; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1303 = 8'h17 == io_state_in_5 ? 8'h87 : _GEN_1302; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1304 = 8'h18 == io_state_in_5 ? 8'h34 : _GEN_1303; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1305 = 8'h19 == io_state_in_5 ? 8'h8e : _GEN_1304; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1306 = 8'h1a == io_state_in_5 ? 8'h43 : _GEN_1305; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1307 = 8'h1b == io_state_in_5 ? 8'h44 : _GEN_1306; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1308 = 8'h1c == io_state_in_5 ? 8'hc4 : _GEN_1307; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1309 = 8'h1d == io_state_in_5 ? 8'hde : _GEN_1308; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1310 = 8'h1e == io_state_in_5 ? 8'he9 : _GEN_1309; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1311 = 8'h1f == io_state_in_5 ? 8'hcb : _GEN_1310; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1312 = 8'h20 == io_state_in_5 ? 8'h54 : _GEN_1311; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1313 = 8'h21 == io_state_in_5 ? 8'h7b : _GEN_1312; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1314 = 8'h22 == io_state_in_5 ? 8'h94 : _GEN_1313; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1315 = 8'h23 == io_state_in_5 ? 8'h32 : _GEN_1314; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1316 = 8'h24 == io_state_in_5 ? 8'ha6 : _GEN_1315; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1317 = 8'h25 == io_state_in_5 ? 8'hc2 : _GEN_1316; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1318 = 8'h26 == io_state_in_5 ? 8'h23 : _GEN_1317; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1319 = 8'h27 == io_state_in_5 ? 8'h3d : _GEN_1318; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1320 = 8'h28 == io_state_in_5 ? 8'hee : _GEN_1319; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1321 = 8'h29 == io_state_in_5 ? 8'h4c : _GEN_1320; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1322 = 8'h2a == io_state_in_5 ? 8'h95 : _GEN_1321; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1323 = 8'h2b == io_state_in_5 ? 8'hb : _GEN_1322; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1324 = 8'h2c == io_state_in_5 ? 8'h42 : _GEN_1323; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1325 = 8'h2d == io_state_in_5 ? 8'hfa : _GEN_1324; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1326 = 8'h2e == io_state_in_5 ? 8'hc3 : _GEN_1325; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1327 = 8'h2f == io_state_in_5 ? 8'h4e : _GEN_1326; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1328 = 8'h30 == io_state_in_5 ? 8'h8 : _GEN_1327; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1329 = 8'h31 == io_state_in_5 ? 8'h2e : _GEN_1328; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1330 = 8'h32 == io_state_in_5 ? 8'ha1 : _GEN_1329; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1331 = 8'h33 == io_state_in_5 ? 8'h66 : _GEN_1330; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1332 = 8'h34 == io_state_in_5 ? 8'h28 : _GEN_1331; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1333 = 8'h35 == io_state_in_5 ? 8'hd9 : _GEN_1332; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1334 = 8'h36 == io_state_in_5 ? 8'h24 : _GEN_1333; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1335 = 8'h37 == io_state_in_5 ? 8'hb2 : _GEN_1334; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1336 = 8'h38 == io_state_in_5 ? 8'h76 : _GEN_1335; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1337 = 8'h39 == io_state_in_5 ? 8'h5b : _GEN_1336; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1338 = 8'h3a == io_state_in_5 ? 8'ha2 : _GEN_1337; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1339 = 8'h3b == io_state_in_5 ? 8'h49 : _GEN_1338; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1340 = 8'h3c == io_state_in_5 ? 8'h6d : _GEN_1339; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1341 = 8'h3d == io_state_in_5 ? 8'h8b : _GEN_1340; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1342 = 8'h3e == io_state_in_5 ? 8'hd1 : _GEN_1341; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1343 = 8'h3f == io_state_in_5 ? 8'h25 : _GEN_1342; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1344 = 8'h40 == io_state_in_5 ? 8'h72 : _GEN_1343; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1345 = 8'h41 == io_state_in_5 ? 8'hf8 : _GEN_1344; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1346 = 8'h42 == io_state_in_5 ? 8'hf6 : _GEN_1345; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1347 = 8'h43 == io_state_in_5 ? 8'h64 : _GEN_1346; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1348 = 8'h44 == io_state_in_5 ? 8'h86 : _GEN_1347; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1349 = 8'h45 == io_state_in_5 ? 8'h68 : _GEN_1348; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1350 = 8'h46 == io_state_in_5 ? 8'h98 : _GEN_1349; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1351 = 8'h47 == io_state_in_5 ? 8'h16 : _GEN_1350; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1352 = 8'h48 == io_state_in_5 ? 8'hd4 : _GEN_1351; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1353 = 8'h49 == io_state_in_5 ? 8'ha4 : _GEN_1352; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1354 = 8'h4a == io_state_in_5 ? 8'h5c : _GEN_1353; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1355 = 8'h4b == io_state_in_5 ? 8'hcc : _GEN_1354; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1356 = 8'h4c == io_state_in_5 ? 8'h5d : _GEN_1355; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1357 = 8'h4d == io_state_in_5 ? 8'h65 : _GEN_1356; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1358 = 8'h4e == io_state_in_5 ? 8'hb6 : _GEN_1357; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1359 = 8'h4f == io_state_in_5 ? 8'h92 : _GEN_1358; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1360 = 8'h50 == io_state_in_5 ? 8'h6c : _GEN_1359; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1361 = 8'h51 == io_state_in_5 ? 8'h70 : _GEN_1360; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1362 = 8'h52 == io_state_in_5 ? 8'h48 : _GEN_1361; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1363 = 8'h53 == io_state_in_5 ? 8'h50 : _GEN_1362; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1364 = 8'h54 == io_state_in_5 ? 8'hfd : _GEN_1363; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1365 = 8'h55 == io_state_in_5 ? 8'hed : _GEN_1364; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1366 = 8'h56 == io_state_in_5 ? 8'hb9 : _GEN_1365; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1367 = 8'h57 == io_state_in_5 ? 8'hda : _GEN_1366; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1368 = 8'h58 == io_state_in_5 ? 8'h5e : _GEN_1367; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1369 = 8'h59 == io_state_in_5 ? 8'h15 : _GEN_1368; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1370 = 8'h5a == io_state_in_5 ? 8'h46 : _GEN_1369; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1371 = 8'h5b == io_state_in_5 ? 8'h57 : _GEN_1370; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1372 = 8'h5c == io_state_in_5 ? 8'ha7 : _GEN_1371; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1373 = 8'h5d == io_state_in_5 ? 8'h8d : _GEN_1372; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1374 = 8'h5e == io_state_in_5 ? 8'h9d : _GEN_1373; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1375 = 8'h5f == io_state_in_5 ? 8'h84 : _GEN_1374; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1376 = 8'h60 == io_state_in_5 ? 8'h90 : _GEN_1375; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1377 = 8'h61 == io_state_in_5 ? 8'hd8 : _GEN_1376; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1378 = 8'h62 == io_state_in_5 ? 8'hab : _GEN_1377; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1379 = 8'h63 == io_state_in_5 ? 8'h0 : _GEN_1378; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1380 = 8'h64 == io_state_in_5 ? 8'h8c : _GEN_1379; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1381 = 8'h65 == io_state_in_5 ? 8'hbc : _GEN_1380; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1382 = 8'h66 == io_state_in_5 ? 8'hd3 : _GEN_1381; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1383 = 8'h67 == io_state_in_5 ? 8'ha : _GEN_1382; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1384 = 8'h68 == io_state_in_5 ? 8'hf7 : _GEN_1383; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1385 = 8'h69 == io_state_in_5 ? 8'he4 : _GEN_1384; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1386 = 8'h6a == io_state_in_5 ? 8'h58 : _GEN_1385; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1387 = 8'h6b == io_state_in_5 ? 8'h5 : _GEN_1386; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1388 = 8'h6c == io_state_in_5 ? 8'hb8 : _GEN_1387; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1389 = 8'h6d == io_state_in_5 ? 8'hb3 : _GEN_1388; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1390 = 8'h6e == io_state_in_5 ? 8'h45 : _GEN_1389; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1391 = 8'h6f == io_state_in_5 ? 8'h6 : _GEN_1390; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1392 = 8'h70 == io_state_in_5 ? 8'hd0 : _GEN_1391; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1393 = 8'h71 == io_state_in_5 ? 8'h2c : _GEN_1392; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1394 = 8'h72 == io_state_in_5 ? 8'h1e : _GEN_1393; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1395 = 8'h73 == io_state_in_5 ? 8'h8f : _GEN_1394; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1396 = 8'h74 == io_state_in_5 ? 8'hca : _GEN_1395; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1397 = 8'h75 == io_state_in_5 ? 8'h3f : _GEN_1396; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1398 = 8'h76 == io_state_in_5 ? 8'hf : _GEN_1397; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1399 = 8'h77 == io_state_in_5 ? 8'h2 : _GEN_1398; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1400 = 8'h78 == io_state_in_5 ? 8'hc1 : _GEN_1399; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1401 = 8'h79 == io_state_in_5 ? 8'haf : _GEN_1400; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1402 = 8'h7a == io_state_in_5 ? 8'hbd : _GEN_1401; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1403 = 8'h7b == io_state_in_5 ? 8'h3 : _GEN_1402; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1404 = 8'h7c == io_state_in_5 ? 8'h1 : _GEN_1403; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1405 = 8'h7d == io_state_in_5 ? 8'h13 : _GEN_1404; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1406 = 8'h7e == io_state_in_5 ? 8'h8a : _GEN_1405; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1407 = 8'h7f == io_state_in_5 ? 8'h6b : _GEN_1406; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1408 = 8'h80 == io_state_in_5 ? 8'h3a : _GEN_1407; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1409 = 8'h81 == io_state_in_5 ? 8'h91 : _GEN_1408; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1410 = 8'h82 == io_state_in_5 ? 8'h11 : _GEN_1409; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1411 = 8'h83 == io_state_in_5 ? 8'h41 : _GEN_1410; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1412 = 8'h84 == io_state_in_5 ? 8'h4f : _GEN_1411; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1413 = 8'h85 == io_state_in_5 ? 8'h67 : _GEN_1412; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1414 = 8'h86 == io_state_in_5 ? 8'hdc : _GEN_1413; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1415 = 8'h87 == io_state_in_5 ? 8'hea : _GEN_1414; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1416 = 8'h88 == io_state_in_5 ? 8'h97 : _GEN_1415; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1417 = 8'h89 == io_state_in_5 ? 8'hf2 : _GEN_1416; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1418 = 8'h8a == io_state_in_5 ? 8'hcf : _GEN_1417; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1419 = 8'h8b == io_state_in_5 ? 8'hce : _GEN_1418; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1420 = 8'h8c == io_state_in_5 ? 8'hf0 : _GEN_1419; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1421 = 8'h8d == io_state_in_5 ? 8'hb4 : _GEN_1420; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1422 = 8'h8e == io_state_in_5 ? 8'he6 : _GEN_1421; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1423 = 8'h8f == io_state_in_5 ? 8'h73 : _GEN_1422; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1424 = 8'h90 == io_state_in_5 ? 8'h96 : _GEN_1423; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1425 = 8'h91 == io_state_in_5 ? 8'hac : _GEN_1424; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1426 = 8'h92 == io_state_in_5 ? 8'h74 : _GEN_1425; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1427 = 8'h93 == io_state_in_5 ? 8'h22 : _GEN_1426; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1428 = 8'h94 == io_state_in_5 ? 8'he7 : _GEN_1427; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1429 = 8'h95 == io_state_in_5 ? 8'had : _GEN_1428; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1430 = 8'h96 == io_state_in_5 ? 8'h35 : _GEN_1429; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1431 = 8'h97 == io_state_in_5 ? 8'h85 : _GEN_1430; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1432 = 8'h98 == io_state_in_5 ? 8'he2 : _GEN_1431; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1433 = 8'h99 == io_state_in_5 ? 8'hf9 : _GEN_1432; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1434 = 8'h9a == io_state_in_5 ? 8'h37 : _GEN_1433; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1435 = 8'h9b == io_state_in_5 ? 8'he8 : _GEN_1434; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1436 = 8'h9c == io_state_in_5 ? 8'h1c : _GEN_1435; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1437 = 8'h9d == io_state_in_5 ? 8'h75 : _GEN_1436; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1438 = 8'h9e == io_state_in_5 ? 8'hdf : _GEN_1437; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1439 = 8'h9f == io_state_in_5 ? 8'h6e : _GEN_1438; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1440 = 8'ha0 == io_state_in_5 ? 8'h47 : _GEN_1439; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1441 = 8'ha1 == io_state_in_5 ? 8'hf1 : _GEN_1440; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1442 = 8'ha2 == io_state_in_5 ? 8'h1a : _GEN_1441; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1443 = 8'ha3 == io_state_in_5 ? 8'h71 : _GEN_1442; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1444 = 8'ha4 == io_state_in_5 ? 8'h1d : _GEN_1443; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1445 = 8'ha5 == io_state_in_5 ? 8'h29 : _GEN_1444; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1446 = 8'ha6 == io_state_in_5 ? 8'hc5 : _GEN_1445; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1447 = 8'ha7 == io_state_in_5 ? 8'h89 : _GEN_1446; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1448 = 8'ha8 == io_state_in_5 ? 8'h6f : _GEN_1447; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1449 = 8'ha9 == io_state_in_5 ? 8'hb7 : _GEN_1448; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1450 = 8'haa == io_state_in_5 ? 8'h62 : _GEN_1449; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1451 = 8'hab == io_state_in_5 ? 8'he : _GEN_1450; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1452 = 8'hac == io_state_in_5 ? 8'haa : _GEN_1451; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1453 = 8'had == io_state_in_5 ? 8'h18 : _GEN_1452; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1454 = 8'hae == io_state_in_5 ? 8'hbe : _GEN_1453; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1455 = 8'haf == io_state_in_5 ? 8'h1b : _GEN_1454; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1456 = 8'hb0 == io_state_in_5 ? 8'hfc : _GEN_1455; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1457 = 8'hb1 == io_state_in_5 ? 8'h56 : _GEN_1456; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1458 = 8'hb2 == io_state_in_5 ? 8'h3e : _GEN_1457; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1459 = 8'hb3 == io_state_in_5 ? 8'h4b : _GEN_1458; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1460 = 8'hb4 == io_state_in_5 ? 8'hc6 : _GEN_1459; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1461 = 8'hb5 == io_state_in_5 ? 8'hd2 : _GEN_1460; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1462 = 8'hb6 == io_state_in_5 ? 8'h79 : _GEN_1461; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1463 = 8'hb7 == io_state_in_5 ? 8'h20 : _GEN_1462; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1464 = 8'hb8 == io_state_in_5 ? 8'h9a : _GEN_1463; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1465 = 8'hb9 == io_state_in_5 ? 8'hdb : _GEN_1464; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1466 = 8'hba == io_state_in_5 ? 8'hc0 : _GEN_1465; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1467 = 8'hbb == io_state_in_5 ? 8'hfe : _GEN_1466; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1468 = 8'hbc == io_state_in_5 ? 8'h78 : _GEN_1467; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1469 = 8'hbd == io_state_in_5 ? 8'hcd : _GEN_1468; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1470 = 8'hbe == io_state_in_5 ? 8'h5a : _GEN_1469; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1471 = 8'hbf == io_state_in_5 ? 8'hf4 : _GEN_1470; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1472 = 8'hc0 == io_state_in_5 ? 8'h1f : _GEN_1471; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1473 = 8'hc1 == io_state_in_5 ? 8'hdd : _GEN_1472; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1474 = 8'hc2 == io_state_in_5 ? 8'ha8 : _GEN_1473; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1475 = 8'hc3 == io_state_in_5 ? 8'h33 : _GEN_1474; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1476 = 8'hc4 == io_state_in_5 ? 8'h88 : _GEN_1475; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1477 = 8'hc5 == io_state_in_5 ? 8'h7 : _GEN_1476; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1478 = 8'hc6 == io_state_in_5 ? 8'hc7 : _GEN_1477; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1479 = 8'hc7 == io_state_in_5 ? 8'h31 : _GEN_1478; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1480 = 8'hc8 == io_state_in_5 ? 8'hb1 : _GEN_1479; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1481 = 8'hc9 == io_state_in_5 ? 8'h12 : _GEN_1480; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1482 = 8'hca == io_state_in_5 ? 8'h10 : _GEN_1481; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1483 = 8'hcb == io_state_in_5 ? 8'h59 : _GEN_1482; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1484 = 8'hcc == io_state_in_5 ? 8'h27 : _GEN_1483; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1485 = 8'hcd == io_state_in_5 ? 8'h80 : _GEN_1484; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1486 = 8'hce == io_state_in_5 ? 8'hec : _GEN_1485; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1487 = 8'hcf == io_state_in_5 ? 8'h5f : _GEN_1486; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1488 = 8'hd0 == io_state_in_5 ? 8'h60 : _GEN_1487; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1489 = 8'hd1 == io_state_in_5 ? 8'h51 : _GEN_1488; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1490 = 8'hd2 == io_state_in_5 ? 8'h7f : _GEN_1489; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1491 = 8'hd3 == io_state_in_5 ? 8'ha9 : _GEN_1490; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1492 = 8'hd4 == io_state_in_5 ? 8'h19 : _GEN_1491; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1493 = 8'hd5 == io_state_in_5 ? 8'hb5 : _GEN_1492; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1494 = 8'hd6 == io_state_in_5 ? 8'h4a : _GEN_1493; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1495 = 8'hd7 == io_state_in_5 ? 8'hd : _GEN_1494; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1496 = 8'hd8 == io_state_in_5 ? 8'h2d : _GEN_1495; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1497 = 8'hd9 == io_state_in_5 ? 8'he5 : _GEN_1496; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1498 = 8'hda == io_state_in_5 ? 8'h7a : _GEN_1497; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1499 = 8'hdb == io_state_in_5 ? 8'h9f : _GEN_1498; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1500 = 8'hdc == io_state_in_5 ? 8'h93 : _GEN_1499; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1501 = 8'hdd == io_state_in_5 ? 8'hc9 : _GEN_1500; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1502 = 8'hde == io_state_in_5 ? 8'h9c : _GEN_1501; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1503 = 8'hdf == io_state_in_5 ? 8'hef : _GEN_1502; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1504 = 8'he0 == io_state_in_5 ? 8'ha0 : _GEN_1503; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1505 = 8'he1 == io_state_in_5 ? 8'he0 : _GEN_1504; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1506 = 8'he2 == io_state_in_5 ? 8'h3b : _GEN_1505; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1507 = 8'he3 == io_state_in_5 ? 8'h4d : _GEN_1506; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1508 = 8'he4 == io_state_in_5 ? 8'hae : _GEN_1507; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1509 = 8'he5 == io_state_in_5 ? 8'h2a : _GEN_1508; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1510 = 8'he6 == io_state_in_5 ? 8'hf5 : _GEN_1509; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1511 = 8'he7 == io_state_in_5 ? 8'hb0 : _GEN_1510; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1512 = 8'he8 == io_state_in_5 ? 8'hc8 : _GEN_1511; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1513 = 8'he9 == io_state_in_5 ? 8'heb : _GEN_1512; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1514 = 8'hea == io_state_in_5 ? 8'hbb : _GEN_1513; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1515 = 8'heb == io_state_in_5 ? 8'h3c : _GEN_1514; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1516 = 8'hec == io_state_in_5 ? 8'h83 : _GEN_1515; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1517 = 8'hed == io_state_in_5 ? 8'h53 : _GEN_1516; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1518 = 8'hee == io_state_in_5 ? 8'h99 : _GEN_1517; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1519 = 8'hef == io_state_in_5 ? 8'h61 : _GEN_1518; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1520 = 8'hf0 == io_state_in_5 ? 8'h17 : _GEN_1519; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1521 = 8'hf1 == io_state_in_5 ? 8'h2b : _GEN_1520; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1522 = 8'hf2 == io_state_in_5 ? 8'h4 : _GEN_1521; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1523 = 8'hf3 == io_state_in_5 ? 8'h7e : _GEN_1522; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1524 = 8'hf4 == io_state_in_5 ? 8'hba : _GEN_1523; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1525 = 8'hf5 == io_state_in_5 ? 8'h77 : _GEN_1524; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1526 = 8'hf6 == io_state_in_5 ? 8'hd6 : _GEN_1525; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1527 = 8'hf7 == io_state_in_5 ? 8'h26 : _GEN_1526; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1528 = 8'hf8 == io_state_in_5 ? 8'he1 : _GEN_1527; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1529 = 8'hf9 == io_state_in_5 ? 8'h69 : _GEN_1528; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1530 = 8'hfa == io_state_in_5 ? 8'h14 : _GEN_1529; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1531 = 8'hfb == io_state_in_5 ? 8'h63 : _GEN_1530; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1532 = 8'hfc == io_state_in_5 ? 8'h55 : _GEN_1531; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1533 = 8'hfd == io_state_in_5 ? 8'h21 : _GEN_1532; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1534 = 8'hfe == io_state_in_5 ? 8'hc : _GEN_1533; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1537 = 8'h1 == io_state_in_6 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1538 = 8'h2 == io_state_in_6 ? 8'h6a : _GEN_1537; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1539 = 8'h3 == io_state_in_6 ? 8'hd5 : _GEN_1538; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1540 = 8'h4 == io_state_in_6 ? 8'h30 : _GEN_1539; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1541 = 8'h5 == io_state_in_6 ? 8'h36 : _GEN_1540; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1542 = 8'h6 == io_state_in_6 ? 8'ha5 : _GEN_1541; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1543 = 8'h7 == io_state_in_6 ? 8'h38 : _GEN_1542; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1544 = 8'h8 == io_state_in_6 ? 8'hbf : _GEN_1543; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1545 = 8'h9 == io_state_in_6 ? 8'h40 : _GEN_1544; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1546 = 8'ha == io_state_in_6 ? 8'ha3 : _GEN_1545; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1547 = 8'hb == io_state_in_6 ? 8'h9e : _GEN_1546; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1548 = 8'hc == io_state_in_6 ? 8'h81 : _GEN_1547; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1549 = 8'hd == io_state_in_6 ? 8'hf3 : _GEN_1548; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1550 = 8'he == io_state_in_6 ? 8'hd7 : _GEN_1549; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1551 = 8'hf == io_state_in_6 ? 8'hfb : _GEN_1550; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1552 = 8'h10 == io_state_in_6 ? 8'h7c : _GEN_1551; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1553 = 8'h11 == io_state_in_6 ? 8'he3 : _GEN_1552; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1554 = 8'h12 == io_state_in_6 ? 8'h39 : _GEN_1553; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1555 = 8'h13 == io_state_in_6 ? 8'h82 : _GEN_1554; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1556 = 8'h14 == io_state_in_6 ? 8'h9b : _GEN_1555; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1557 = 8'h15 == io_state_in_6 ? 8'h2f : _GEN_1556; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1558 = 8'h16 == io_state_in_6 ? 8'hff : _GEN_1557; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1559 = 8'h17 == io_state_in_6 ? 8'h87 : _GEN_1558; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1560 = 8'h18 == io_state_in_6 ? 8'h34 : _GEN_1559; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1561 = 8'h19 == io_state_in_6 ? 8'h8e : _GEN_1560; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1562 = 8'h1a == io_state_in_6 ? 8'h43 : _GEN_1561; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1563 = 8'h1b == io_state_in_6 ? 8'h44 : _GEN_1562; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1564 = 8'h1c == io_state_in_6 ? 8'hc4 : _GEN_1563; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1565 = 8'h1d == io_state_in_6 ? 8'hde : _GEN_1564; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1566 = 8'h1e == io_state_in_6 ? 8'he9 : _GEN_1565; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1567 = 8'h1f == io_state_in_6 ? 8'hcb : _GEN_1566; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1568 = 8'h20 == io_state_in_6 ? 8'h54 : _GEN_1567; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1569 = 8'h21 == io_state_in_6 ? 8'h7b : _GEN_1568; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1570 = 8'h22 == io_state_in_6 ? 8'h94 : _GEN_1569; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1571 = 8'h23 == io_state_in_6 ? 8'h32 : _GEN_1570; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1572 = 8'h24 == io_state_in_6 ? 8'ha6 : _GEN_1571; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1573 = 8'h25 == io_state_in_6 ? 8'hc2 : _GEN_1572; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1574 = 8'h26 == io_state_in_6 ? 8'h23 : _GEN_1573; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1575 = 8'h27 == io_state_in_6 ? 8'h3d : _GEN_1574; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1576 = 8'h28 == io_state_in_6 ? 8'hee : _GEN_1575; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1577 = 8'h29 == io_state_in_6 ? 8'h4c : _GEN_1576; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1578 = 8'h2a == io_state_in_6 ? 8'h95 : _GEN_1577; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1579 = 8'h2b == io_state_in_6 ? 8'hb : _GEN_1578; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1580 = 8'h2c == io_state_in_6 ? 8'h42 : _GEN_1579; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1581 = 8'h2d == io_state_in_6 ? 8'hfa : _GEN_1580; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1582 = 8'h2e == io_state_in_6 ? 8'hc3 : _GEN_1581; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1583 = 8'h2f == io_state_in_6 ? 8'h4e : _GEN_1582; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1584 = 8'h30 == io_state_in_6 ? 8'h8 : _GEN_1583; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1585 = 8'h31 == io_state_in_6 ? 8'h2e : _GEN_1584; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1586 = 8'h32 == io_state_in_6 ? 8'ha1 : _GEN_1585; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1587 = 8'h33 == io_state_in_6 ? 8'h66 : _GEN_1586; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1588 = 8'h34 == io_state_in_6 ? 8'h28 : _GEN_1587; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1589 = 8'h35 == io_state_in_6 ? 8'hd9 : _GEN_1588; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1590 = 8'h36 == io_state_in_6 ? 8'h24 : _GEN_1589; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1591 = 8'h37 == io_state_in_6 ? 8'hb2 : _GEN_1590; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1592 = 8'h38 == io_state_in_6 ? 8'h76 : _GEN_1591; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1593 = 8'h39 == io_state_in_6 ? 8'h5b : _GEN_1592; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1594 = 8'h3a == io_state_in_6 ? 8'ha2 : _GEN_1593; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1595 = 8'h3b == io_state_in_6 ? 8'h49 : _GEN_1594; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1596 = 8'h3c == io_state_in_6 ? 8'h6d : _GEN_1595; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1597 = 8'h3d == io_state_in_6 ? 8'h8b : _GEN_1596; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1598 = 8'h3e == io_state_in_6 ? 8'hd1 : _GEN_1597; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1599 = 8'h3f == io_state_in_6 ? 8'h25 : _GEN_1598; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1600 = 8'h40 == io_state_in_6 ? 8'h72 : _GEN_1599; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1601 = 8'h41 == io_state_in_6 ? 8'hf8 : _GEN_1600; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1602 = 8'h42 == io_state_in_6 ? 8'hf6 : _GEN_1601; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1603 = 8'h43 == io_state_in_6 ? 8'h64 : _GEN_1602; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1604 = 8'h44 == io_state_in_6 ? 8'h86 : _GEN_1603; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1605 = 8'h45 == io_state_in_6 ? 8'h68 : _GEN_1604; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1606 = 8'h46 == io_state_in_6 ? 8'h98 : _GEN_1605; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1607 = 8'h47 == io_state_in_6 ? 8'h16 : _GEN_1606; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1608 = 8'h48 == io_state_in_6 ? 8'hd4 : _GEN_1607; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1609 = 8'h49 == io_state_in_6 ? 8'ha4 : _GEN_1608; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1610 = 8'h4a == io_state_in_6 ? 8'h5c : _GEN_1609; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1611 = 8'h4b == io_state_in_6 ? 8'hcc : _GEN_1610; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1612 = 8'h4c == io_state_in_6 ? 8'h5d : _GEN_1611; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1613 = 8'h4d == io_state_in_6 ? 8'h65 : _GEN_1612; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1614 = 8'h4e == io_state_in_6 ? 8'hb6 : _GEN_1613; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1615 = 8'h4f == io_state_in_6 ? 8'h92 : _GEN_1614; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1616 = 8'h50 == io_state_in_6 ? 8'h6c : _GEN_1615; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1617 = 8'h51 == io_state_in_6 ? 8'h70 : _GEN_1616; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1618 = 8'h52 == io_state_in_6 ? 8'h48 : _GEN_1617; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1619 = 8'h53 == io_state_in_6 ? 8'h50 : _GEN_1618; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1620 = 8'h54 == io_state_in_6 ? 8'hfd : _GEN_1619; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1621 = 8'h55 == io_state_in_6 ? 8'hed : _GEN_1620; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1622 = 8'h56 == io_state_in_6 ? 8'hb9 : _GEN_1621; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1623 = 8'h57 == io_state_in_6 ? 8'hda : _GEN_1622; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1624 = 8'h58 == io_state_in_6 ? 8'h5e : _GEN_1623; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1625 = 8'h59 == io_state_in_6 ? 8'h15 : _GEN_1624; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1626 = 8'h5a == io_state_in_6 ? 8'h46 : _GEN_1625; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1627 = 8'h5b == io_state_in_6 ? 8'h57 : _GEN_1626; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1628 = 8'h5c == io_state_in_6 ? 8'ha7 : _GEN_1627; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1629 = 8'h5d == io_state_in_6 ? 8'h8d : _GEN_1628; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1630 = 8'h5e == io_state_in_6 ? 8'h9d : _GEN_1629; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1631 = 8'h5f == io_state_in_6 ? 8'h84 : _GEN_1630; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1632 = 8'h60 == io_state_in_6 ? 8'h90 : _GEN_1631; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1633 = 8'h61 == io_state_in_6 ? 8'hd8 : _GEN_1632; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1634 = 8'h62 == io_state_in_6 ? 8'hab : _GEN_1633; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1635 = 8'h63 == io_state_in_6 ? 8'h0 : _GEN_1634; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1636 = 8'h64 == io_state_in_6 ? 8'h8c : _GEN_1635; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1637 = 8'h65 == io_state_in_6 ? 8'hbc : _GEN_1636; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1638 = 8'h66 == io_state_in_6 ? 8'hd3 : _GEN_1637; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1639 = 8'h67 == io_state_in_6 ? 8'ha : _GEN_1638; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1640 = 8'h68 == io_state_in_6 ? 8'hf7 : _GEN_1639; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1641 = 8'h69 == io_state_in_6 ? 8'he4 : _GEN_1640; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1642 = 8'h6a == io_state_in_6 ? 8'h58 : _GEN_1641; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1643 = 8'h6b == io_state_in_6 ? 8'h5 : _GEN_1642; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1644 = 8'h6c == io_state_in_6 ? 8'hb8 : _GEN_1643; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1645 = 8'h6d == io_state_in_6 ? 8'hb3 : _GEN_1644; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1646 = 8'h6e == io_state_in_6 ? 8'h45 : _GEN_1645; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1647 = 8'h6f == io_state_in_6 ? 8'h6 : _GEN_1646; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1648 = 8'h70 == io_state_in_6 ? 8'hd0 : _GEN_1647; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1649 = 8'h71 == io_state_in_6 ? 8'h2c : _GEN_1648; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1650 = 8'h72 == io_state_in_6 ? 8'h1e : _GEN_1649; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1651 = 8'h73 == io_state_in_6 ? 8'h8f : _GEN_1650; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1652 = 8'h74 == io_state_in_6 ? 8'hca : _GEN_1651; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1653 = 8'h75 == io_state_in_6 ? 8'h3f : _GEN_1652; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1654 = 8'h76 == io_state_in_6 ? 8'hf : _GEN_1653; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1655 = 8'h77 == io_state_in_6 ? 8'h2 : _GEN_1654; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1656 = 8'h78 == io_state_in_6 ? 8'hc1 : _GEN_1655; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1657 = 8'h79 == io_state_in_6 ? 8'haf : _GEN_1656; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1658 = 8'h7a == io_state_in_6 ? 8'hbd : _GEN_1657; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1659 = 8'h7b == io_state_in_6 ? 8'h3 : _GEN_1658; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1660 = 8'h7c == io_state_in_6 ? 8'h1 : _GEN_1659; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1661 = 8'h7d == io_state_in_6 ? 8'h13 : _GEN_1660; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1662 = 8'h7e == io_state_in_6 ? 8'h8a : _GEN_1661; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1663 = 8'h7f == io_state_in_6 ? 8'h6b : _GEN_1662; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1664 = 8'h80 == io_state_in_6 ? 8'h3a : _GEN_1663; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1665 = 8'h81 == io_state_in_6 ? 8'h91 : _GEN_1664; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1666 = 8'h82 == io_state_in_6 ? 8'h11 : _GEN_1665; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1667 = 8'h83 == io_state_in_6 ? 8'h41 : _GEN_1666; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1668 = 8'h84 == io_state_in_6 ? 8'h4f : _GEN_1667; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1669 = 8'h85 == io_state_in_6 ? 8'h67 : _GEN_1668; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1670 = 8'h86 == io_state_in_6 ? 8'hdc : _GEN_1669; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1671 = 8'h87 == io_state_in_6 ? 8'hea : _GEN_1670; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1672 = 8'h88 == io_state_in_6 ? 8'h97 : _GEN_1671; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1673 = 8'h89 == io_state_in_6 ? 8'hf2 : _GEN_1672; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1674 = 8'h8a == io_state_in_6 ? 8'hcf : _GEN_1673; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1675 = 8'h8b == io_state_in_6 ? 8'hce : _GEN_1674; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1676 = 8'h8c == io_state_in_6 ? 8'hf0 : _GEN_1675; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1677 = 8'h8d == io_state_in_6 ? 8'hb4 : _GEN_1676; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1678 = 8'h8e == io_state_in_6 ? 8'he6 : _GEN_1677; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1679 = 8'h8f == io_state_in_6 ? 8'h73 : _GEN_1678; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1680 = 8'h90 == io_state_in_6 ? 8'h96 : _GEN_1679; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1681 = 8'h91 == io_state_in_6 ? 8'hac : _GEN_1680; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1682 = 8'h92 == io_state_in_6 ? 8'h74 : _GEN_1681; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1683 = 8'h93 == io_state_in_6 ? 8'h22 : _GEN_1682; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1684 = 8'h94 == io_state_in_6 ? 8'he7 : _GEN_1683; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1685 = 8'h95 == io_state_in_6 ? 8'had : _GEN_1684; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1686 = 8'h96 == io_state_in_6 ? 8'h35 : _GEN_1685; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1687 = 8'h97 == io_state_in_6 ? 8'h85 : _GEN_1686; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1688 = 8'h98 == io_state_in_6 ? 8'he2 : _GEN_1687; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1689 = 8'h99 == io_state_in_6 ? 8'hf9 : _GEN_1688; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1690 = 8'h9a == io_state_in_6 ? 8'h37 : _GEN_1689; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1691 = 8'h9b == io_state_in_6 ? 8'he8 : _GEN_1690; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1692 = 8'h9c == io_state_in_6 ? 8'h1c : _GEN_1691; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1693 = 8'h9d == io_state_in_6 ? 8'h75 : _GEN_1692; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1694 = 8'h9e == io_state_in_6 ? 8'hdf : _GEN_1693; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1695 = 8'h9f == io_state_in_6 ? 8'h6e : _GEN_1694; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1696 = 8'ha0 == io_state_in_6 ? 8'h47 : _GEN_1695; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1697 = 8'ha1 == io_state_in_6 ? 8'hf1 : _GEN_1696; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1698 = 8'ha2 == io_state_in_6 ? 8'h1a : _GEN_1697; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1699 = 8'ha3 == io_state_in_6 ? 8'h71 : _GEN_1698; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1700 = 8'ha4 == io_state_in_6 ? 8'h1d : _GEN_1699; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1701 = 8'ha5 == io_state_in_6 ? 8'h29 : _GEN_1700; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1702 = 8'ha6 == io_state_in_6 ? 8'hc5 : _GEN_1701; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1703 = 8'ha7 == io_state_in_6 ? 8'h89 : _GEN_1702; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1704 = 8'ha8 == io_state_in_6 ? 8'h6f : _GEN_1703; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1705 = 8'ha9 == io_state_in_6 ? 8'hb7 : _GEN_1704; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1706 = 8'haa == io_state_in_6 ? 8'h62 : _GEN_1705; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1707 = 8'hab == io_state_in_6 ? 8'he : _GEN_1706; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1708 = 8'hac == io_state_in_6 ? 8'haa : _GEN_1707; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1709 = 8'had == io_state_in_6 ? 8'h18 : _GEN_1708; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1710 = 8'hae == io_state_in_6 ? 8'hbe : _GEN_1709; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1711 = 8'haf == io_state_in_6 ? 8'h1b : _GEN_1710; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1712 = 8'hb0 == io_state_in_6 ? 8'hfc : _GEN_1711; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1713 = 8'hb1 == io_state_in_6 ? 8'h56 : _GEN_1712; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1714 = 8'hb2 == io_state_in_6 ? 8'h3e : _GEN_1713; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1715 = 8'hb3 == io_state_in_6 ? 8'h4b : _GEN_1714; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1716 = 8'hb4 == io_state_in_6 ? 8'hc6 : _GEN_1715; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1717 = 8'hb5 == io_state_in_6 ? 8'hd2 : _GEN_1716; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1718 = 8'hb6 == io_state_in_6 ? 8'h79 : _GEN_1717; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1719 = 8'hb7 == io_state_in_6 ? 8'h20 : _GEN_1718; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1720 = 8'hb8 == io_state_in_6 ? 8'h9a : _GEN_1719; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1721 = 8'hb9 == io_state_in_6 ? 8'hdb : _GEN_1720; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1722 = 8'hba == io_state_in_6 ? 8'hc0 : _GEN_1721; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1723 = 8'hbb == io_state_in_6 ? 8'hfe : _GEN_1722; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1724 = 8'hbc == io_state_in_6 ? 8'h78 : _GEN_1723; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1725 = 8'hbd == io_state_in_6 ? 8'hcd : _GEN_1724; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1726 = 8'hbe == io_state_in_6 ? 8'h5a : _GEN_1725; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1727 = 8'hbf == io_state_in_6 ? 8'hf4 : _GEN_1726; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1728 = 8'hc0 == io_state_in_6 ? 8'h1f : _GEN_1727; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1729 = 8'hc1 == io_state_in_6 ? 8'hdd : _GEN_1728; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1730 = 8'hc2 == io_state_in_6 ? 8'ha8 : _GEN_1729; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1731 = 8'hc3 == io_state_in_6 ? 8'h33 : _GEN_1730; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1732 = 8'hc4 == io_state_in_6 ? 8'h88 : _GEN_1731; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1733 = 8'hc5 == io_state_in_6 ? 8'h7 : _GEN_1732; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1734 = 8'hc6 == io_state_in_6 ? 8'hc7 : _GEN_1733; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1735 = 8'hc7 == io_state_in_6 ? 8'h31 : _GEN_1734; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1736 = 8'hc8 == io_state_in_6 ? 8'hb1 : _GEN_1735; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1737 = 8'hc9 == io_state_in_6 ? 8'h12 : _GEN_1736; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1738 = 8'hca == io_state_in_6 ? 8'h10 : _GEN_1737; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1739 = 8'hcb == io_state_in_6 ? 8'h59 : _GEN_1738; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1740 = 8'hcc == io_state_in_6 ? 8'h27 : _GEN_1739; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1741 = 8'hcd == io_state_in_6 ? 8'h80 : _GEN_1740; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1742 = 8'hce == io_state_in_6 ? 8'hec : _GEN_1741; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1743 = 8'hcf == io_state_in_6 ? 8'h5f : _GEN_1742; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1744 = 8'hd0 == io_state_in_6 ? 8'h60 : _GEN_1743; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1745 = 8'hd1 == io_state_in_6 ? 8'h51 : _GEN_1744; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1746 = 8'hd2 == io_state_in_6 ? 8'h7f : _GEN_1745; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1747 = 8'hd3 == io_state_in_6 ? 8'ha9 : _GEN_1746; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1748 = 8'hd4 == io_state_in_6 ? 8'h19 : _GEN_1747; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1749 = 8'hd5 == io_state_in_6 ? 8'hb5 : _GEN_1748; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1750 = 8'hd6 == io_state_in_6 ? 8'h4a : _GEN_1749; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1751 = 8'hd7 == io_state_in_6 ? 8'hd : _GEN_1750; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1752 = 8'hd8 == io_state_in_6 ? 8'h2d : _GEN_1751; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1753 = 8'hd9 == io_state_in_6 ? 8'he5 : _GEN_1752; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1754 = 8'hda == io_state_in_6 ? 8'h7a : _GEN_1753; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1755 = 8'hdb == io_state_in_6 ? 8'h9f : _GEN_1754; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1756 = 8'hdc == io_state_in_6 ? 8'h93 : _GEN_1755; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1757 = 8'hdd == io_state_in_6 ? 8'hc9 : _GEN_1756; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1758 = 8'hde == io_state_in_6 ? 8'h9c : _GEN_1757; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1759 = 8'hdf == io_state_in_6 ? 8'hef : _GEN_1758; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1760 = 8'he0 == io_state_in_6 ? 8'ha0 : _GEN_1759; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1761 = 8'he1 == io_state_in_6 ? 8'he0 : _GEN_1760; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1762 = 8'he2 == io_state_in_6 ? 8'h3b : _GEN_1761; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1763 = 8'he3 == io_state_in_6 ? 8'h4d : _GEN_1762; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1764 = 8'he4 == io_state_in_6 ? 8'hae : _GEN_1763; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1765 = 8'he5 == io_state_in_6 ? 8'h2a : _GEN_1764; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1766 = 8'he6 == io_state_in_6 ? 8'hf5 : _GEN_1765; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1767 = 8'he7 == io_state_in_6 ? 8'hb0 : _GEN_1766; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1768 = 8'he8 == io_state_in_6 ? 8'hc8 : _GEN_1767; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1769 = 8'he9 == io_state_in_6 ? 8'heb : _GEN_1768; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1770 = 8'hea == io_state_in_6 ? 8'hbb : _GEN_1769; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1771 = 8'heb == io_state_in_6 ? 8'h3c : _GEN_1770; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1772 = 8'hec == io_state_in_6 ? 8'h83 : _GEN_1771; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1773 = 8'hed == io_state_in_6 ? 8'h53 : _GEN_1772; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1774 = 8'hee == io_state_in_6 ? 8'h99 : _GEN_1773; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1775 = 8'hef == io_state_in_6 ? 8'h61 : _GEN_1774; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1776 = 8'hf0 == io_state_in_6 ? 8'h17 : _GEN_1775; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1777 = 8'hf1 == io_state_in_6 ? 8'h2b : _GEN_1776; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1778 = 8'hf2 == io_state_in_6 ? 8'h4 : _GEN_1777; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1779 = 8'hf3 == io_state_in_6 ? 8'h7e : _GEN_1778; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1780 = 8'hf4 == io_state_in_6 ? 8'hba : _GEN_1779; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1781 = 8'hf5 == io_state_in_6 ? 8'h77 : _GEN_1780; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1782 = 8'hf6 == io_state_in_6 ? 8'hd6 : _GEN_1781; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1783 = 8'hf7 == io_state_in_6 ? 8'h26 : _GEN_1782; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1784 = 8'hf8 == io_state_in_6 ? 8'he1 : _GEN_1783; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1785 = 8'hf9 == io_state_in_6 ? 8'h69 : _GEN_1784; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1786 = 8'hfa == io_state_in_6 ? 8'h14 : _GEN_1785; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1787 = 8'hfb == io_state_in_6 ? 8'h63 : _GEN_1786; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1788 = 8'hfc == io_state_in_6 ? 8'h55 : _GEN_1787; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1789 = 8'hfd == io_state_in_6 ? 8'h21 : _GEN_1788; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1790 = 8'hfe == io_state_in_6 ? 8'hc : _GEN_1789; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1793 = 8'h1 == io_state_in_7 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1794 = 8'h2 == io_state_in_7 ? 8'h6a : _GEN_1793; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1795 = 8'h3 == io_state_in_7 ? 8'hd5 : _GEN_1794; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1796 = 8'h4 == io_state_in_7 ? 8'h30 : _GEN_1795; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1797 = 8'h5 == io_state_in_7 ? 8'h36 : _GEN_1796; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1798 = 8'h6 == io_state_in_7 ? 8'ha5 : _GEN_1797; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1799 = 8'h7 == io_state_in_7 ? 8'h38 : _GEN_1798; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1800 = 8'h8 == io_state_in_7 ? 8'hbf : _GEN_1799; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1801 = 8'h9 == io_state_in_7 ? 8'h40 : _GEN_1800; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1802 = 8'ha == io_state_in_7 ? 8'ha3 : _GEN_1801; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1803 = 8'hb == io_state_in_7 ? 8'h9e : _GEN_1802; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1804 = 8'hc == io_state_in_7 ? 8'h81 : _GEN_1803; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1805 = 8'hd == io_state_in_7 ? 8'hf3 : _GEN_1804; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1806 = 8'he == io_state_in_7 ? 8'hd7 : _GEN_1805; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1807 = 8'hf == io_state_in_7 ? 8'hfb : _GEN_1806; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1808 = 8'h10 == io_state_in_7 ? 8'h7c : _GEN_1807; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1809 = 8'h11 == io_state_in_7 ? 8'he3 : _GEN_1808; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1810 = 8'h12 == io_state_in_7 ? 8'h39 : _GEN_1809; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1811 = 8'h13 == io_state_in_7 ? 8'h82 : _GEN_1810; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1812 = 8'h14 == io_state_in_7 ? 8'h9b : _GEN_1811; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1813 = 8'h15 == io_state_in_7 ? 8'h2f : _GEN_1812; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1814 = 8'h16 == io_state_in_7 ? 8'hff : _GEN_1813; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1815 = 8'h17 == io_state_in_7 ? 8'h87 : _GEN_1814; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1816 = 8'h18 == io_state_in_7 ? 8'h34 : _GEN_1815; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1817 = 8'h19 == io_state_in_7 ? 8'h8e : _GEN_1816; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1818 = 8'h1a == io_state_in_7 ? 8'h43 : _GEN_1817; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1819 = 8'h1b == io_state_in_7 ? 8'h44 : _GEN_1818; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1820 = 8'h1c == io_state_in_7 ? 8'hc4 : _GEN_1819; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1821 = 8'h1d == io_state_in_7 ? 8'hde : _GEN_1820; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1822 = 8'h1e == io_state_in_7 ? 8'he9 : _GEN_1821; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1823 = 8'h1f == io_state_in_7 ? 8'hcb : _GEN_1822; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1824 = 8'h20 == io_state_in_7 ? 8'h54 : _GEN_1823; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1825 = 8'h21 == io_state_in_7 ? 8'h7b : _GEN_1824; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1826 = 8'h22 == io_state_in_7 ? 8'h94 : _GEN_1825; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1827 = 8'h23 == io_state_in_7 ? 8'h32 : _GEN_1826; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1828 = 8'h24 == io_state_in_7 ? 8'ha6 : _GEN_1827; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1829 = 8'h25 == io_state_in_7 ? 8'hc2 : _GEN_1828; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1830 = 8'h26 == io_state_in_7 ? 8'h23 : _GEN_1829; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1831 = 8'h27 == io_state_in_7 ? 8'h3d : _GEN_1830; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1832 = 8'h28 == io_state_in_7 ? 8'hee : _GEN_1831; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1833 = 8'h29 == io_state_in_7 ? 8'h4c : _GEN_1832; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1834 = 8'h2a == io_state_in_7 ? 8'h95 : _GEN_1833; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1835 = 8'h2b == io_state_in_7 ? 8'hb : _GEN_1834; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1836 = 8'h2c == io_state_in_7 ? 8'h42 : _GEN_1835; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1837 = 8'h2d == io_state_in_7 ? 8'hfa : _GEN_1836; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1838 = 8'h2e == io_state_in_7 ? 8'hc3 : _GEN_1837; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1839 = 8'h2f == io_state_in_7 ? 8'h4e : _GEN_1838; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1840 = 8'h30 == io_state_in_7 ? 8'h8 : _GEN_1839; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1841 = 8'h31 == io_state_in_7 ? 8'h2e : _GEN_1840; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1842 = 8'h32 == io_state_in_7 ? 8'ha1 : _GEN_1841; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1843 = 8'h33 == io_state_in_7 ? 8'h66 : _GEN_1842; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1844 = 8'h34 == io_state_in_7 ? 8'h28 : _GEN_1843; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1845 = 8'h35 == io_state_in_7 ? 8'hd9 : _GEN_1844; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1846 = 8'h36 == io_state_in_7 ? 8'h24 : _GEN_1845; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1847 = 8'h37 == io_state_in_7 ? 8'hb2 : _GEN_1846; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1848 = 8'h38 == io_state_in_7 ? 8'h76 : _GEN_1847; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1849 = 8'h39 == io_state_in_7 ? 8'h5b : _GEN_1848; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1850 = 8'h3a == io_state_in_7 ? 8'ha2 : _GEN_1849; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1851 = 8'h3b == io_state_in_7 ? 8'h49 : _GEN_1850; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1852 = 8'h3c == io_state_in_7 ? 8'h6d : _GEN_1851; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1853 = 8'h3d == io_state_in_7 ? 8'h8b : _GEN_1852; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1854 = 8'h3e == io_state_in_7 ? 8'hd1 : _GEN_1853; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1855 = 8'h3f == io_state_in_7 ? 8'h25 : _GEN_1854; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1856 = 8'h40 == io_state_in_7 ? 8'h72 : _GEN_1855; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1857 = 8'h41 == io_state_in_7 ? 8'hf8 : _GEN_1856; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1858 = 8'h42 == io_state_in_7 ? 8'hf6 : _GEN_1857; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1859 = 8'h43 == io_state_in_7 ? 8'h64 : _GEN_1858; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1860 = 8'h44 == io_state_in_7 ? 8'h86 : _GEN_1859; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1861 = 8'h45 == io_state_in_7 ? 8'h68 : _GEN_1860; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1862 = 8'h46 == io_state_in_7 ? 8'h98 : _GEN_1861; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1863 = 8'h47 == io_state_in_7 ? 8'h16 : _GEN_1862; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1864 = 8'h48 == io_state_in_7 ? 8'hd4 : _GEN_1863; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1865 = 8'h49 == io_state_in_7 ? 8'ha4 : _GEN_1864; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1866 = 8'h4a == io_state_in_7 ? 8'h5c : _GEN_1865; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1867 = 8'h4b == io_state_in_7 ? 8'hcc : _GEN_1866; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1868 = 8'h4c == io_state_in_7 ? 8'h5d : _GEN_1867; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1869 = 8'h4d == io_state_in_7 ? 8'h65 : _GEN_1868; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1870 = 8'h4e == io_state_in_7 ? 8'hb6 : _GEN_1869; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1871 = 8'h4f == io_state_in_7 ? 8'h92 : _GEN_1870; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1872 = 8'h50 == io_state_in_7 ? 8'h6c : _GEN_1871; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1873 = 8'h51 == io_state_in_7 ? 8'h70 : _GEN_1872; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1874 = 8'h52 == io_state_in_7 ? 8'h48 : _GEN_1873; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1875 = 8'h53 == io_state_in_7 ? 8'h50 : _GEN_1874; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1876 = 8'h54 == io_state_in_7 ? 8'hfd : _GEN_1875; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1877 = 8'h55 == io_state_in_7 ? 8'hed : _GEN_1876; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1878 = 8'h56 == io_state_in_7 ? 8'hb9 : _GEN_1877; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1879 = 8'h57 == io_state_in_7 ? 8'hda : _GEN_1878; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1880 = 8'h58 == io_state_in_7 ? 8'h5e : _GEN_1879; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1881 = 8'h59 == io_state_in_7 ? 8'h15 : _GEN_1880; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1882 = 8'h5a == io_state_in_7 ? 8'h46 : _GEN_1881; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1883 = 8'h5b == io_state_in_7 ? 8'h57 : _GEN_1882; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1884 = 8'h5c == io_state_in_7 ? 8'ha7 : _GEN_1883; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1885 = 8'h5d == io_state_in_7 ? 8'h8d : _GEN_1884; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1886 = 8'h5e == io_state_in_7 ? 8'h9d : _GEN_1885; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1887 = 8'h5f == io_state_in_7 ? 8'h84 : _GEN_1886; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1888 = 8'h60 == io_state_in_7 ? 8'h90 : _GEN_1887; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1889 = 8'h61 == io_state_in_7 ? 8'hd8 : _GEN_1888; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1890 = 8'h62 == io_state_in_7 ? 8'hab : _GEN_1889; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1891 = 8'h63 == io_state_in_7 ? 8'h0 : _GEN_1890; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1892 = 8'h64 == io_state_in_7 ? 8'h8c : _GEN_1891; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1893 = 8'h65 == io_state_in_7 ? 8'hbc : _GEN_1892; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1894 = 8'h66 == io_state_in_7 ? 8'hd3 : _GEN_1893; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1895 = 8'h67 == io_state_in_7 ? 8'ha : _GEN_1894; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1896 = 8'h68 == io_state_in_7 ? 8'hf7 : _GEN_1895; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1897 = 8'h69 == io_state_in_7 ? 8'he4 : _GEN_1896; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1898 = 8'h6a == io_state_in_7 ? 8'h58 : _GEN_1897; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1899 = 8'h6b == io_state_in_7 ? 8'h5 : _GEN_1898; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1900 = 8'h6c == io_state_in_7 ? 8'hb8 : _GEN_1899; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1901 = 8'h6d == io_state_in_7 ? 8'hb3 : _GEN_1900; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1902 = 8'h6e == io_state_in_7 ? 8'h45 : _GEN_1901; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1903 = 8'h6f == io_state_in_7 ? 8'h6 : _GEN_1902; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1904 = 8'h70 == io_state_in_7 ? 8'hd0 : _GEN_1903; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1905 = 8'h71 == io_state_in_7 ? 8'h2c : _GEN_1904; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1906 = 8'h72 == io_state_in_7 ? 8'h1e : _GEN_1905; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1907 = 8'h73 == io_state_in_7 ? 8'h8f : _GEN_1906; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1908 = 8'h74 == io_state_in_7 ? 8'hca : _GEN_1907; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1909 = 8'h75 == io_state_in_7 ? 8'h3f : _GEN_1908; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1910 = 8'h76 == io_state_in_7 ? 8'hf : _GEN_1909; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1911 = 8'h77 == io_state_in_7 ? 8'h2 : _GEN_1910; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1912 = 8'h78 == io_state_in_7 ? 8'hc1 : _GEN_1911; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1913 = 8'h79 == io_state_in_7 ? 8'haf : _GEN_1912; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1914 = 8'h7a == io_state_in_7 ? 8'hbd : _GEN_1913; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1915 = 8'h7b == io_state_in_7 ? 8'h3 : _GEN_1914; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1916 = 8'h7c == io_state_in_7 ? 8'h1 : _GEN_1915; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1917 = 8'h7d == io_state_in_7 ? 8'h13 : _GEN_1916; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1918 = 8'h7e == io_state_in_7 ? 8'h8a : _GEN_1917; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1919 = 8'h7f == io_state_in_7 ? 8'h6b : _GEN_1918; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1920 = 8'h80 == io_state_in_7 ? 8'h3a : _GEN_1919; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1921 = 8'h81 == io_state_in_7 ? 8'h91 : _GEN_1920; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1922 = 8'h82 == io_state_in_7 ? 8'h11 : _GEN_1921; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1923 = 8'h83 == io_state_in_7 ? 8'h41 : _GEN_1922; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1924 = 8'h84 == io_state_in_7 ? 8'h4f : _GEN_1923; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1925 = 8'h85 == io_state_in_7 ? 8'h67 : _GEN_1924; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1926 = 8'h86 == io_state_in_7 ? 8'hdc : _GEN_1925; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1927 = 8'h87 == io_state_in_7 ? 8'hea : _GEN_1926; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1928 = 8'h88 == io_state_in_7 ? 8'h97 : _GEN_1927; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1929 = 8'h89 == io_state_in_7 ? 8'hf2 : _GEN_1928; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1930 = 8'h8a == io_state_in_7 ? 8'hcf : _GEN_1929; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1931 = 8'h8b == io_state_in_7 ? 8'hce : _GEN_1930; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1932 = 8'h8c == io_state_in_7 ? 8'hf0 : _GEN_1931; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1933 = 8'h8d == io_state_in_7 ? 8'hb4 : _GEN_1932; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1934 = 8'h8e == io_state_in_7 ? 8'he6 : _GEN_1933; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1935 = 8'h8f == io_state_in_7 ? 8'h73 : _GEN_1934; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1936 = 8'h90 == io_state_in_7 ? 8'h96 : _GEN_1935; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1937 = 8'h91 == io_state_in_7 ? 8'hac : _GEN_1936; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1938 = 8'h92 == io_state_in_7 ? 8'h74 : _GEN_1937; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1939 = 8'h93 == io_state_in_7 ? 8'h22 : _GEN_1938; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1940 = 8'h94 == io_state_in_7 ? 8'he7 : _GEN_1939; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1941 = 8'h95 == io_state_in_7 ? 8'had : _GEN_1940; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1942 = 8'h96 == io_state_in_7 ? 8'h35 : _GEN_1941; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1943 = 8'h97 == io_state_in_7 ? 8'h85 : _GEN_1942; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1944 = 8'h98 == io_state_in_7 ? 8'he2 : _GEN_1943; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1945 = 8'h99 == io_state_in_7 ? 8'hf9 : _GEN_1944; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1946 = 8'h9a == io_state_in_7 ? 8'h37 : _GEN_1945; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1947 = 8'h9b == io_state_in_7 ? 8'he8 : _GEN_1946; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1948 = 8'h9c == io_state_in_7 ? 8'h1c : _GEN_1947; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1949 = 8'h9d == io_state_in_7 ? 8'h75 : _GEN_1948; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1950 = 8'h9e == io_state_in_7 ? 8'hdf : _GEN_1949; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1951 = 8'h9f == io_state_in_7 ? 8'h6e : _GEN_1950; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1952 = 8'ha0 == io_state_in_7 ? 8'h47 : _GEN_1951; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1953 = 8'ha1 == io_state_in_7 ? 8'hf1 : _GEN_1952; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1954 = 8'ha2 == io_state_in_7 ? 8'h1a : _GEN_1953; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1955 = 8'ha3 == io_state_in_7 ? 8'h71 : _GEN_1954; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1956 = 8'ha4 == io_state_in_7 ? 8'h1d : _GEN_1955; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1957 = 8'ha5 == io_state_in_7 ? 8'h29 : _GEN_1956; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1958 = 8'ha6 == io_state_in_7 ? 8'hc5 : _GEN_1957; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1959 = 8'ha7 == io_state_in_7 ? 8'h89 : _GEN_1958; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1960 = 8'ha8 == io_state_in_7 ? 8'h6f : _GEN_1959; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1961 = 8'ha9 == io_state_in_7 ? 8'hb7 : _GEN_1960; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1962 = 8'haa == io_state_in_7 ? 8'h62 : _GEN_1961; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1963 = 8'hab == io_state_in_7 ? 8'he : _GEN_1962; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1964 = 8'hac == io_state_in_7 ? 8'haa : _GEN_1963; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1965 = 8'had == io_state_in_7 ? 8'h18 : _GEN_1964; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1966 = 8'hae == io_state_in_7 ? 8'hbe : _GEN_1965; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1967 = 8'haf == io_state_in_7 ? 8'h1b : _GEN_1966; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1968 = 8'hb0 == io_state_in_7 ? 8'hfc : _GEN_1967; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1969 = 8'hb1 == io_state_in_7 ? 8'h56 : _GEN_1968; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1970 = 8'hb2 == io_state_in_7 ? 8'h3e : _GEN_1969; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1971 = 8'hb3 == io_state_in_7 ? 8'h4b : _GEN_1970; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1972 = 8'hb4 == io_state_in_7 ? 8'hc6 : _GEN_1971; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1973 = 8'hb5 == io_state_in_7 ? 8'hd2 : _GEN_1972; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1974 = 8'hb6 == io_state_in_7 ? 8'h79 : _GEN_1973; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1975 = 8'hb7 == io_state_in_7 ? 8'h20 : _GEN_1974; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1976 = 8'hb8 == io_state_in_7 ? 8'h9a : _GEN_1975; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1977 = 8'hb9 == io_state_in_7 ? 8'hdb : _GEN_1976; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1978 = 8'hba == io_state_in_7 ? 8'hc0 : _GEN_1977; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1979 = 8'hbb == io_state_in_7 ? 8'hfe : _GEN_1978; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1980 = 8'hbc == io_state_in_7 ? 8'h78 : _GEN_1979; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1981 = 8'hbd == io_state_in_7 ? 8'hcd : _GEN_1980; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1982 = 8'hbe == io_state_in_7 ? 8'h5a : _GEN_1981; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1983 = 8'hbf == io_state_in_7 ? 8'hf4 : _GEN_1982; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1984 = 8'hc0 == io_state_in_7 ? 8'h1f : _GEN_1983; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1985 = 8'hc1 == io_state_in_7 ? 8'hdd : _GEN_1984; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1986 = 8'hc2 == io_state_in_7 ? 8'ha8 : _GEN_1985; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1987 = 8'hc3 == io_state_in_7 ? 8'h33 : _GEN_1986; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1988 = 8'hc4 == io_state_in_7 ? 8'h88 : _GEN_1987; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1989 = 8'hc5 == io_state_in_7 ? 8'h7 : _GEN_1988; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1990 = 8'hc6 == io_state_in_7 ? 8'hc7 : _GEN_1989; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1991 = 8'hc7 == io_state_in_7 ? 8'h31 : _GEN_1990; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1992 = 8'hc8 == io_state_in_7 ? 8'hb1 : _GEN_1991; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1993 = 8'hc9 == io_state_in_7 ? 8'h12 : _GEN_1992; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1994 = 8'hca == io_state_in_7 ? 8'h10 : _GEN_1993; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1995 = 8'hcb == io_state_in_7 ? 8'h59 : _GEN_1994; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1996 = 8'hcc == io_state_in_7 ? 8'h27 : _GEN_1995; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1997 = 8'hcd == io_state_in_7 ? 8'h80 : _GEN_1996; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1998 = 8'hce == io_state_in_7 ? 8'hec : _GEN_1997; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_1999 = 8'hcf == io_state_in_7 ? 8'h5f : _GEN_1998; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2000 = 8'hd0 == io_state_in_7 ? 8'h60 : _GEN_1999; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2001 = 8'hd1 == io_state_in_7 ? 8'h51 : _GEN_2000; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2002 = 8'hd2 == io_state_in_7 ? 8'h7f : _GEN_2001; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2003 = 8'hd3 == io_state_in_7 ? 8'ha9 : _GEN_2002; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2004 = 8'hd4 == io_state_in_7 ? 8'h19 : _GEN_2003; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2005 = 8'hd5 == io_state_in_7 ? 8'hb5 : _GEN_2004; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2006 = 8'hd6 == io_state_in_7 ? 8'h4a : _GEN_2005; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2007 = 8'hd7 == io_state_in_7 ? 8'hd : _GEN_2006; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2008 = 8'hd8 == io_state_in_7 ? 8'h2d : _GEN_2007; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2009 = 8'hd9 == io_state_in_7 ? 8'he5 : _GEN_2008; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2010 = 8'hda == io_state_in_7 ? 8'h7a : _GEN_2009; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2011 = 8'hdb == io_state_in_7 ? 8'h9f : _GEN_2010; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2012 = 8'hdc == io_state_in_7 ? 8'h93 : _GEN_2011; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2013 = 8'hdd == io_state_in_7 ? 8'hc9 : _GEN_2012; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2014 = 8'hde == io_state_in_7 ? 8'h9c : _GEN_2013; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2015 = 8'hdf == io_state_in_7 ? 8'hef : _GEN_2014; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2016 = 8'he0 == io_state_in_7 ? 8'ha0 : _GEN_2015; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2017 = 8'he1 == io_state_in_7 ? 8'he0 : _GEN_2016; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2018 = 8'he2 == io_state_in_7 ? 8'h3b : _GEN_2017; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2019 = 8'he3 == io_state_in_7 ? 8'h4d : _GEN_2018; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2020 = 8'he4 == io_state_in_7 ? 8'hae : _GEN_2019; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2021 = 8'he5 == io_state_in_7 ? 8'h2a : _GEN_2020; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2022 = 8'he6 == io_state_in_7 ? 8'hf5 : _GEN_2021; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2023 = 8'he7 == io_state_in_7 ? 8'hb0 : _GEN_2022; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2024 = 8'he8 == io_state_in_7 ? 8'hc8 : _GEN_2023; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2025 = 8'he9 == io_state_in_7 ? 8'heb : _GEN_2024; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2026 = 8'hea == io_state_in_7 ? 8'hbb : _GEN_2025; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2027 = 8'heb == io_state_in_7 ? 8'h3c : _GEN_2026; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2028 = 8'hec == io_state_in_7 ? 8'h83 : _GEN_2027; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2029 = 8'hed == io_state_in_7 ? 8'h53 : _GEN_2028; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2030 = 8'hee == io_state_in_7 ? 8'h99 : _GEN_2029; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2031 = 8'hef == io_state_in_7 ? 8'h61 : _GEN_2030; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2032 = 8'hf0 == io_state_in_7 ? 8'h17 : _GEN_2031; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2033 = 8'hf1 == io_state_in_7 ? 8'h2b : _GEN_2032; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2034 = 8'hf2 == io_state_in_7 ? 8'h4 : _GEN_2033; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2035 = 8'hf3 == io_state_in_7 ? 8'h7e : _GEN_2034; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2036 = 8'hf4 == io_state_in_7 ? 8'hba : _GEN_2035; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2037 = 8'hf5 == io_state_in_7 ? 8'h77 : _GEN_2036; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2038 = 8'hf6 == io_state_in_7 ? 8'hd6 : _GEN_2037; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2039 = 8'hf7 == io_state_in_7 ? 8'h26 : _GEN_2038; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2040 = 8'hf8 == io_state_in_7 ? 8'he1 : _GEN_2039; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2041 = 8'hf9 == io_state_in_7 ? 8'h69 : _GEN_2040; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2042 = 8'hfa == io_state_in_7 ? 8'h14 : _GEN_2041; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2043 = 8'hfb == io_state_in_7 ? 8'h63 : _GEN_2042; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2044 = 8'hfc == io_state_in_7 ? 8'h55 : _GEN_2043; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2045 = 8'hfd == io_state_in_7 ? 8'h21 : _GEN_2044; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2046 = 8'hfe == io_state_in_7 ? 8'hc : _GEN_2045; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2049 = 8'h1 == io_state_in_8 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2050 = 8'h2 == io_state_in_8 ? 8'h6a : _GEN_2049; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2051 = 8'h3 == io_state_in_8 ? 8'hd5 : _GEN_2050; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2052 = 8'h4 == io_state_in_8 ? 8'h30 : _GEN_2051; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2053 = 8'h5 == io_state_in_8 ? 8'h36 : _GEN_2052; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2054 = 8'h6 == io_state_in_8 ? 8'ha5 : _GEN_2053; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2055 = 8'h7 == io_state_in_8 ? 8'h38 : _GEN_2054; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2056 = 8'h8 == io_state_in_8 ? 8'hbf : _GEN_2055; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2057 = 8'h9 == io_state_in_8 ? 8'h40 : _GEN_2056; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2058 = 8'ha == io_state_in_8 ? 8'ha3 : _GEN_2057; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2059 = 8'hb == io_state_in_8 ? 8'h9e : _GEN_2058; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2060 = 8'hc == io_state_in_8 ? 8'h81 : _GEN_2059; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2061 = 8'hd == io_state_in_8 ? 8'hf3 : _GEN_2060; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2062 = 8'he == io_state_in_8 ? 8'hd7 : _GEN_2061; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2063 = 8'hf == io_state_in_8 ? 8'hfb : _GEN_2062; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2064 = 8'h10 == io_state_in_8 ? 8'h7c : _GEN_2063; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2065 = 8'h11 == io_state_in_8 ? 8'he3 : _GEN_2064; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2066 = 8'h12 == io_state_in_8 ? 8'h39 : _GEN_2065; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2067 = 8'h13 == io_state_in_8 ? 8'h82 : _GEN_2066; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2068 = 8'h14 == io_state_in_8 ? 8'h9b : _GEN_2067; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2069 = 8'h15 == io_state_in_8 ? 8'h2f : _GEN_2068; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2070 = 8'h16 == io_state_in_8 ? 8'hff : _GEN_2069; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2071 = 8'h17 == io_state_in_8 ? 8'h87 : _GEN_2070; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2072 = 8'h18 == io_state_in_8 ? 8'h34 : _GEN_2071; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2073 = 8'h19 == io_state_in_8 ? 8'h8e : _GEN_2072; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2074 = 8'h1a == io_state_in_8 ? 8'h43 : _GEN_2073; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2075 = 8'h1b == io_state_in_8 ? 8'h44 : _GEN_2074; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2076 = 8'h1c == io_state_in_8 ? 8'hc4 : _GEN_2075; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2077 = 8'h1d == io_state_in_8 ? 8'hde : _GEN_2076; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2078 = 8'h1e == io_state_in_8 ? 8'he9 : _GEN_2077; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2079 = 8'h1f == io_state_in_8 ? 8'hcb : _GEN_2078; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2080 = 8'h20 == io_state_in_8 ? 8'h54 : _GEN_2079; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2081 = 8'h21 == io_state_in_8 ? 8'h7b : _GEN_2080; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2082 = 8'h22 == io_state_in_8 ? 8'h94 : _GEN_2081; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2083 = 8'h23 == io_state_in_8 ? 8'h32 : _GEN_2082; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2084 = 8'h24 == io_state_in_8 ? 8'ha6 : _GEN_2083; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2085 = 8'h25 == io_state_in_8 ? 8'hc2 : _GEN_2084; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2086 = 8'h26 == io_state_in_8 ? 8'h23 : _GEN_2085; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2087 = 8'h27 == io_state_in_8 ? 8'h3d : _GEN_2086; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2088 = 8'h28 == io_state_in_8 ? 8'hee : _GEN_2087; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2089 = 8'h29 == io_state_in_8 ? 8'h4c : _GEN_2088; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2090 = 8'h2a == io_state_in_8 ? 8'h95 : _GEN_2089; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2091 = 8'h2b == io_state_in_8 ? 8'hb : _GEN_2090; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2092 = 8'h2c == io_state_in_8 ? 8'h42 : _GEN_2091; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2093 = 8'h2d == io_state_in_8 ? 8'hfa : _GEN_2092; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2094 = 8'h2e == io_state_in_8 ? 8'hc3 : _GEN_2093; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2095 = 8'h2f == io_state_in_8 ? 8'h4e : _GEN_2094; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2096 = 8'h30 == io_state_in_8 ? 8'h8 : _GEN_2095; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2097 = 8'h31 == io_state_in_8 ? 8'h2e : _GEN_2096; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2098 = 8'h32 == io_state_in_8 ? 8'ha1 : _GEN_2097; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2099 = 8'h33 == io_state_in_8 ? 8'h66 : _GEN_2098; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2100 = 8'h34 == io_state_in_8 ? 8'h28 : _GEN_2099; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2101 = 8'h35 == io_state_in_8 ? 8'hd9 : _GEN_2100; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2102 = 8'h36 == io_state_in_8 ? 8'h24 : _GEN_2101; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2103 = 8'h37 == io_state_in_8 ? 8'hb2 : _GEN_2102; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2104 = 8'h38 == io_state_in_8 ? 8'h76 : _GEN_2103; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2105 = 8'h39 == io_state_in_8 ? 8'h5b : _GEN_2104; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2106 = 8'h3a == io_state_in_8 ? 8'ha2 : _GEN_2105; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2107 = 8'h3b == io_state_in_8 ? 8'h49 : _GEN_2106; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2108 = 8'h3c == io_state_in_8 ? 8'h6d : _GEN_2107; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2109 = 8'h3d == io_state_in_8 ? 8'h8b : _GEN_2108; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2110 = 8'h3e == io_state_in_8 ? 8'hd1 : _GEN_2109; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2111 = 8'h3f == io_state_in_8 ? 8'h25 : _GEN_2110; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2112 = 8'h40 == io_state_in_8 ? 8'h72 : _GEN_2111; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2113 = 8'h41 == io_state_in_8 ? 8'hf8 : _GEN_2112; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2114 = 8'h42 == io_state_in_8 ? 8'hf6 : _GEN_2113; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2115 = 8'h43 == io_state_in_8 ? 8'h64 : _GEN_2114; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2116 = 8'h44 == io_state_in_8 ? 8'h86 : _GEN_2115; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2117 = 8'h45 == io_state_in_8 ? 8'h68 : _GEN_2116; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2118 = 8'h46 == io_state_in_8 ? 8'h98 : _GEN_2117; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2119 = 8'h47 == io_state_in_8 ? 8'h16 : _GEN_2118; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2120 = 8'h48 == io_state_in_8 ? 8'hd4 : _GEN_2119; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2121 = 8'h49 == io_state_in_8 ? 8'ha4 : _GEN_2120; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2122 = 8'h4a == io_state_in_8 ? 8'h5c : _GEN_2121; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2123 = 8'h4b == io_state_in_8 ? 8'hcc : _GEN_2122; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2124 = 8'h4c == io_state_in_8 ? 8'h5d : _GEN_2123; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2125 = 8'h4d == io_state_in_8 ? 8'h65 : _GEN_2124; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2126 = 8'h4e == io_state_in_8 ? 8'hb6 : _GEN_2125; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2127 = 8'h4f == io_state_in_8 ? 8'h92 : _GEN_2126; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2128 = 8'h50 == io_state_in_8 ? 8'h6c : _GEN_2127; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2129 = 8'h51 == io_state_in_8 ? 8'h70 : _GEN_2128; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2130 = 8'h52 == io_state_in_8 ? 8'h48 : _GEN_2129; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2131 = 8'h53 == io_state_in_8 ? 8'h50 : _GEN_2130; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2132 = 8'h54 == io_state_in_8 ? 8'hfd : _GEN_2131; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2133 = 8'h55 == io_state_in_8 ? 8'hed : _GEN_2132; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2134 = 8'h56 == io_state_in_8 ? 8'hb9 : _GEN_2133; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2135 = 8'h57 == io_state_in_8 ? 8'hda : _GEN_2134; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2136 = 8'h58 == io_state_in_8 ? 8'h5e : _GEN_2135; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2137 = 8'h59 == io_state_in_8 ? 8'h15 : _GEN_2136; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2138 = 8'h5a == io_state_in_8 ? 8'h46 : _GEN_2137; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2139 = 8'h5b == io_state_in_8 ? 8'h57 : _GEN_2138; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2140 = 8'h5c == io_state_in_8 ? 8'ha7 : _GEN_2139; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2141 = 8'h5d == io_state_in_8 ? 8'h8d : _GEN_2140; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2142 = 8'h5e == io_state_in_8 ? 8'h9d : _GEN_2141; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2143 = 8'h5f == io_state_in_8 ? 8'h84 : _GEN_2142; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2144 = 8'h60 == io_state_in_8 ? 8'h90 : _GEN_2143; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2145 = 8'h61 == io_state_in_8 ? 8'hd8 : _GEN_2144; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2146 = 8'h62 == io_state_in_8 ? 8'hab : _GEN_2145; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2147 = 8'h63 == io_state_in_8 ? 8'h0 : _GEN_2146; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2148 = 8'h64 == io_state_in_8 ? 8'h8c : _GEN_2147; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2149 = 8'h65 == io_state_in_8 ? 8'hbc : _GEN_2148; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2150 = 8'h66 == io_state_in_8 ? 8'hd3 : _GEN_2149; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2151 = 8'h67 == io_state_in_8 ? 8'ha : _GEN_2150; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2152 = 8'h68 == io_state_in_8 ? 8'hf7 : _GEN_2151; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2153 = 8'h69 == io_state_in_8 ? 8'he4 : _GEN_2152; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2154 = 8'h6a == io_state_in_8 ? 8'h58 : _GEN_2153; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2155 = 8'h6b == io_state_in_8 ? 8'h5 : _GEN_2154; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2156 = 8'h6c == io_state_in_8 ? 8'hb8 : _GEN_2155; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2157 = 8'h6d == io_state_in_8 ? 8'hb3 : _GEN_2156; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2158 = 8'h6e == io_state_in_8 ? 8'h45 : _GEN_2157; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2159 = 8'h6f == io_state_in_8 ? 8'h6 : _GEN_2158; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2160 = 8'h70 == io_state_in_8 ? 8'hd0 : _GEN_2159; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2161 = 8'h71 == io_state_in_8 ? 8'h2c : _GEN_2160; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2162 = 8'h72 == io_state_in_8 ? 8'h1e : _GEN_2161; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2163 = 8'h73 == io_state_in_8 ? 8'h8f : _GEN_2162; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2164 = 8'h74 == io_state_in_8 ? 8'hca : _GEN_2163; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2165 = 8'h75 == io_state_in_8 ? 8'h3f : _GEN_2164; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2166 = 8'h76 == io_state_in_8 ? 8'hf : _GEN_2165; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2167 = 8'h77 == io_state_in_8 ? 8'h2 : _GEN_2166; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2168 = 8'h78 == io_state_in_8 ? 8'hc1 : _GEN_2167; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2169 = 8'h79 == io_state_in_8 ? 8'haf : _GEN_2168; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2170 = 8'h7a == io_state_in_8 ? 8'hbd : _GEN_2169; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2171 = 8'h7b == io_state_in_8 ? 8'h3 : _GEN_2170; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2172 = 8'h7c == io_state_in_8 ? 8'h1 : _GEN_2171; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2173 = 8'h7d == io_state_in_8 ? 8'h13 : _GEN_2172; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2174 = 8'h7e == io_state_in_8 ? 8'h8a : _GEN_2173; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2175 = 8'h7f == io_state_in_8 ? 8'h6b : _GEN_2174; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2176 = 8'h80 == io_state_in_8 ? 8'h3a : _GEN_2175; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2177 = 8'h81 == io_state_in_8 ? 8'h91 : _GEN_2176; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2178 = 8'h82 == io_state_in_8 ? 8'h11 : _GEN_2177; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2179 = 8'h83 == io_state_in_8 ? 8'h41 : _GEN_2178; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2180 = 8'h84 == io_state_in_8 ? 8'h4f : _GEN_2179; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2181 = 8'h85 == io_state_in_8 ? 8'h67 : _GEN_2180; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2182 = 8'h86 == io_state_in_8 ? 8'hdc : _GEN_2181; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2183 = 8'h87 == io_state_in_8 ? 8'hea : _GEN_2182; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2184 = 8'h88 == io_state_in_8 ? 8'h97 : _GEN_2183; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2185 = 8'h89 == io_state_in_8 ? 8'hf2 : _GEN_2184; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2186 = 8'h8a == io_state_in_8 ? 8'hcf : _GEN_2185; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2187 = 8'h8b == io_state_in_8 ? 8'hce : _GEN_2186; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2188 = 8'h8c == io_state_in_8 ? 8'hf0 : _GEN_2187; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2189 = 8'h8d == io_state_in_8 ? 8'hb4 : _GEN_2188; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2190 = 8'h8e == io_state_in_8 ? 8'he6 : _GEN_2189; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2191 = 8'h8f == io_state_in_8 ? 8'h73 : _GEN_2190; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2192 = 8'h90 == io_state_in_8 ? 8'h96 : _GEN_2191; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2193 = 8'h91 == io_state_in_8 ? 8'hac : _GEN_2192; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2194 = 8'h92 == io_state_in_8 ? 8'h74 : _GEN_2193; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2195 = 8'h93 == io_state_in_8 ? 8'h22 : _GEN_2194; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2196 = 8'h94 == io_state_in_8 ? 8'he7 : _GEN_2195; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2197 = 8'h95 == io_state_in_8 ? 8'had : _GEN_2196; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2198 = 8'h96 == io_state_in_8 ? 8'h35 : _GEN_2197; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2199 = 8'h97 == io_state_in_8 ? 8'h85 : _GEN_2198; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2200 = 8'h98 == io_state_in_8 ? 8'he2 : _GEN_2199; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2201 = 8'h99 == io_state_in_8 ? 8'hf9 : _GEN_2200; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2202 = 8'h9a == io_state_in_8 ? 8'h37 : _GEN_2201; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2203 = 8'h9b == io_state_in_8 ? 8'he8 : _GEN_2202; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2204 = 8'h9c == io_state_in_8 ? 8'h1c : _GEN_2203; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2205 = 8'h9d == io_state_in_8 ? 8'h75 : _GEN_2204; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2206 = 8'h9e == io_state_in_8 ? 8'hdf : _GEN_2205; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2207 = 8'h9f == io_state_in_8 ? 8'h6e : _GEN_2206; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2208 = 8'ha0 == io_state_in_8 ? 8'h47 : _GEN_2207; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2209 = 8'ha1 == io_state_in_8 ? 8'hf1 : _GEN_2208; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2210 = 8'ha2 == io_state_in_8 ? 8'h1a : _GEN_2209; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2211 = 8'ha3 == io_state_in_8 ? 8'h71 : _GEN_2210; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2212 = 8'ha4 == io_state_in_8 ? 8'h1d : _GEN_2211; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2213 = 8'ha5 == io_state_in_8 ? 8'h29 : _GEN_2212; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2214 = 8'ha6 == io_state_in_8 ? 8'hc5 : _GEN_2213; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2215 = 8'ha7 == io_state_in_8 ? 8'h89 : _GEN_2214; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2216 = 8'ha8 == io_state_in_8 ? 8'h6f : _GEN_2215; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2217 = 8'ha9 == io_state_in_8 ? 8'hb7 : _GEN_2216; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2218 = 8'haa == io_state_in_8 ? 8'h62 : _GEN_2217; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2219 = 8'hab == io_state_in_8 ? 8'he : _GEN_2218; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2220 = 8'hac == io_state_in_8 ? 8'haa : _GEN_2219; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2221 = 8'had == io_state_in_8 ? 8'h18 : _GEN_2220; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2222 = 8'hae == io_state_in_8 ? 8'hbe : _GEN_2221; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2223 = 8'haf == io_state_in_8 ? 8'h1b : _GEN_2222; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2224 = 8'hb0 == io_state_in_8 ? 8'hfc : _GEN_2223; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2225 = 8'hb1 == io_state_in_8 ? 8'h56 : _GEN_2224; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2226 = 8'hb2 == io_state_in_8 ? 8'h3e : _GEN_2225; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2227 = 8'hb3 == io_state_in_8 ? 8'h4b : _GEN_2226; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2228 = 8'hb4 == io_state_in_8 ? 8'hc6 : _GEN_2227; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2229 = 8'hb5 == io_state_in_8 ? 8'hd2 : _GEN_2228; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2230 = 8'hb6 == io_state_in_8 ? 8'h79 : _GEN_2229; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2231 = 8'hb7 == io_state_in_8 ? 8'h20 : _GEN_2230; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2232 = 8'hb8 == io_state_in_8 ? 8'h9a : _GEN_2231; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2233 = 8'hb9 == io_state_in_8 ? 8'hdb : _GEN_2232; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2234 = 8'hba == io_state_in_8 ? 8'hc0 : _GEN_2233; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2235 = 8'hbb == io_state_in_8 ? 8'hfe : _GEN_2234; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2236 = 8'hbc == io_state_in_8 ? 8'h78 : _GEN_2235; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2237 = 8'hbd == io_state_in_8 ? 8'hcd : _GEN_2236; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2238 = 8'hbe == io_state_in_8 ? 8'h5a : _GEN_2237; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2239 = 8'hbf == io_state_in_8 ? 8'hf4 : _GEN_2238; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2240 = 8'hc0 == io_state_in_8 ? 8'h1f : _GEN_2239; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2241 = 8'hc1 == io_state_in_8 ? 8'hdd : _GEN_2240; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2242 = 8'hc2 == io_state_in_8 ? 8'ha8 : _GEN_2241; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2243 = 8'hc3 == io_state_in_8 ? 8'h33 : _GEN_2242; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2244 = 8'hc4 == io_state_in_8 ? 8'h88 : _GEN_2243; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2245 = 8'hc5 == io_state_in_8 ? 8'h7 : _GEN_2244; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2246 = 8'hc6 == io_state_in_8 ? 8'hc7 : _GEN_2245; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2247 = 8'hc7 == io_state_in_8 ? 8'h31 : _GEN_2246; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2248 = 8'hc8 == io_state_in_8 ? 8'hb1 : _GEN_2247; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2249 = 8'hc9 == io_state_in_8 ? 8'h12 : _GEN_2248; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2250 = 8'hca == io_state_in_8 ? 8'h10 : _GEN_2249; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2251 = 8'hcb == io_state_in_8 ? 8'h59 : _GEN_2250; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2252 = 8'hcc == io_state_in_8 ? 8'h27 : _GEN_2251; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2253 = 8'hcd == io_state_in_8 ? 8'h80 : _GEN_2252; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2254 = 8'hce == io_state_in_8 ? 8'hec : _GEN_2253; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2255 = 8'hcf == io_state_in_8 ? 8'h5f : _GEN_2254; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2256 = 8'hd0 == io_state_in_8 ? 8'h60 : _GEN_2255; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2257 = 8'hd1 == io_state_in_8 ? 8'h51 : _GEN_2256; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2258 = 8'hd2 == io_state_in_8 ? 8'h7f : _GEN_2257; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2259 = 8'hd3 == io_state_in_8 ? 8'ha9 : _GEN_2258; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2260 = 8'hd4 == io_state_in_8 ? 8'h19 : _GEN_2259; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2261 = 8'hd5 == io_state_in_8 ? 8'hb5 : _GEN_2260; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2262 = 8'hd6 == io_state_in_8 ? 8'h4a : _GEN_2261; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2263 = 8'hd7 == io_state_in_8 ? 8'hd : _GEN_2262; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2264 = 8'hd8 == io_state_in_8 ? 8'h2d : _GEN_2263; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2265 = 8'hd9 == io_state_in_8 ? 8'he5 : _GEN_2264; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2266 = 8'hda == io_state_in_8 ? 8'h7a : _GEN_2265; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2267 = 8'hdb == io_state_in_8 ? 8'h9f : _GEN_2266; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2268 = 8'hdc == io_state_in_8 ? 8'h93 : _GEN_2267; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2269 = 8'hdd == io_state_in_8 ? 8'hc9 : _GEN_2268; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2270 = 8'hde == io_state_in_8 ? 8'h9c : _GEN_2269; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2271 = 8'hdf == io_state_in_8 ? 8'hef : _GEN_2270; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2272 = 8'he0 == io_state_in_8 ? 8'ha0 : _GEN_2271; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2273 = 8'he1 == io_state_in_8 ? 8'he0 : _GEN_2272; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2274 = 8'he2 == io_state_in_8 ? 8'h3b : _GEN_2273; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2275 = 8'he3 == io_state_in_8 ? 8'h4d : _GEN_2274; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2276 = 8'he4 == io_state_in_8 ? 8'hae : _GEN_2275; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2277 = 8'he5 == io_state_in_8 ? 8'h2a : _GEN_2276; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2278 = 8'he6 == io_state_in_8 ? 8'hf5 : _GEN_2277; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2279 = 8'he7 == io_state_in_8 ? 8'hb0 : _GEN_2278; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2280 = 8'he8 == io_state_in_8 ? 8'hc8 : _GEN_2279; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2281 = 8'he9 == io_state_in_8 ? 8'heb : _GEN_2280; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2282 = 8'hea == io_state_in_8 ? 8'hbb : _GEN_2281; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2283 = 8'heb == io_state_in_8 ? 8'h3c : _GEN_2282; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2284 = 8'hec == io_state_in_8 ? 8'h83 : _GEN_2283; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2285 = 8'hed == io_state_in_8 ? 8'h53 : _GEN_2284; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2286 = 8'hee == io_state_in_8 ? 8'h99 : _GEN_2285; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2287 = 8'hef == io_state_in_8 ? 8'h61 : _GEN_2286; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2288 = 8'hf0 == io_state_in_8 ? 8'h17 : _GEN_2287; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2289 = 8'hf1 == io_state_in_8 ? 8'h2b : _GEN_2288; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2290 = 8'hf2 == io_state_in_8 ? 8'h4 : _GEN_2289; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2291 = 8'hf3 == io_state_in_8 ? 8'h7e : _GEN_2290; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2292 = 8'hf4 == io_state_in_8 ? 8'hba : _GEN_2291; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2293 = 8'hf5 == io_state_in_8 ? 8'h77 : _GEN_2292; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2294 = 8'hf6 == io_state_in_8 ? 8'hd6 : _GEN_2293; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2295 = 8'hf7 == io_state_in_8 ? 8'h26 : _GEN_2294; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2296 = 8'hf8 == io_state_in_8 ? 8'he1 : _GEN_2295; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2297 = 8'hf9 == io_state_in_8 ? 8'h69 : _GEN_2296; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2298 = 8'hfa == io_state_in_8 ? 8'h14 : _GEN_2297; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2299 = 8'hfb == io_state_in_8 ? 8'h63 : _GEN_2298; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2300 = 8'hfc == io_state_in_8 ? 8'h55 : _GEN_2299; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2301 = 8'hfd == io_state_in_8 ? 8'h21 : _GEN_2300; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2302 = 8'hfe == io_state_in_8 ? 8'hc : _GEN_2301; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2305 = 8'h1 == io_state_in_9 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2306 = 8'h2 == io_state_in_9 ? 8'h6a : _GEN_2305; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2307 = 8'h3 == io_state_in_9 ? 8'hd5 : _GEN_2306; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2308 = 8'h4 == io_state_in_9 ? 8'h30 : _GEN_2307; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2309 = 8'h5 == io_state_in_9 ? 8'h36 : _GEN_2308; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2310 = 8'h6 == io_state_in_9 ? 8'ha5 : _GEN_2309; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2311 = 8'h7 == io_state_in_9 ? 8'h38 : _GEN_2310; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2312 = 8'h8 == io_state_in_9 ? 8'hbf : _GEN_2311; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2313 = 8'h9 == io_state_in_9 ? 8'h40 : _GEN_2312; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2314 = 8'ha == io_state_in_9 ? 8'ha3 : _GEN_2313; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2315 = 8'hb == io_state_in_9 ? 8'h9e : _GEN_2314; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2316 = 8'hc == io_state_in_9 ? 8'h81 : _GEN_2315; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2317 = 8'hd == io_state_in_9 ? 8'hf3 : _GEN_2316; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2318 = 8'he == io_state_in_9 ? 8'hd7 : _GEN_2317; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2319 = 8'hf == io_state_in_9 ? 8'hfb : _GEN_2318; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2320 = 8'h10 == io_state_in_9 ? 8'h7c : _GEN_2319; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2321 = 8'h11 == io_state_in_9 ? 8'he3 : _GEN_2320; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2322 = 8'h12 == io_state_in_9 ? 8'h39 : _GEN_2321; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2323 = 8'h13 == io_state_in_9 ? 8'h82 : _GEN_2322; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2324 = 8'h14 == io_state_in_9 ? 8'h9b : _GEN_2323; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2325 = 8'h15 == io_state_in_9 ? 8'h2f : _GEN_2324; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2326 = 8'h16 == io_state_in_9 ? 8'hff : _GEN_2325; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2327 = 8'h17 == io_state_in_9 ? 8'h87 : _GEN_2326; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2328 = 8'h18 == io_state_in_9 ? 8'h34 : _GEN_2327; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2329 = 8'h19 == io_state_in_9 ? 8'h8e : _GEN_2328; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2330 = 8'h1a == io_state_in_9 ? 8'h43 : _GEN_2329; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2331 = 8'h1b == io_state_in_9 ? 8'h44 : _GEN_2330; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2332 = 8'h1c == io_state_in_9 ? 8'hc4 : _GEN_2331; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2333 = 8'h1d == io_state_in_9 ? 8'hde : _GEN_2332; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2334 = 8'h1e == io_state_in_9 ? 8'he9 : _GEN_2333; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2335 = 8'h1f == io_state_in_9 ? 8'hcb : _GEN_2334; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2336 = 8'h20 == io_state_in_9 ? 8'h54 : _GEN_2335; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2337 = 8'h21 == io_state_in_9 ? 8'h7b : _GEN_2336; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2338 = 8'h22 == io_state_in_9 ? 8'h94 : _GEN_2337; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2339 = 8'h23 == io_state_in_9 ? 8'h32 : _GEN_2338; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2340 = 8'h24 == io_state_in_9 ? 8'ha6 : _GEN_2339; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2341 = 8'h25 == io_state_in_9 ? 8'hc2 : _GEN_2340; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2342 = 8'h26 == io_state_in_9 ? 8'h23 : _GEN_2341; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2343 = 8'h27 == io_state_in_9 ? 8'h3d : _GEN_2342; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2344 = 8'h28 == io_state_in_9 ? 8'hee : _GEN_2343; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2345 = 8'h29 == io_state_in_9 ? 8'h4c : _GEN_2344; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2346 = 8'h2a == io_state_in_9 ? 8'h95 : _GEN_2345; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2347 = 8'h2b == io_state_in_9 ? 8'hb : _GEN_2346; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2348 = 8'h2c == io_state_in_9 ? 8'h42 : _GEN_2347; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2349 = 8'h2d == io_state_in_9 ? 8'hfa : _GEN_2348; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2350 = 8'h2e == io_state_in_9 ? 8'hc3 : _GEN_2349; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2351 = 8'h2f == io_state_in_9 ? 8'h4e : _GEN_2350; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2352 = 8'h30 == io_state_in_9 ? 8'h8 : _GEN_2351; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2353 = 8'h31 == io_state_in_9 ? 8'h2e : _GEN_2352; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2354 = 8'h32 == io_state_in_9 ? 8'ha1 : _GEN_2353; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2355 = 8'h33 == io_state_in_9 ? 8'h66 : _GEN_2354; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2356 = 8'h34 == io_state_in_9 ? 8'h28 : _GEN_2355; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2357 = 8'h35 == io_state_in_9 ? 8'hd9 : _GEN_2356; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2358 = 8'h36 == io_state_in_9 ? 8'h24 : _GEN_2357; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2359 = 8'h37 == io_state_in_9 ? 8'hb2 : _GEN_2358; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2360 = 8'h38 == io_state_in_9 ? 8'h76 : _GEN_2359; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2361 = 8'h39 == io_state_in_9 ? 8'h5b : _GEN_2360; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2362 = 8'h3a == io_state_in_9 ? 8'ha2 : _GEN_2361; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2363 = 8'h3b == io_state_in_9 ? 8'h49 : _GEN_2362; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2364 = 8'h3c == io_state_in_9 ? 8'h6d : _GEN_2363; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2365 = 8'h3d == io_state_in_9 ? 8'h8b : _GEN_2364; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2366 = 8'h3e == io_state_in_9 ? 8'hd1 : _GEN_2365; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2367 = 8'h3f == io_state_in_9 ? 8'h25 : _GEN_2366; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2368 = 8'h40 == io_state_in_9 ? 8'h72 : _GEN_2367; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2369 = 8'h41 == io_state_in_9 ? 8'hf8 : _GEN_2368; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2370 = 8'h42 == io_state_in_9 ? 8'hf6 : _GEN_2369; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2371 = 8'h43 == io_state_in_9 ? 8'h64 : _GEN_2370; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2372 = 8'h44 == io_state_in_9 ? 8'h86 : _GEN_2371; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2373 = 8'h45 == io_state_in_9 ? 8'h68 : _GEN_2372; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2374 = 8'h46 == io_state_in_9 ? 8'h98 : _GEN_2373; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2375 = 8'h47 == io_state_in_9 ? 8'h16 : _GEN_2374; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2376 = 8'h48 == io_state_in_9 ? 8'hd4 : _GEN_2375; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2377 = 8'h49 == io_state_in_9 ? 8'ha4 : _GEN_2376; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2378 = 8'h4a == io_state_in_9 ? 8'h5c : _GEN_2377; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2379 = 8'h4b == io_state_in_9 ? 8'hcc : _GEN_2378; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2380 = 8'h4c == io_state_in_9 ? 8'h5d : _GEN_2379; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2381 = 8'h4d == io_state_in_9 ? 8'h65 : _GEN_2380; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2382 = 8'h4e == io_state_in_9 ? 8'hb6 : _GEN_2381; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2383 = 8'h4f == io_state_in_9 ? 8'h92 : _GEN_2382; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2384 = 8'h50 == io_state_in_9 ? 8'h6c : _GEN_2383; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2385 = 8'h51 == io_state_in_9 ? 8'h70 : _GEN_2384; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2386 = 8'h52 == io_state_in_9 ? 8'h48 : _GEN_2385; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2387 = 8'h53 == io_state_in_9 ? 8'h50 : _GEN_2386; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2388 = 8'h54 == io_state_in_9 ? 8'hfd : _GEN_2387; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2389 = 8'h55 == io_state_in_9 ? 8'hed : _GEN_2388; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2390 = 8'h56 == io_state_in_9 ? 8'hb9 : _GEN_2389; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2391 = 8'h57 == io_state_in_9 ? 8'hda : _GEN_2390; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2392 = 8'h58 == io_state_in_9 ? 8'h5e : _GEN_2391; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2393 = 8'h59 == io_state_in_9 ? 8'h15 : _GEN_2392; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2394 = 8'h5a == io_state_in_9 ? 8'h46 : _GEN_2393; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2395 = 8'h5b == io_state_in_9 ? 8'h57 : _GEN_2394; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2396 = 8'h5c == io_state_in_9 ? 8'ha7 : _GEN_2395; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2397 = 8'h5d == io_state_in_9 ? 8'h8d : _GEN_2396; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2398 = 8'h5e == io_state_in_9 ? 8'h9d : _GEN_2397; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2399 = 8'h5f == io_state_in_9 ? 8'h84 : _GEN_2398; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2400 = 8'h60 == io_state_in_9 ? 8'h90 : _GEN_2399; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2401 = 8'h61 == io_state_in_9 ? 8'hd8 : _GEN_2400; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2402 = 8'h62 == io_state_in_9 ? 8'hab : _GEN_2401; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2403 = 8'h63 == io_state_in_9 ? 8'h0 : _GEN_2402; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2404 = 8'h64 == io_state_in_9 ? 8'h8c : _GEN_2403; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2405 = 8'h65 == io_state_in_9 ? 8'hbc : _GEN_2404; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2406 = 8'h66 == io_state_in_9 ? 8'hd3 : _GEN_2405; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2407 = 8'h67 == io_state_in_9 ? 8'ha : _GEN_2406; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2408 = 8'h68 == io_state_in_9 ? 8'hf7 : _GEN_2407; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2409 = 8'h69 == io_state_in_9 ? 8'he4 : _GEN_2408; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2410 = 8'h6a == io_state_in_9 ? 8'h58 : _GEN_2409; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2411 = 8'h6b == io_state_in_9 ? 8'h5 : _GEN_2410; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2412 = 8'h6c == io_state_in_9 ? 8'hb8 : _GEN_2411; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2413 = 8'h6d == io_state_in_9 ? 8'hb3 : _GEN_2412; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2414 = 8'h6e == io_state_in_9 ? 8'h45 : _GEN_2413; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2415 = 8'h6f == io_state_in_9 ? 8'h6 : _GEN_2414; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2416 = 8'h70 == io_state_in_9 ? 8'hd0 : _GEN_2415; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2417 = 8'h71 == io_state_in_9 ? 8'h2c : _GEN_2416; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2418 = 8'h72 == io_state_in_9 ? 8'h1e : _GEN_2417; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2419 = 8'h73 == io_state_in_9 ? 8'h8f : _GEN_2418; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2420 = 8'h74 == io_state_in_9 ? 8'hca : _GEN_2419; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2421 = 8'h75 == io_state_in_9 ? 8'h3f : _GEN_2420; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2422 = 8'h76 == io_state_in_9 ? 8'hf : _GEN_2421; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2423 = 8'h77 == io_state_in_9 ? 8'h2 : _GEN_2422; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2424 = 8'h78 == io_state_in_9 ? 8'hc1 : _GEN_2423; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2425 = 8'h79 == io_state_in_9 ? 8'haf : _GEN_2424; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2426 = 8'h7a == io_state_in_9 ? 8'hbd : _GEN_2425; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2427 = 8'h7b == io_state_in_9 ? 8'h3 : _GEN_2426; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2428 = 8'h7c == io_state_in_9 ? 8'h1 : _GEN_2427; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2429 = 8'h7d == io_state_in_9 ? 8'h13 : _GEN_2428; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2430 = 8'h7e == io_state_in_9 ? 8'h8a : _GEN_2429; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2431 = 8'h7f == io_state_in_9 ? 8'h6b : _GEN_2430; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2432 = 8'h80 == io_state_in_9 ? 8'h3a : _GEN_2431; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2433 = 8'h81 == io_state_in_9 ? 8'h91 : _GEN_2432; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2434 = 8'h82 == io_state_in_9 ? 8'h11 : _GEN_2433; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2435 = 8'h83 == io_state_in_9 ? 8'h41 : _GEN_2434; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2436 = 8'h84 == io_state_in_9 ? 8'h4f : _GEN_2435; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2437 = 8'h85 == io_state_in_9 ? 8'h67 : _GEN_2436; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2438 = 8'h86 == io_state_in_9 ? 8'hdc : _GEN_2437; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2439 = 8'h87 == io_state_in_9 ? 8'hea : _GEN_2438; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2440 = 8'h88 == io_state_in_9 ? 8'h97 : _GEN_2439; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2441 = 8'h89 == io_state_in_9 ? 8'hf2 : _GEN_2440; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2442 = 8'h8a == io_state_in_9 ? 8'hcf : _GEN_2441; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2443 = 8'h8b == io_state_in_9 ? 8'hce : _GEN_2442; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2444 = 8'h8c == io_state_in_9 ? 8'hf0 : _GEN_2443; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2445 = 8'h8d == io_state_in_9 ? 8'hb4 : _GEN_2444; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2446 = 8'h8e == io_state_in_9 ? 8'he6 : _GEN_2445; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2447 = 8'h8f == io_state_in_9 ? 8'h73 : _GEN_2446; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2448 = 8'h90 == io_state_in_9 ? 8'h96 : _GEN_2447; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2449 = 8'h91 == io_state_in_9 ? 8'hac : _GEN_2448; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2450 = 8'h92 == io_state_in_9 ? 8'h74 : _GEN_2449; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2451 = 8'h93 == io_state_in_9 ? 8'h22 : _GEN_2450; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2452 = 8'h94 == io_state_in_9 ? 8'he7 : _GEN_2451; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2453 = 8'h95 == io_state_in_9 ? 8'had : _GEN_2452; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2454 = 8'h96 == io_state_in_9 ? 8'h35 : _GEN_2453; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2455 = 8'h97 == io_state_in_9 ? 8'h85 : _GEN_2454; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2456 = 8'h98 == io_state_in_9 ? 8'he2 : _GEN_2455; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2457 = 8'h99 == io_state_in_9 ? 8'hf9 : _GEN_2456; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2458 = 8'h9a == io_state_in_9 ? 8'h37 : _GEN_2457; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2459 = 8'h9b == io_state_in_9 ? 8'he8 : _GEN_2458; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2460 = 8'h9c == io_state_in_9 ? 8'h1c : _GEN_2459; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2461 = 8'h9d == io_state_in_9 ? 8'h75 : _GEN_2460; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2462 = 8'h9e == io_state_in_9 ? 8'hdf : _GEN_2461; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2463 = 8'h9f == io_state_in_9 ? 8'h6e : _GEN_2462; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2464 = 8'ha0 == io_state_in_9 ? 8'h47 : _GEN_2463; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2465 = 8'ha1 == io_state_in_9 ? 8'hf1 : _GEN_2464; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2466 = 8'ha2 == io_state_in_9 ? 8'h1a : _GEN_2465; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2467 = 8'ha3 == io_state_in_9 ? 8'h71 : _GEN_2466; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2468 = 8'ha4 == io_state_in_9 ? 8'h1d : _GEN_2467; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2469 = 8'ha5 == io_state_in_9 ? 8'h29 : _GEN_2468; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2470 = 8'ha6 == io_state_in_9 ? 8'hc5 : _GEN_2469; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2471 = 8'ha7 == io_state_in_9 ? 8'h89 : _GEN_2470; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2472 = 8'ha8 == io_state_in_9 ? 8'h6f : _GEN_2471; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2473 = 8'ha9 == io_state_in_9 ? 8'hb7 : _GEN_2472; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2474 = 8'haa == io_state_in_9 ? 8'h62 : _GEN_2473; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2475 = 8'hab == io_state_in_9 ? 8'he : _GEN_2474; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2476 = 8'hac == io_state_in_9 ? 8'haa : _GEN_2475; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2477 = 8'had == io_state_in_9 ? 8'h18 : _GEN_2476; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2478 = 8'hae == io_state_in_9 ? 8'hbe : _GEN_2477; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2479 = 8'haf == io_state_in_9 ? 8'h1b : _GEN_2478; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2480 = 8'hb0 == io_state_in_9 ? 8'hfc : _GEN_2479; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2481 = 8'hb1 == io_state_in_9 ? 8'h56 : _GEN_2480; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2482 = 8'hb2 == io_state_in_9 ? 8'h3e : _GEN_2481; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2483 = 8'hb3 == io_state_in_9 ? 8'h4b : _GEN_2482; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2484 = 8'hb4 == io_state_in_9 ? 8'hc6 : _GEN_2483; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2485 = 8'hb5 == io_state_in_9 ? 8'hd2 : _GEN_2484; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2486 = 8'hb6 == io_state_in_9 ? 8'h79 : _GEN_2485; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2487 = 8'hb7 == io_state_in_9 ? 8'h20 : _GEN_2486; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2488 = 8'hb8 == io_state_in_9 ? 8'h9a : _GEN_2487; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2489 = 8'hb9 == io_state_in_9 ? 8'hdb : _GEN_2488; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2490 = 8'hba == io_state_in_9 ? 8'hc0 : _GEN_2489; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2491 = 8'hbb == io_state_in_9 ? 8'hfe : _GEN_2490; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2492 = 8'hbc == io_state_in_9 ? 8'h78 : _GEN_2491; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2493 = 8'hbd == io_state_in_9 ? 8'hcd : _GEN_2492; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2494 = 8'hbe == io_state_in_9 ? 8'h5a : _GEN_2493; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2495 = 8'hbf == io_state_in_9 ? 8'hf4 : _GEN_2494; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2496 = 8'hc0 == io_state_in_9 ? 8'h1f : _GEN_2495; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2497 = 8'hc1 == io_state_in_9 ? 8'hdd : _GEN_2496; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2498 = 8'hc2 == io_state_in_9 ? 8'ha8 : _GEN_2497; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2499 = 8'hc3 == io_state_in_9 ? 8'h33 : _GEN_2498; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2500 = 8'hc4 == io_state_in_9 ? 8'h88 : _GEN_2499; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2501 = 8'hc5 == io_state_in_9 ? 8'h7 : _GEN_2500; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2502 = 8'hc6 == io_state_in_9 ? 8'hc7 : _GEN_2501; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2503 = 8'hc7 == io_state_in_9 ? 8'h31 : _GEN_2502; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2504 = 8'hc8 == io_state_in_9 ? 8'hb1 : _GEN_2503; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2505 = 8'hc9 == io_state_in_9 ? 8'h12 : _GEN_2504; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2506 = 8'hca == io_state_in_9 ? 8'h10 : _GEN_2505; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2507 = 8'hcb == io_state_in_9 ? 8'h59 : _GEN_2506; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2508 = 8'hcc == io_state_in_9 ? 8'h27 : _GEN_2507; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2509 = 8'hcd == io_state_in_9 ? 8'h80 : _GEN_2508; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2510 = 8'hce == io_state_in_9 ? 8'hec : _GEN_2509; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2511 = 8'hcf == io_state_in_9 ? 8'h5f : _GEN_2510; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2512 = 8'hd0 == io_state_in_9 ? 8'h60 : _GEN_2511; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2513 = 8'hd1 == io_state_in_9 ? 8'h51 : _GEN_2512; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2514 = 8'hd2 == io_state_in_9 ? 8'h7f : _GEN_2513; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2515 = 8'hd3 == io_state_in_9 ? 8'ha9 : _GEN_2514; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2516 = 8'hd4 == io_state_in_9 ? 8'h19 : _GEN_2515; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2517 = 8'hd5 == io_state_in_9 ? 8'hb5 : _GEN_2516; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2518 = 8'hd6 == io_state_in_9 ? 8'h4a : _GEN_2517; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2519 = 8'hd7 == io_state_in_9 ? 8'hd : _GEN_2518; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2520 = 8'hd8 == io_state_in_9 ? 8'h2d : _GEN_2519; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2521 = 8'hd9 == io_state_in_9 ? 8'he5 : _GEN_2520; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2522 = 8'hda == io_state_in_9 ? 8'h7a : _GEN_2521; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2523 = 8'hdb == io_state_in_9 ? 8'h9f : _GEN_2522; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2524 = 8'hdc == io_state_in_9 ? 8'h93 : _GEN_2523; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2525 = 8'hdd == io_state_in_9 ? 8'hc9 : _GEN_2524; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2526 = 8'hde == io_state_in_9 ? 8'h9c : _GEN_2525; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2527 = 8'hdf == io_state_in_9 ? 8'hef : _GEN_2526; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2528 = 8'he0 == io_state_in_9 ? 8'ha0 : _GEN_2527; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2529 = 8'he1 == io_state_in_9 ? 8'he0 : _GEN_2528; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2530 = 8'he2 == io_state_in_9 ? 8'h3b : _GEN_2529; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2531 = 8'he3 == io_state_in_9 ? 8'h4d : _GEN_2530; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2532 = 8'he4 == io_state_in_9 ? 8'hae : _GEN_2531; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2533 = 8'he5 == io_state_in_9 ? 8'h2a : _GEN_2532; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2534 = 8'he6 == io_state_in_9 ? 8'hf5 : _GEN_2533; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2535 = 8'he7 == io_state_in_9 ? 8'hb0 : _GEN_2534; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2536 = 8'he8 == io_state_in_9 ? 8'hc8 : _GEN_2535; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2537 = 8'he9 == io_state_in_9 ? 8'heb : _GEN_2536; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2538 = 8'hea == io_state_in_9 ? 8'hbb : _GEN_2537; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2539 = 8'heb == io_state_in_9 ? 8'h3c : _GEN_2538; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2540 = 8'hec == io_state_in_9 ? 8'h83 : _GEN_2539; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2541 = 8'hed == io_state_in_9 ? 8'h53 : _GEN_2540; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2542 = 8'hee == io_state_in_9 ? 8'h99 : _GEN_2541; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2543 = 8'hef == io_state_in_9 ? 8'h61 : _GEN_2542; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2544 = 8'hf0 == io_state_in_9 ? 8'h17 : _GEN_2543; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2545 = 8'hf1 == io_state_in_9 ? 8'h2b : _GEN_2544; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2546 = 8'hf2 == io_state_in_9 ? 8'h4 : _GEN_2545; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2547 = 8'hf3 == io_state_in_9 ? 8'h7e : _GEN_2546; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2548 = 8'hf4 == io_state_in_9 ? 8'hba : _GEN_2547; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2549 = 8'hf5 == io_state_in_9 ? 8'h77 : _GEN_2548; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2550 = 8'hf6 == io_state_in_9 ? 8'hd6 : _GEN_2549; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2551 = 8'hf7 == io_state_in_9 ? 8'h26 : _GEN_2550; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2552 = 8'hf8 == io_state_in_9 ? 8'he1 : _GEN_2551; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2553 = 8'hf9 == io_state_in_9 ? 8'h69 : _GEN_2552; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2554 = 8'hfa == io_state_in_9 ? 8'h14 : _GEN_2553; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2555 = 8'hfb == io_state_in_9 ? 8'h63 : _GEN_2554; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2556 = 8'hfc == io_state_in_9 ? 8'h55 : _GEN_2555; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2557 = 8'hfd == io_state_in_9 ? 8'h21 : _GEN_2556; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2558 = 8'hfe == io_state_in_9 ? 8'hc : _GEN_2557; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2561 = 8'h1 == io_state_in_10 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2562 = 8'h2 == io_state_in_10 ? 8'h6a : _GEN_2561; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2563 = 8'h3 == io_state_in_10 ? 8'hd5 : _GEN_2562; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2564 = 8'h4 == io_state_in_10 ? 8'h30 : _GEN_2563; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2565 = 8'h5 == io_state_in_10 ? 8'h36 : _GEN_2564; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2566 = 8'h6 == io_state_in_10 ? 8'ha5 : _GEN_2565; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2567 = 8'h7 == io_state_in_10 ? 8'h38 : _GEN_2566; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2568 = 8'h8 == io_state_in_10 ? 8'hbf : _GEN_2567; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2569 = 8'h9 == io_state_in_10 ? 8'h40 : _GEN_2568; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2570 = 8'ha == io_state_in_10 ? 8'ha3 : _GEN_2569; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2571 = 8'hb == io_state_in_10 ? 8'h9e : _GEN_2570; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2572 = 8'hc == io_state_in_10 ? 8'h81 : _GEN_2571; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2573 = 8'hd == io_state_in_10 ? 8'hf3 : _GEN_2572; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2574 = 8'he == io_state_in_10 ? 8'hd7 : _GEN_2573; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2575 = 8'hf == io_state_in_10 ? 8'hfb : _GEN_2574; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2576 = 8'h10 == io_state_in_10 ? 8'h7c : _GEN_2575; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2577 = 8'h11 == io_state_in_10 ? 8'he3 : _GEN_2576; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2578 = 8'h12 == io_state_in_10 ? 8'h39 : _GEN_2577; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2579 = 8'h13 == io_state_in_10 ? 8'h82 : _GEN_2578; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2580 = 8'h14 == io_state_in_10 ? 8'h9b : _GEN_2579; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2581 = 8'h15 == io_state_in_10 ? 8'h2f : _GEN_2580; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2582 = 8'h16 == io_state_in_10 ? 8'hff : _GEN_2581; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2583 = 8'h17 == io_state_in_10 ? 8'h87 : _GEN_2582; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2584 = 8'h18 == io_state_in_10 ? 8'h34 : _GEN_2583; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2585 = 8'h19 == io_state_in_10 ? 8'h8e : _GEN_2584; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2586 = 8'h1a == io_state_in_10 ? 8'h43 : _GEN_2585; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2587 = 8'h1b == io_state_in_10 ? 8'h44 : _GEN_2586; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2588 = 8'h1c == io_state_in_10 ? 8'hc4 : _GEN_2587; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2589 = 8'h1d == io_state_in_10 ? 8'hde : _GEN_2588; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2590 = 8'h1e == io_state_in_10 ? 8'he9 : _GEN_2589; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2591 = 8'h1f == io_state_in_10 ? 8'hcb : _GEN_2590; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2592 = 8'h20 == io_state_in_10 ? 8'h54 : _GEN_2591; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2593 = 8'h21 == io_state_in_10 ? 8'h7b : _GEN_2592; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2594 = 8'h22 == io_state_in_10 ? 8'h94 : _GEN_2593; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2595 = 8'h23 == io_state_in_10 ? 8'h32 : _GEN_2594; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2596 = 8'h24 == io_state_in_10 ? 8'ha6 : _GEN_2595; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2597 = 8'h25 == io_state_in_10 ? 8'hc2 : _GEN_2596; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2598 = 8'h26 == io_state_in_10 ? 8'h23 : _GEN_2597; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2599 = 8'h27 == io_state_in_10 ? 8'h3d : _GEN_2598; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2600 = 8'h28 == io_state_in_10 ? 8'hee : _GEN_2599; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2601 = 8'h29 == io_state_in_10 ? 8'h4c : _GEN_2600; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2602 = 8'h2a == io_state_in_10 ? 8'h95 : _GEN_2601; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2603 = 8'h2b == io_state_in_10 ? 8'hb : _GEN_2602; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2604 = 8'h2c == io_state_in_10 ? 8'h42 : _GEN_2603; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2605 = 8'h2d == io_state_in_10 ? 8'hfa : _GEN_2604; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2606 = 8'h2e == io_state_in_10 ? 8'hc3 : _GEN_2605; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2607 = 8'h2f == io_state_in_10 ? 8'h4e : _GEN_2606; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2608 = 8'h30 == io_state_in_10 ? 8'h8 : _GEN_2607; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2609 = 8'h31 == io_state_in_10 ? 8'h2e : _GEN_2608; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2610 = 8'h32 == io_state_in_10 ? 8'ha1 : _GEN_2609; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2611 = 8'h33 == io_state_in_10 ? 8'h66 : _GEN_2610; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2612 = 8'h34 == io_state_in_10 ? 8'h28 : _GEN_2611; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2613 = 8'h35 == io_state_in_10 ? 8'hd9 : _GEN_2612; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2614 = 8'h36 == io_state_in_10 ? 8'h24 : _GEN_2613; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2615 = 8'h37 == io_state_in_10 ? 8'hb2 : _GEN_2614; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2616 = 8'h38 == io_state_in_10 ? 8'h76 : _GEN_2615; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2617 = 8'h39 == io_state_in_10 ? 8'h5b : _GEN_2616; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2618 = 8'h3a == io_state_in_10 ? 8'ha2 : _GEN_2617; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2619 = 8'h3b == io_state_in_10 ? 8'h49 : _GEN_2618; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2620 = 8'h3c == io_state_in_10 ? 8'h6d : _GEN_2619; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2621 = 8'h3d == io_state_in_10 ? 8'h8b : _GEN_2620; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2622 = 8'h3e == io_state_in_10 ? 8'hd1 : _GEN_2621; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2623 = 8'h3f == io_state_in_10 ? 8'h25 : _GEN_2622; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2624 = 8'h40 == io_state_in_10 ? 8'h72 : _GEN_2623; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2625 = 8'h41 == io_state_in_10 ? 8'hf8 : _GEN_2624; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2626 = 8'h42 == io_state_in_10 ? 8'hf6 : _GEN_2625; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2627 = 8'h43 == io_state_in_10 ? 8'h64 : _GEN_2626; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2628 = 8'h44 == io_state_in_10 ? 8'h86 : _GEN_2627; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2629 = 8'h45 == io_state_in_10 ? 8'h68 : _GEN_2628; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2630 = 8'h46 == io_state_in_10 ? 8'h98 : _GEN_2629; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2631 = 8'h47 == io_state_in_10 ? 8'h16 : _GEN_2630; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2632 = 8'h48 == io_state_in_10 ? 8'hd4 : _GEN_2631; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2633 = 8'h49 == io_state_in_10 ? 8'ha4 : _GEN_2632; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2634 = 8'h4a == io_state_in_10 ? 8'h5c : _GEN_2633; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2635 = 8'h4b == io_state_in_10 ? 8'hcc : _GEN_2634; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2636 = 8'h4c == io_state_in_10 ? 8'h5d : _GEN_2635; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2637 = 8'h4d == io_state_in_10 ? 8'h65 : _GEN_2636; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2638 = 8'h4e == io_state_in_10 ? 8'hb6 : _GEN_2637; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2639 = 8'h4f == io_state_in_10 ? 8'h92 : _GEN_2638; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2640 = 8'h50 == io_state_in_10 ? 8'h6c : _GEN_2639; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2641 = 8'h51 == io_state_in_10 ? 8'h70 : _GEN_2640; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2642 = 8'h52 == io_state_in_10 ? 8'h48 : _GEN_2641; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2643 = 8'h53 == io_state_in_10 ? 8'h50 : _GEN_2642; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2644 = 8'h54 == io_state_in_10 ? 8'hfd : _GEN_2643; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2645 = 8'h55 == io_state_in_10 ? 8'hed : _GEN_2644; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2646 = 8'h56 == io_state_in_10 ? 8'hb9 : _GEN_2645; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2647 = 8'h57 == io_state_in_10 ? 8'hda : _GEN_2646; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2648 = 8'h58 == io_state_in_10 ? 8'h5e : _GEN_2647; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2649 = 8'h59 == io_state_in_10 ? 8'h15 : _GEN_2648; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2650 = 8'h5a == io_state_in_10 ? 8'h46 : _GEN_2649; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2651 = 8'h5b == io_state_in_10 ? 8'h57 : _GEN_2650; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2652 = 8'h5c == io_state_in_10 ? 8'ha7 : _GEN_2651; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2653 = 8'h5d == io_state_in_10 ? 8'h8d : _GEN_2652; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2654 = 8'h5e == io_state_in_10 ? 8'h9d : _GEN_2653; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2655 = 8'h5f == io_state_in_10 ? 8'h84 : _GEN_2654; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2656 = 8'h60 == io_state_in_10 ? 8'h90 : _GEN_2655; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2657 = 8'h61 == io_state_in_10 ? 8'hd8 : _GEN_2656; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2658 = 8'h62 == io_state_in_10 ? 8'hab : _GEN_2657; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2659 = 8'h63 == io_state_in_10 ? 8'h0 : _GEN_2658; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2660 = 8'h64 == io_state_in_10 ? 8'h8c : _GEN_2659; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2661 = 8'h65 == io_state_in_10 ? 8'hbc : _GEN_2660; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2662 = 8'h66 == io_state_in_10 ? 8'hd3 : _GEN_2661; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2663 = 8'h67 == io_state_in_10 ? 8'ha : _GEN_2662; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2664 = 8'h68 == io_state_in_10 ? 8'hf7 : _GEN_2663; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2665 = 8'h69 == io_state_in_10 ? 8'he4 : _GEN_2664; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2666 = 8'h6a == io_state_in_10 ? 8'h58 : _GEN_2665; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2667 = 8'h6b == io_state_in_10 ? 8'h5 : _GEN_2666; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2668 = 8'h6c == io_state_in_10 ? 8'hb8 : _GEN_2667; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2669 = 8'h6d == io_state_in_10 ? 8'hb3 : _GEN_2668; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2670 = 8'h6e == io_state_in_10 ? 8'h45 : _GEN_2669; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2671 = 8'h6f == io_state_in_10 ? 8'h6 : _GEN_2670; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2672 = 8'h70 == io_state_in_10 ? 8'hd0 : _GEN_2671; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2673 = 8'h71 == io_state_in_10 ? 8'h2c : _GEN_2672; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2674 = 8'h72 == io_state_in_10 ? 8'h1e : _GEN_2673; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2675 = 8'h73 == io_state_in_10 ? 8'h8f : _GEN_2674; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2676 = 8'h74 == io_state_in_10 ? 8'hca : _GEN_2675; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2677 = 8'h75 == io_state_in_10 ? 8'h3f : _GEN_2676; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2678 = 8'h76 == io_state_in_10 ? 8'hf : _GEN_2677; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2679 = 8'h77 == io_state_in_10 ? 8'h2 : _GEN_2678; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2680 = 8'h78 == io_state_in_10 ? 8'hc1 : _GEN_2679; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2681 = 8'h79 == io_state_in_10 ? 8'haf : _GEN_2680; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2682 = 8'h7a == io_state_in_10 ? 8'hbd : _GEN_2681; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2683 = 8'h7b == io_state_in_10 ? 8'h3 : _GEN_2682; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2684 = 8'h7c == io_state_in_10 ? 8'h1 : _GEN_2683; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2685 = 8'h7d == io_state_in_10 ? 8'h13 : _GEN_2684; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2686 = 8'h7e == io_state_in_10 ? 8'h8a : _GEN_2685; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2687 = 8'h7f == io_state_in_10 ? 8'h6b : _GEN_2686; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2688 = 8'h80 == io_state_in_10 ? 8'h3a : _GEN_2687; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2689 = 8'h81 == io_state_in_10 ? 8'h91 : _GEN_2688; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2690 = 8'h82 == io_state_in_10 ? 8'h11 : _GEN_2689; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2691 = 8'h83 == io_state_in_10 ? 8'h41 : _GEN_2690; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2692 = 8'h84 == io_state_in_10 ? 8'h4f : _GEN_2691; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2693 = 8'h85 == io_state_in_10 ? 8'h67 : _GEN_2692; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2694 = 8'h86 == io_state_in_10 ? 8'hdc : _GEN_2693; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2695 = 8'h87 == io_state_in_10 ? 8'hea : _GEN_2694; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2696 = 8'h88 == io_state_in_10 ? 8'h97 : _GEN_2695; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2697 = 8'h89 == io_state_in_10 ? 8'hf2 : _GEN_2696; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2698 = 8'h8a == io_state_in_10 ? 8'hcf : _GEN_2697; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2699 = 8'h8b == io_state_in_10 ? 8'hce : _GEN_2698; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2700 = 8'h8c == io_state_in_10 ? 8'hf0 : _GEN_2699; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2701 = 8'h8d == io_state_in_10 ? 8'hb4 : _GEN_2700; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2702 = 8'h8e == io_state_in_10 ? 8'he6 : _GEN_2701; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2703 = 8'h8f == io_state_in_10 ? 8'h73 : _GEN_2702; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2704 = 8'h90 == io_state_in_10 ? 8'h96 : _GEN_2703; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2705 = 8'h91 == io_state_in_10 ? 8'hac : _GEN_2704; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2706 = 8'h92 == io_state_in_10 ? 8'h74 : _GEN_2705; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2707 = 8'h93 == io_state_in_10 ? 8'h22 : _GEN_2706; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2708 = 8'h94 == io_state_in_10 ? 8'he7 : _GEN_2707; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2709 = 8'h95 == io_state_in_10 ? 8'had : _GEN_2708; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2710 = 8'h96 == io_state_in_10 ? 8'h35 : _GEN_2709; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2711 = 8'h97 == io_state_in_10 ? 8'h85 : _GEN_2710; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2712 = 8'h98 == io_state_in_10 ? 8'he2 : _GEN_2711; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2713 = 8'h99 == io_state_in_10 ? 8'hf9 : _GEN_2712; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2714 = 8'h9a == io_state_in_10 ? 8'h37 : _GEN_2713; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2715 = 8'h9b == io_state_in_10 ? 8'he8 : _GEN_2714; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2716 = 8'h9c == io_state_in_10 ? 8'h1c : _GEN_2715; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2717 = 8'h9d == io_state_in_10 ? 8'h75 : _GEN_2716; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2718 = 8'h9e == io_state_in_10 ? 8'hdf : _GEN_2717; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2719 = 8'h9f == io_state_in_10 ? 8'h6e : _GEN_2718; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2720 = 8'ha0 == io_state_in_10 ? 8'h47 : _GEN_2719; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2721 = 8'ha1 == io_state_in_10 ? 8'hf1 : _GEN_2720; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2722 = 8'ha2 == io_state_in_10 ? 8'h1a : _GEN_2721; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2723 = 8'ha3 == io_state_in_10 ? 8'h71 : _GEN_2722; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2724 = 8'ha4 == io_state_in_10 ? 8'h1d : _GEN_2723; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2725 = 8'ha5 == io_state_in_10 ? 8'h29 : _GEN_2724; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2726 = 8'ha6 == io_state_in_10 ? 8'hc5 : _GEN_2725; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2727 = 8'ha7 == io_state_in_10 ? 8'h89 : _GEN_2726; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2728 = 8'ha8 == io_state_in_10 ? 8'h6f : _GEN_2727; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2729 = 8'ha9 == io_state_in_10 ? 8'hb7 : _GEN_2728; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2730 = 8'haa == io_state_in_10 ? 8'h62 : _GEN_2729; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2731 = 8'hab == io_state_in_10 ? 8'he : _GEN_2730; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2732 = 8'hac == io_state_in_10 ? 8'haa : _GEN_2731; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2733 = 8'had == io_state_in_10 ? 8'h18 : _GEN_2732; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2734 = 8'hae == io_state_in_10 ? 8'hbe : _GEN_2733; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2735 = 8'haf == io_state_in_10 ? 8'h1b : _GEN_2734; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2736 = 8'hb0 == io_state_in_10 ? 8'hfc : _GEN_2735; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2737 = 8'hb1 == io_state_in_10 ? 8'h56 : _GEN_2736; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2738 = 8'hb2 == io_state_in_10 ? 8'h3e : _GEN_2737; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2739 = 8'hb3 == io_state_in_10 ? 8'h4b : _GEN_2738; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2740 = 8'hb4 == io_state_in_10 ? 8'hc6 : _GEN_2739; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2741 = 8'hb5 == io_state_in_10 ? 8'hd2 : _GEN_2740; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2742 = 8'hb6 == io_state_in_10 ? 8'h79 : _GEN_2741; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2743 = 8'hb7 == io_state_in_10 ? 8'h20 : _GEN_2742; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2744 = 8'hb8 == io_state_in_10 ? 8'h9a : _GEN_2743; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2745 = 8'hb9 == io_state_in_10 ? 8'hdb : _GEN_2744; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2746 = 8'hba == io_state_in_10 ? 8'hc0 : _GEN_2745; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2747 = 8'hbb == io_state_in_10 ? 8'hfe : _GEN_2746; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2748 = 8'hbc == io_state_in_10 ? 8'h78 : _GEN_2747; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2749 = 8'hbd == io_state_in_10 ? 8'hcd : _GEN_2748; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2750 = 8'hbe == io_state_in_10 ? 8'h5a : _GEN_2749; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2751 = 8'hbf == io_state_in_10 ? 8'hf4 : _GEN_2750; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2752 = 8'hc0 == io_state_in_10 ? 8'h1f : _GEN_2751; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2753 = 8'hc1 == io_state_in_10 ? 8'hdd : _GEN_2752; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2754 = 8'hc2 == io_state_in_10 ? 8'ha8 : _GEN_2753; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2755 = 8'hc3 == io_state_in_10 ? 8'h33 : _GEN_2754; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2756 = 8'hc4 == io_state_in_10 ? 8'h88 : _GEN_2755; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2757 = 8'hc5 == io_state_in_10 ? 8'h7 : _GEN_2756; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2758 = 8'hc6 == io_state_in_10 ? 8'hc7 : _GEN_2757; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2759 = 8'hc7 == io_state_in_10 ? 8'h31 : _GEN_2758; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2760 = 8'hc8 == io_state_in_10 ? 8'hb1 : _GEN_2759; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2761 = 8'hc9 == io_state_in_10 ? 8'h12 : _GEN_2760; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2762 = 8'hca == io_state_in_10 ? 8'h10 : _GEN_2761; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2763 = 8'hcb == io_state_in_10 ? 8'h59 : _GEN_2762; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2764 = 8'hcc == io_state_in_10 ? 8'h27 : _GEN_2763; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2765 = 8'hcd == io_state_in_10 ? 8'h80 : _GEN_2764; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2766 = 8'hce == io_state_in_10 ? 8'hec : _GEN_2765; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2767 = 8'hcf == io_state_in_10 ? 8'h5f : _GEN_2766; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2768 = 8'hd0 == io_state_in_10 ? 8'h60 : _GEN_2767; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2769 = 8'hd1 == io_state_in_10 ? 8'h51 : _GEN_2768; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2770 = 8'hd2 == io_state_in_10 ? 8'h7f : _GEN_2769; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2771 = 8'hd3 == io_state_in_10 ? 8'ha9 : _GEN_2770; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2772 = 8'hd4 == io_state_in_10 ? 8'h19 : _GEN_2771; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2773 = 8'hd5 == io_state_in_10 ? 8'hb5 : _GEN_2772; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2774 = 8'hd6 == io_state_in_10 ? 8'h4a : _GEN_2773; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2775 = 8'hd7 == io_state_in_10 ? 8'hd : _GEN_2774; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2776 = 8'hd8 == io_state_in_10 ? 8'h2d : _GEN_2775; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2777 = 8'hd9 == io_state_in_10 ? 8'he5 : _GEN_2776; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2778 = 8'hda == io_state_in_10 ? 8'h7a : _GEN_2777; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2779 = 8'hdb == io_state_in_10 ? 8'h9f : _GEN_2778; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2780 = 8'hdc == io_state_in_10 ? 8'h93 : _GEN_2779; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2781 = 8'hdd == io_state_in_10 ? 8'hc9 : _GEN_2780; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2782 = 8'hde == io_state_in_10 ? 8'h9c : _GEN_2781; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2783 = 8'hdf == io_state_in_10 ? 8'hef : _GEN_2782; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2784 = 8'he0 == io_state_in_10 ? 8'ha0 : _GEN_2783; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2785 = 8'he1 == io_state_in_10 ? 8'he0 : _GEN_2784; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2786 = 8'he2 == io_state_in_10 ? 8'h3b : _GEN_2785; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2787 = 8'he3 == io_state_in_10 ? 8'h4d : _GEN_2786; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2788 = 8'he4 == io_state_in_10 ? 8'hae : _GEN_2787; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2789 = 8'he5 == io_state_in_10 ? 8'h2a : _GEN_2788; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2790 = 8'he6 == io_state_in_10 ? 8'hf5 : _GEN_2789; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2791 = 8'he7 == io_state_in_10 ? 8'hb0 : _GEN_2790; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2792 = 8'he8 == io_state_in_10 ? 8'hc8 : _GEN_2791; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2793 = 8'he9 == io_state_in_10 ? 8'heb : _GEN_2792; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2794 = 8'hea == io_state_in_10 ? 8'hbb : _GEN_2793; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2795 = 8'heb == io_state_in_10 ? 8'h3c : _GEN_2794; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2796 = 8'hec == io_state_in_10 ? 8'h83 : _GEN_2795; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2797 = 8'hed == io_state_in_10 ? 8'h53 : _GEN_2796; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2798 = 8'hee == io_state_in_10 ? 8'h99 : _GEN_2797; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2799 = 8'hef == io_state_in_10 ? 8'h61 : _GEN_2798; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2800 = 8'hf0 == io_state_in_10 ? 8'h17 : _GEN_2799; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2801 = 8'hf1 == io_state_in_10 ? 8'h2b : _GEN_2800; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2802 = 8'hf2 == io_state_in_10 ? 8'h4 : _GEN_2801; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2803 = 8'hf3 == io_state_in_10 ? 8'h7e : _GEN_2802; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2804 = 8'hf4 == io_state_in_10 ? 8'hba : _GEN_2803; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2805 = 8'hf5 == io_state_in_10 ? 8'h77 : _GEN_2804; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2806 = 8'hf6 == io_state_in_10 ? 8'hd6 : _GEN_2805; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2807 = 8'hf7 == io_state_in_10 ? 8'h26 : _GEN_2806; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2808 = 8'hf8 == io_state_in_10 ? 8'he1 : _GEN_2807; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2809 = 8'hf9 == io_state_in_10 ? 8'h69 : _GEN_2808; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2810 = 8'hfa == io_state_in_10 ? 8'h14 : _GEN_2809; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2811 = 8'hfb == io_state_in_10 ? 8'h63 : _GEN_2810; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2812 = 8'hfc == io_state_in_10 ? 8'h55 : _GEN_2811; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2813 = 8'hfd == io_state_in_10 ? 8'h21 : _GEN_2812; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2814 = 8'hfe == io_state_in_10 ? 8'hc : _GEN_2813; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2817 = 8'h1 == io_state_in_11 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2818 = 8'h2 == io_state_in_11 ? 8'h6a : _GEN_2817; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2819 = 8'h3 == io_state_in_11 ? 8'hd5 : _GEN_2818; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2820 = 8'h4 == io_state_in_11 ? 8'h30 : _GEN_2819; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2821 = 8'h5 == io_state_in_11 ? 8'h36 : _GEN_2820; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2822 = 8'h6 == io_state_in_11 ? 8'ha5 : _GEN_2821; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2823 = 8'h7 == io_state_in_11 ? 8'h38 : _GEN_2822; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2824 = 8'h8 == io_state_in_11 ? 8'hbf : _GEN_2823; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2825 = 8'h9 == io_state_in_11 ? 8'h40 : _GEN_2824; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2826 = 8'ha == io_state_in_11 ? 8'ha3 : _GEN_2825; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2827 = 8'hb == io_state_in_11 ? 8'h9e : _GEN_2826; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2828 = 8'hc == io_state_in_11 ? 8'h81 : _GEN_2827; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2829 = 8'hd == io_state_in_11 ? 8'hf3 : _GEN_2828; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2830 = 8'he == io_state_in_11 ? 8'hd7 : _GEN_2829; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2831 = 8'hf == io_state_in_11 ? 8'hfb : _GEN_2830; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2832 = 8'h10 == io_state_in_11 ? 8'h7c : _GEN_2831; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2833 = 8'h11 == io_state_in_11 ? 8'he3 : _GEN_2832; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2834 = 8'h12 == io_state_in_11 ? 8'h39 : _GEN_2833; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2835 = 8'h13 == io_state_in_11 ? 8'h82 : _GEN_2834; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2836 = 8'h14 == io_state_in_11 ? 8'h9b : _GEN_2835; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2837 = 8'h15 == io_state_in_11 ? 8'h2f : _GEN_2836; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2838 = 8'h16 == io_state_in_11 ? 8'hff : _GEN_2837; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2839 = 8'h17 == io_state_in_11 ? 8'h87 : _GEN_2838; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2840 = 8'h18 == io_state_in_11 ? 8'h34 : _GEN_2839; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2841 = 8'h19 == io_state_in_11 ? 8'h8e : _GEN_2840; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2842 = 8'h1a == io_state_in_11 ? 8'h43 : _GEN_2841; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2843 = 8'h1b == io_state_in_11 ? 8'h44 : _GEN_2842; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2844 = 8'h1c == io_state_in_11 ? 8'hc4 : _GEN_2843; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2845 = 8'h1d == io_state_in_11 ? 8'hde : _GEN_2844; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2846 = 8'h1e == io_state_in_11 ? 8'he9 : _GEN_2845; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2847 = 8'h1f == io_state_in_11 ? 8'hcb : _GEN_2846; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2848 = 8'h20 == io_state_in_11 ? 8'h54 : _GEN_2847; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2849 = 8'h21 == io_state_in_11 ? 8'h7b : _GEN_2848; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2850 = 8'h22 == io_state_in_11 ? 8'h94 : _GEN_2849; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2851 = 8'h23 == io_state_in_11 ? 8'h32 : _GEN_2850; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2852 = 8'h24 == io_state_in_11 ? 8'ha6 : _GEN_2851; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2853 = 8'h25 == io_state_in_11 ? 8'hc2 : _GEN_2852; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2854 = 8'h26 == io_state_in_11 ? 8'h23 : _GEN_2853; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2855 = 8'h27 == io_state_in_11 ? 8'h3d : _GEN_2854; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2856 = 8'h28 == io_state_in_11 ? 8'hee : _GEN_2855; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2857 = 8'h29 == io_state_in_11 ? 8'h4c : _GEN_2856; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2858 = 8'h2a == io_state_in_11 ? 8'h95 : _GEN_2857; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2859 = 8'h2b == io_state_in_11 ? 8'hb : _GEN_2858; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2860 = 8'h2c == io_state_in_11 ? 8'h42 : _GEN_2859; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2861 = 8'h2d == io_state_in_11 ? 8'hfa : _GEN_2860; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2862 = 8'h2e == io_state_in_11 ? 8'hc3 : _GEN_2861; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2863 = 8'h2f == io_state_in_11 ? 8'h4e : _GEN_2862; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2864 = 8'h30 == io_state_in_11 ? 8'h8 : _GEN_2863; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2865 = 8'h31 == io_state_in_11 ? 8'h2e : _GEN_2864; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2866 = 8'h32 == io_state_in_11 ? 8'ha1 : _GEN_2865; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2867 = 8'h33 == io_state_in_11 ? 8'h66 : _GEN_2866; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2868 = 8'h34 == io_state_in_11 ? 8'h28 : _GEN_2867; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2869 = 8'h35 == io_state_in_11 ? 8'hd9 : _GEN_2868; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2870 = 8'h36 == io_state_in_11 ? 8'h24 : _GEN_2869; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2871 = 8'h37 == io_state_in_11 ? 8'hb2 : _GEN_2870; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2872 = 8'h38 == io_state_in_11 ? 8'h76 : _GEN_2871; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2873 = 8'h39 == io_state_in_11 ? 8'h5b : _GEN_2872; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2874 = 8'h3a == io_state_in_11 ? 8'ha2 : _GEN_2873; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2875 = 8'h3b == io_state_in_11 ? 8'h49 : _GEN_2874; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2876 = 8'h3c == io_state_in_11 ? 8'h6d : _GEN_2875; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2877 = 8'h3d == io_state_in_11 ? 8'h8b : _GEN_2876; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2878 = 8'h3e == io_state_in_11 ? 8'hd1 : _GEN_2877; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2879 = 8'h3f == io_state_in_11 ? 8'h25 : _GEN_2878; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2880 = 8'h40 == io_state_in_11 ? 8'h72 : _GEN_2879; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2881 = 8'h41 == io_state_in_11 ? 8'hf8 : _GEN_2880; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2882 = 8'h42 == io_state_in_11 ? 8'hf6 : _GEN_2881; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2883 = 8'h43 == io_state_in_11 ? 8'h64 : _GEN_2882; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2884 = 8'h44 == io_state_in_11 ? 8'h86 : _GEN_2883; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2885 = 8'h45 == io_state_in_11 ? 8'h68 : _GEN_2884; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2886 = 8'h46 == io_state_in_11 ? 8'h98 : _GEN_2885; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2887 = 8'h47 == io_state_in_11 ? 8'h16 : _GEN_2886; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2888 = 8'h48 == io_state_in_11 ? 8'hd4 : _GEN_2887; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2889 = 8'h49 == io_state_in_11 ? 8'ha4 : _GEN_2888; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2890 = 8'h4a == io_state_in_11 ? 8'h5c : _GEN_2889; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2891 = 8'h4b == io_state_in_11 ? 8'hcc : _GEN_2890; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2892 = 8'h4c == io_state_in_11 ? 8'h5d : _GEN_2891; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2893 = 8'h4d == io_state_in_11 ? 8'h65 : _GEN_2892; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2894 = 8'h4e == io_state_in_11 ? 8'hb6 : _GEN_2893; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2895 = 8'h4f == io_state_in_11 ? 8'h92 : _GEN_2894; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2896 = 8'h50 == io_state_in_11 ? 8'h6c : _GEN_2895; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2897 = 8'h51 == io_state_in_11 ? 8'h70 : _GEN_2896; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2898 = 8'h52 == io_state_in_11 ? 8'h48 : _GEN_2897; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2899 = 8'h53 == io_state_in_11 ? 8'h50 : _GEN_2898; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2900 = 8'h54 == io_state_in_11 ? 8'hfd : _GEN_2899; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2901 = 8'h55 == io_state_in_11 ? 8'hed : _GEN_2900; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2902 = 8'h56 == io_state_in_11 ? 8'hb9 : _GEN_2901; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2903 = 8'h57 == io_state_in_11 ? 8'hda : _GEN_2902; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2904 = 8'h58 == io_state_in_11 ? 8'h5e : _GEN_2903; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2905 = 8'h59 == io_state_in_11 ? 8'h15 : _GEN_2904; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2906 = 8'h5a == io_state_in_11 ? 8'h46 : _GEN_2905; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2907 = 8'h5b == io_state_in_11 ? 8'h57 : _GEN_2906; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2908 = 8'h5c == io_state_in_11 ? 8'ha7 : _GEN_2907; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2909 = 8'h5d == io_state_in_11 ? 8'h8d : _GEN_2908; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2910 = 8'h5e == io_state_in_11 ? 8'h9d : _GEN_2909; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2911 = 8'h5f == io_state_in_11 ? 8'h84 : _GEN_2910; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2912 = 8'h60 == io_state_in_11 ? 8'h90 : _GEN_2911; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2913 = 8'h61 == io_state_in_11 ? 8'hd8 : _GEN_2912; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2914 = 8'h62 == io_state_in_11 ? 8'hab : _GEN_2913; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2915 = 8'h63 == io_state_in_11 ? 8'h0 : _GEN_2914; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2916 = 8'h64 == io_state_in_11 ? 8'h8c : _GEN_2915; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2917 = 8'h65 == io_state_in_11 ? 8'hbc : _GEN_2916; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2918 = 8'h66 == io_state_in_11 ? 8'hd3 : _GEN_2917; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2919 = 8'h67 == io_state_in_11 ? 8'ha : _GEN_2918; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2920 = 8'h68 == io_state_in_11 ? 8'hf7 : _GEN_2919; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2921 = 8'h69 == io_state_in_11 ? 8'he4 : _GEN_2920; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2922 = 8'h6a == io_state_in_11 ? 8'h58 : _GEN_2921; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2923 = 8'h6b == io_state_in_11 ? 8'h5 : _GEN_2922; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2924 = 8'h6c == io_state_in_11 ? 8'hb8 : _GEN_2923; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2925 = 8'h6d == io_state_in_11 ? 8'hb3 : _GEN_2924; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2926 = 8'h6e == io_state_in_11 ? 8'h45 : _GEN_2925; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2927 = 8'h6f == io_state_in_11 ? 8'h6 : _GEN_2926; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2928 = 8'h70 == io_state_in_11 ? 8'hd0 : _GEN_2927; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2929 = 8'h71 == io_state_in_11 ? 8'h2c : _GEN_2928; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2930 = 8'h72 == io_state_in_11 ? 8'h1e : _GEN_2929; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2931 = 8'h73 == io_state_in_11 ? 8'h8f : _GEN_2930; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2932 = 8'h74 == io_state_in_11 ? 8'hca : _GEN_2931; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2933 = 8'h75 == io_state_in_11 ? 8'h3f : _GEN_2932; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2934 = 8'h76 == io_state_in_11 ? 8'hf : _GEN_2933; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2935 = 8'h77 == io_state_in_11 ? 8'h2 : _GEN_2934; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2936 = 8'h78 == io_state_in_11 ? 8'hc1 : _GEN_2935; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2937 = 8'h79 == io_state_in_11 ? 8'haf : _GEN_2936; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2938 = 8'h7a == io_state_in_11 ? 8'hbd : _GEN_2937; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2939 = 8'h7b == io_state_in_11 ? 8'h3 : _GEN_2938; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2940 = 8'h7c == io_state_in_11 ? 8'h1 : _GEN_2939; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2941 = 8'h7d == io_state_in_11 ? 8'h13 : _GEN_2940; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2942 = 8'h7e == io_state_in_11 ? 8'h8a : _GEN_2941; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2943 = 8'h7f == io_state_in_11 ? 8'h6b : _GEN_2942; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2944 = 8'h80 == io_state_in_11 ? 8'h3a : _GEN_2943; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2945 = 8'h81 == io_state_in_11 ? 8'h91 : _GEN_2944; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2946 = 8'h82 == io_state_in_11 ? 8'h11 : _GEN_2945; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2947 = 8'h83 == io_state_in_11 ? 8'h41 : _GEN_2946; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2948 = 8'h84 == io_state_in_11 ? 8'h4f : _GEN_2947; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2949 = 8'h85 == io_state_in_11 ? 8'h67 : _GEN_2948; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2950 = 8'h86 == io_state_in_11 ? 8'hdc : _GEN_2949; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2951 = 8'h87 == io_state_in_11 ? 8'hea : _GEN_2950; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2952 = 8'h88 == io_state_in_11 ? 8'h97 : _GEN_2951; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2953 = 8'h89 == io_state_in_11 ? 8'hf2 : _GEN_2952; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2954 = 8'h8a == io_state_in_11 ? 8'hcf : _GEN_2953; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2955 = 8'h8b == io_state_in_11 ? 8'hce : _GEN_2954; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2956 = 8'h8c == io_state_in_11 ? 8'hf0 : _GEN_2955; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2957 = 8'h8d == io_state_in_11 ? 8'hb4 : _GEN_2956; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2958 = 8'h8e == io_state_in_11 ? 8'he6 : _GEN_2957; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2959 = 8'h8f == io_state_in_11 ? 8'h73 : _GEN_2958; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2960 = 8'h90 == io_state_in_11 ? 8'h96 : _GEN_2959; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2961 = 8'h91 == io_state_in_11 ? 8'hac : _GEN_2960; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2962 = 8'h92 == io_state_in_11 ? 8'h74 : _GEN_2961; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2963 = 8'h93 == io_state_in_11 ? 8'h22 : _GEN_2962; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2964 = 8'h94 == io_state_in_11 ? 8'he7 : _GEN_2963; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2965 = 8'h95 == io_state_in_11 ? 8'had : _GEN_2964; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2966 = 8'h96 == io_state_in_11 ? 8'h35 : _GEN_2965; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2967 = 8'h97 == io_state_in_11 ? 8'h85 : _GEN_2966; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2968 = 8'h98 == io_state_in_11 ? 8'he2 : _GEN_2967; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2969 = 8'h99 == io_state_in_11 ? 8'hf9 : _GEN_2968; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2970 = 8'h9a == io_state_in_11 ? 8'h37 : _GEN_2969; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2971 = 8'h9b == io_state_in_11 ? 8'he8 : _GEN_2970; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2972 = 8'h9c == io_state_in_11 ? 8'h1c : _GEN_2971; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2973 = 8'h9d == io_state_in_11 ? 8'h75 : _GEN_2972; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2974 = 8'h9e == io_state_in_11 ? 8'hdf : _GEN_2973; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2975 = 8'h9f == io_state_in_11 ? 8'h6e : _GEN_2974; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2976 = 8'ha0 == io_state_in_11 ? 8'h47 : _GEN_2975; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2977 = 8'ha1 == io_state_in_11 ? 8'hf1 : _GEN_2976; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2978 = 8'ha2 == io_state_in_11 ? 8'h1a : _GEN_2977; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2979 = 8'ha3 == io_state_in_11 ? 8'h71 : _GEN_2978; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2980 = 8'ha4 == io_state_in_11 ? 8'h1d : _GEN_2979; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2981 = 8'ha5 == io_state_in_11 ? 8'h29 : _GEN_2980; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2982 = 8'ha6 == io_state_in_11 ? 8'hc5 : _GEN_2981; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2983 = 8'ha7 == io_state_in_11 ? 8'h89 : _GEN_2982; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2984 = 8'ha8 == io_state_in_11 ? 8'h6f : _GEN_2983; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2985 = 8'ha9 == io_state_in_11 ? 8'hb7 : _GEN_2984; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2986 = 8'haa == io_state_in_11 ? 8'h62 : _GEN_2985; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2987 = 8'hab == io_state_in_11 ? 8'he : _GEN_2986; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2988 = 8'hac == io_state_in_11 ? 8'haa : _GEN_2987; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2989 = 8'had == io_state_in_11 ? 8'h18 : _GEN_2988; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2990 = 8'hae == io_state_in_11 ? 8'hbe : _GEN_2989; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2991 = 8'haf == io_state_in_11 ? 8'h1b : _GEN_2990; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2992 = 8'hb0 == io_state_in_11 ? 8'hfc : _GEN_2991; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2993 = 8'hb1 == io_state_in_11 ? 8'h56 : _GEN_2992; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2994 = 8'hb2 == io_state_in_11 ? 8'h3e : _GEN_2993; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2995 = 8'hb3 == io_state_in_11 ? 8'h4b : _GEN_2994; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2996 = 8'hb4 == io_state_in_11 ? 8'hc6 : _GEN_2995; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2997 = 8'hb5 == io_state_in_11 ? 8'hd2 : _GEN_2996; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2998 = 8'hb6 == io_state_in_11 ? 8'h79 : _GEN_2997; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_2999 = 8'hb7 == io_state_in_11 ? 8'h20 : _GEN_2998; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3000 = 8'hb8 == io_state_in_11 ? 8'h9a : _GEN_2999; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3001 = 8'hb9 == io_state_in_11 ? 8'hdb : _GEN_3000; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3002 = 8'hba == io_state_in_11 ? 8'hc0 : _GEN_3001; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3003 = 8'hbb == io_state_in_11 ? 8'hfe : _GEN_3002; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3004 = 8'hbc == io_state_in_11 ? 8'h78 : _GEN_3003; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3005 = 8'hbd == io_state_in_11 ? 8'hcd : _GEN_3004; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3006 = 8'hbe == io_state_in_11 ? 8'h5a : _GEN_3005; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3007 = 8'hbf == io_state_in_11 ? 8'hf4 : _GEN_3006; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3008 = 8'hc0 == io_state_in_11 ? 8'h1f : _GEN_3007; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3009 = 8'hc1 == io_state_in_11 ? 8'hdd : _GEN_3008; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3010 = 8'hc2 == io_state_in_11 ? 8'ha8 : _GEN_3009; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3011 = 8'hc3 == io_state_in_11 ? 8'h33 : _GEN_3010; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3012 = 8'hc4 == io_state_in_11 ? 8'h88 : _GEN_3011; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3013 = 8'hc5 == io_state_in_11 ? 8'h7 : _GEN_3012; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3014 = 8'hc6 == io_state_in_11 ? 8'hc7 : _GEN_3013; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3015 = 8'hc7 == io_state_in_11 ? 8'h31 : _GEN_3014; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3016 = 8'hc8 == io_state_in_11 ? 8'hb1 : _GEN_3015; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3017 = 8'hc9 == io_state_in_11 ? 8'h12 : _GEN_3016; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3018 = 8'hca == io_state_in_11 ? 8'h10 : _GEN_3017; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3019 = 8'hcb == io_state_in_11 ? 8'h59 : _GEN_3018; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3020 = 8'hcc == io_state_in_11 ? 8'h27 : _GEN_3019; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3021 = 8'hcd == io_state_in_11 ? 8'h80 : _GEN_3020; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3022 = 8'hce == io_state_in_11 ? 8'hec : _GEN_3021; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3023 = 8'hcf == io_state_in_11 ? 8'h5f : _GEN_3022; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3024 = 8'hd0 == io_state_in_11 ? 8'h60 : _GEN_3023; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3025 = 8'hd1 == io_state_in_11 ? 8'h51 : _GEN_3024; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3026 = 8'hd2 == io_state_in_11 ? 8'h7f : _GEN_3025; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3027 = 8'hd3 == io_state_in_11 ? 8'ha9 : _GEN_3026; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3028 = 8'hd4 == io_state_in_11 ? 8'h19 : _GEN_3027; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3029 = 8'hd5 == io_state_in_11 ? 8'hb5 : _GEN_3028; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3030 = 8'hd6 == io_state_in_11 ? 8'h4a : _GEN_3029; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3031 = 8'hd7 == io_state_in_11 ? 8'hd : _GEN_3030; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3032 = 8'hd8 == io_state_in_11 ? 8'h2d : _GEN_3031; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3033 = 8'hd9 == io_state_in_11 ? 8'he5 : _GEN_3032; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3034 = 8'hda == io_state_in_11 ? 8'h7a : _GEN_3033; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3035 = 8'hdb == io_state_in_11 ? 8'h9f : _GEN_3034; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3036 = 8'hdc == io_state_in_11 ? 8'h93 : _GEN_3035; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3037 = 8'hdd == io_state_in_11 ? 8'hc9 : _GEN_3036; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3038 = 8'hde == io_state_in_11 ? 8'h9c : _GEN_3037; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3039 = 8'hdf == io_state_in_11 ? 8'hef : _GEN_3038; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3040 = 8'he0 == io_state_in_11 ? 8'ha0 : _GEN_3039; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3041 = 8'he1 == io_state_in_11 ? 8'he0 : _GEN_3040; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3042 = 8'he2 == io_state_in_11 ? 8'h3b : _GEN_3041; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3043 = 8'he3 == io_state_in_11 ? 8'h4d : _GEN_3042; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3044 = 8'he4 == io_state_in_11 ? 8'hae : _GEN_3043; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3045 = 8'he5 == io_state_in_11 ? 8'h2a : _GEN_3044; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3046 = 8'he6 == io_state_in_11 ? 8'hf5 : _GEN_3045; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3047 = 8'he7 == io_state_in_11 ? 8'hb0 : _GEN_3046; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3048 = 8'he8 == io_state_in_11 ? 8'hc8 : _GEN_3047; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3049 = 8'he9 == io_state_in_11 ? 8'heb : _GEN_3048; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3050 = 8'hea == io_state_in_11 ? 8'hbb : _GEN_3049; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3051 = 8'heb == io_state_in_11 ? 8'h3c : _GEN_3050; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3052 = 8'hec == io_state_in_11 ? 8'h83 : _GEN_3051; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3053 = 8'hed == io_state_in_11 ? 8'h53 : _GEN_3052; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3054 = 8'hee == io_state_in_11 ? 8'h99 : _GEN_3053; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3055 = 8'hef == io_state_in_11 ? 8'h61 : _GEN_3054; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3056 = 8'hf0 == io_state_in_11 ? 8'h17 : _GEN_3055; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3057 = 8'hf1 == io_state_in_11 ? 8'h2b : _GEN_3056; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3058 = 8'hf2 == io_state_in_11 ? 8'h4 : _GEN_3057; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3059 = 8'hf3 == io_state_in_11 ? 8'h7e : _GEN_3058; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3060 = 8'hf4 == io_state_in_11 ? 8'hba : _GEN_3059; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3061 = 8'hf5 == io_state_in_11 ? 8'h77 : _GEN_3060; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3062 = 8'hf6 == io_state_in_11 ? 8'hd6 : _GEN_3061; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3063 = 8'hf7 == io_state_in_11 ? 8'h26 : _GEN_3062; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3064 = 8'hf8 == io_state_in_11 ? 8'he1 : _GEN_3063; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3065 = 8'hf9 == io_state_in_11 ? 8'h69 : _GEN_3064; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3066 = 8'hfa == io_state_in_11 ? 8'h14 : _GEN_3065; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3067 = 8'hfb == io_state_in_11 ? 8'h63 : _GEN_3066; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3068 = 8'hfc == io_state_in_11 ? 8'h55 : _GEN_3067; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3069 = 8'hfd == io_state_in_11 ? 8'h21 : _GEN_3068; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3070 = 8'hfe == io_state_in_11 ? 8'hc : _GEN_3069; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3073 = 8'h1 == io_state_in_12 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3074 = 8'h2 == io_state_in_12 ? 8'h6a : _GEN_3073; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3075 = 8'h3 == io_state_in_12 ? 8'hd5 : _GEN_3074; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3076 = 8'h4 == io_state_in_12 ? 8'h30 : _GEN_3075; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3077 = 8'h5 == io_state_in_12 ? 8'h36 : _GEN_3076; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3078 = 8'h6 == io_state_in_12 ? 8'ha5 : _GEN_3077; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3079 = 8'h7 == io_state_in_12 ? 8'h38 : _GEN_3078; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3080 = 8'h8 == io_state_in_12 ? 8'hbf : _GEN_3079; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3081 = 8'h9 == io_state_in_12 ? 8'h40 : _GEN_3080; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3082 = 8'ha == io_state_in_12 ? 8'ha3 : _GEN_3081; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3083 = 8'hb == io_state_in_12 ? 8'h9e : _GEN_3082; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3084 = 8'hc == io_state_in_12 ? 8'h81 : _GEN_3083; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3085 = 8'hd == io_state_in_12 ? 8'hf3 : _GEN_3084; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3086 = 8'he == io_state_in_12 ? 8'hd7 : _GEN_3085; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3087 = 8'hf == io_state_in_12 ? 8'hfb : _GEN_3086; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3088 = 8'h10 == io_state_in_12 ? 8'h7c : _GEN_3087; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3089 = 8'h11 == io_state_in_12 ? 8'he3 : _GEN_3088; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3090 = 8'h12 == io_state_in_12 ? 8'h39 : _GEN_3089; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3091 = 8'h13 == io_state_in_12 ? 8'h82 : _GEN_3090; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3092 = 8'h14 == io_state_in_12 ? 8'h9b : _GEN_3091; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3093 = 8'h15 == io_state_in_12 ? 8'h2f : _GEN_3092; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3094 = 8'h16 == io_state_in_12 ? 8'hff : _GEN_3093; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3095 = 8'h17 == io_state_in_12 ? 8'h87 : _GEN_3094; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3096 = 8'h18 == io_state_in_12 ? 8'h34 : _GEN_3095; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3097 = 8'h19 == io_state_in_12 ? 8'h8e : _GEN_3096; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3098 = 8'h1a == io_state_in_12 ? 8'h43 : _GEN_3097; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3099 = 8'h1b == io_state_in_12 ? 8'h44 : _GEN_3098; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3100 = 8'h1c == io_state_in_12 ? 8'hc4 : _GEN_3099; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3101 = 8'h1d == io_state_in_12 ? 8'hde : _GEN_3100; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3102 = 8'h1e == io_state_in_12 ? 8'he9 : _GEN_3101; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3103 = 8'h1f == io_state_in_12 ? 8'hcb : _GEN_3102; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3104 = 8'h20 == io_state_in_12 ? 8'h54 : _GEN_3103; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3105 = 8'h21 == io_state_in_12 ? 8'h7b : _GEN_3104; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3106 = 8'h22 == io_state_in_12 ? 8'h94 : _GEN_3105; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3107 = 8'h23 == io_state_in_12 ? 8'h32 : _GEN_3106; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3108 = 8'h24 == io_state_in_12 ? 8'ha6 : _GEN_3107; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3109 = 8'h25 == io_state_in_12 ? 8'hc2 : _GEN_3108; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3110 = 8'h26 == io_state_in_12 ? 8'h23 : _GEN_3109; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3111 = 8'h27 == io_state_in_12 ? 8'h3d : _GEN_3110; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3112 = 8'h28 == io_state_in_12 ? 8'hee : _GEN_3111; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3113 = 8'h29 == io_state_in_12 ? 8'h4c : _GEN_3112; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3114 = 8'h2a == io_state_in_12 ? 8'h95 : _GEN_3113; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3115 = 8'h2b == io_state_in_12 ? 8'hb : _GEN_3114; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3116 = 8'h2c == io_state_in_12 ? 8'h42 : _GEN_3115; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3117 = 8'h2d == io_state_in_12 ? 8'hfa : _GEN_3116; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3118 = 8'h2e == io_state_in_12 ? 8'hc3 : _GEN_3117; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3119 = 8'h2f == io_state_in_12 ? 8'h4e : _GEN_3118; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3120 = 8'h30 == io_state_in_12 ? 8'h8 : _GEN_3119; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3121 = 8'h31 == io_state_in_12 ? 8'h2e : _GEN_3120; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3122 = 8'h32 == io_state_in_12 ? 8'ha1 : _GEN_3121; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3123 = 8'h33 == io_state_in_12 ? 8'h66 : _GEN_3122; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3124 = 8'h34 == io_state_in_12 ? 8'h28 : _GEN_3123; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3125 = 8'h35 == io_state_in_12 ? 8'hd9 : _GEN_3124; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3126 = 8'h36 == io_state_in_12 ? 8'h24 : _GEN_3125; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3127 = 8'h37 == io_state_in_12 ? 8'hb2 : _GEN_3126; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3128 = 8'h38 == io_state_in_12 ? 8'h76 : _GEN_3127; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3129 = 8'h39 == io_state_in_12 ? 8'h5b : _GEN_3128; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3130 = 8'h3a == io_state_in_12 ? 8'ha2 : _GEN_3129; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3131 = 8'h3b == io_state_in_12 ? 8'h49 : _GEN_3130; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3132 = 8'h3c == io_state_in_12 ? 8'h6d : _GEN_3131; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3133 = 8'h3d == io_state_in_12 ? 8'h8b : _GEN_3132; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3134 = 8'h3e == io_state_in_12 ? 8'hd1 : _GEN_3133; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3135 = 8'h3f == io_state_in_12 ? 8'h25 : _GEN_3134; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3136 = 8'h40 == io_state_in_12 ? 8'h72 : _GEN_3135; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3137 = 8'h41 == io_state_in_12 ? 8'hf8 : _GEN_3136; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3138 = 8'h42 == io_state_in_12 ? 8'hf6 : _GEN_3137; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3139 = 8'h43 == io_state_in_12 ? 8'h64 : _GEN_3138; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3140 = 8'h44 == io_state_in_12 ? 8'h86 : _GEN_3139; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3141 = 8'h45 == io_state_in_12 ? 8'h68 : _GEN_3140; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3142 = 8'h46 == io_state_in_12 ? 8'h98 : _GEN_3141; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3143 = 8'h47 == io_state_in_12 ? 8'h16 : _GEN_3142; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3144 = 8'h48 == io_state_in_12 ? 8'hd4 : _GEN_3143; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3145 = 8'h49 == io_state_in_12 ? 8'ha4 : _GEN_3144; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3146 = 8'h4a == io_state_in_12 ? 8'h5c : _GEN_3145; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3147 = 8'h4b == io_state_in_12 ? 8'hcc : _GEN_3146; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3148 = 8'h4c == io_state_in_12 ? 8'h5d : _GEN_3147; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3149 = 8'h4d == io_state_in_12 ? 8'h65 : _GEN_3148; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3150 = 8'h4e == io_state_in_12 ? 8'hb6 : _GEN_3149; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3151 = 8'h4f == io_state_in_12 ? 8'h92 : _GEN_3150; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3152 = 8'h50 == io_state_in_12 ? 8'h6c : _GEN_3151; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3153 = 8'h51 == io_state_in_12 ? 8'h70 : _GEN_3152; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3154 = 8'h52 == io_state_in_12 ? 8'h48 : _GEN_3153; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3155 = 8'h53 == io_state_in_12 ? 8'h50 : _GEN_3154; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3156 = 8'h54 == io_state_in_12 ? 8'hfd : _GEN_3155; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3157 = 8'h55 == io_state_in_12 ? 8'hed : _GEN_3156; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3158 = 8'h56 == io_state_in_12 ? 8'hb9 : _GEN_3157; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3159 = 8'h57 == io_state_in_12 ? 8'hda : _GEN_3158; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3160 = 8'h58 == io_state_in_12 ? 8'h5e : _GEN_3159; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3161 = 8'h59 == io_state_in_12 ? 8'h15 : _GEN_3160; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3162 = 8'h5a == io_state_in_12 ? 8'h46 : _GEN_3161; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3163 = 8'h5b == io_state_in_12 ? 8'h57 : _GEN_3162; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3164 = 8'h5c == io_state_in_12 ? 8'ha7 : _GEN_3163; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3165 = 8'h5d == io_state_in_12 ? 8'h8d : _GEN_3164; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3166 = 8'h5e == io_state_in_12 ? 8'h9d : _GEN_3165; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3167 = 8'h5f == io_state_in_12 ? 8'h84 : _GEN_3166; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3168 = 8'h60 == io_state_in_12 ? 8'h90 : _GEN_3167; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3169 = 8'h61 == io_state_in_12 ? 8'hd8 : _GEN_3168; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3170 = 8'h62 == io_state_in_12 ? 8'hab : _GEN_3169; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3171 = 8'h63 == io_state_in_12 ? 8'h0 : _GEN_3170; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3172 = 8'h64 == io_state_in_12 ? 8'h8c : _GEN_3171; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3173 = 8'h65 == io_state_in_12 ? 8'hbc : _GEN_3172; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3174 = 8'h66 == io_state_in_12 ? 8'hd3 : _GEN_3173; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3175 = 8'h67 == io_state_in_12 ? 8'ha : _GEN_3174; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3176 = 8'h68 == io_state_in_12 ? 8'hf7 : _GEN_3175; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3177 = 8'h69 == io_state_in_12 ? 8'he4 : _GEN_3176; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3178 = 8'h6a == io_state_in_12 ? 8'h58 : _GEN_3177; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3179 = 8'h6b == io_state_in_12 ? 8'h5 : _GEN_3178; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3180 = 8'h6c == io_state_in_12 ? 8'hb8 : _GEN_3179; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3181 = 8'h6d == io_state_in_12 ? 8'hb3 : _GEN_3180; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3182 = 8'h6e == io_state_in_12 ? 8'h45 : _GEN_3181; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3183 = 8'h6f == io_state_in_12 ? 8'h6 : _GEN_3182; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3184 = 8'h70 == io_state_in_12 ? 8'hd0 : _GEN_3183; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3185 = 8'h71 == io_state_in_12 ? 8'h2c : _GEN_3184; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3186 = 8'h72 == io_state_in_12 ? 8'h1e : _GEN_3185; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3187 = 8'h73 == io_state_in_12 ? 8'h8f : _GEN_3186; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3188 = 8'h74 == io_state_in_12 ? 8'hca : _GEN_3187; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3189 = 8'h75 == io_state_in_12 ? 8'h3f : _GEN_3188; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3190 = 8'h76 == io_state_in_12 ? 8'hf : _GEN_3189; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3191 = 8'h77 == io_state_in_12 ? 8'h2 : _GEN_3190; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3192 = 8'h78 == io_state_in_12 ? 8'hc1 : _GEN_3191; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3193 = 8'h79 == io_state_in_12 ? 8'haf : _GEN_3192; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3194 = 8'h7a == io_state_in_12 ? 8'hbd : _GEN_3193; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3195 = 8'h7b == io_state_in_12 ? 8'h3 : _GEN_3194; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3196 = 8'h7c == io_state_in_12 ? 8'h1 : _GEN_3195; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3197 = 8'h7d == io_state_in_12 ? 8'h13 : _GEN_3196; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3198 = 8'h7e == io_state_in_12 ? 8'h8a : _GEN_3197; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3199 = 8'h7f == io_state_in_12 ? 8'h6b : _GEN_3198; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3200 = 8'h80 == io_state_in_12 ? 8'h3a : _GEN_3199; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3201 = 8'h81 == io_state_in_12 ? 8'h91 : _GEN_3200; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3202 = 8'h82 == io_state_in_12 ? 8'h11 : _GEN_3201; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3203 = 8'h83 == io_state_in_12 ? 8'h41 : _GEN_3202; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3204 = 8'h84 == io_state_in_12 ? 8'h4f : _GEN_3203; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3205 = 8'h85 == io_state_in_12 ? 8'h67 : _GEN_3204; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3206 = 8'h86 == io_state_in_12 ? 8'hdc : _GEN_3205; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3207 = 8'h87 == io_state_in_12 ? 8'hea : _GEN_3206; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3208 = 8'h88 == io_state_in_12 ? 8'h97 : _GEN_3207; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3209 = 8'h89 == io_state_in_12 ? 8'hf2 : _GEN_3208; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3210 = 8'h8a == io_state_in_12 ? 8'hcf : _GEN_3209; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3211 = 8'h8b == io_state_in_12 ? 8'hce : _GEN_3210; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3212 = 8'h8c == io_state_in_12 ? 8'hf0 : _GEN_3211; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3213 = 8'h8d == io_state_in_12 ? 8'hb4 : _GEN_3212; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3214 = 8'h8e == io_state_in_12 ? 8'he6 : _GEN_3213; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3215 = 8'h8f == io_state_in_12 ? 8'h73 : _GEN_3214; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3216 = 8'h90 == io_state_in_12 ? 8'h96 : _GEN_3215; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3217 = 8'h91 == io_state_in_12 ? 8'hac : _GEN_3216; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3218 = 8'h92 == io_state_in_12 ? 8'h74 : _GEN_3217; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3219 = 8'h93 == io_state_in_12 ? 8'h22 : _GEN_3218; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3220 = 8'h94 == io_state_in_12 ? 8'he7 : _GEN_3219; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3221 = 8'h95 == io_state_in_12 ? 8'had : _GEN_3220; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3222 = 8'h96 == io_state_in_12 ? 8'h35 : _GEN_3221; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3223 = 8'h97 == io_state_in_12 ? 8'h85 : _GEN_3222; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3224 = 8'h98 == io_state_in_12 ? 8'he2 : _GEN_3223; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3225 = 8'h99 == io_state_in_12 ? 8'hf9 : _GEN_3224; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3226 = 8'h9a == io_state_in_12 ? 8'h37 : _GEN_3225; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3227 = 8'h9b == io_state_in_12 ? 8'he8 : _GEN_3226; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3228 = 8'h9c == io_state_in_12 ? 8'h1c : _GEN_3227; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3229 = 8'h9d == io_state_in_12 ? 8'h75 : _GEN_3228; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3230 = 8'h9e == io_state_in_12 ? 8'hdf : _GEN_3229; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3231 = 8'h9f == io_state_in_12 ? 8'h6e : _GEN_3230; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3232 = 8'ha0 == io_state_in_12 ? 8'h47 : _GEN_3231; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3233 = 8'ha1 == io_state_in_12 ? 8'hf1 : _GEN_3232; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3234 = 8'ha2 == io_state_in_12 ? 8'h1a : _GEN_3233; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3235 = 8'ha3 == io_state_in_12 ? 8'h71 : _GEN_3234; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3236 = 8'ha4 == io_state_in_12 ? 8'h1d : _GEN_3235; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3237 = 8'ha5 == io_state_in_12 ? 8'h29 : _GEN_3236; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3238 = 8'ha6 == io_state_in_12 ? 8'hc5 : _GEN_3237; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3239 = 8'ha7 == io_state_in_12 ? 8'h89 : _GEN_3238; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3240 = 8'ha8 == io_state_in_12 ? 8'h6f : _GEN_3239; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3241 = 8'ha9 == io_state_in_12 ? 8'hb7 : _GEN_3240; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3242 = 8'haa == io_state_in_12 ? 8'h62 : _GEN_3241; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3243 = 8'hab == io_state_in_12 ? 8'he : _GEN_3242; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3244 = 8'hac == io_state_in_12 ? 8'haa : _GEN_3243; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3245 = 8'had == io_state_in_12 ? 8'h18 : _GEN_3244; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3246 = 8'hae == io_state_in_12 ? 8'hbe : _GEN_3245; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3247 = 8'haf == io_state_in_12 ? 8'h1b : _GEN_3246; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3248 = 8'hb0 == io_state_in_12 ? 8'hfc : _GEN_3247; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3249 = 8'hb1 == io_state_in_12 ? 8'h56 : _GEN_3248; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3250 = 8'hb2 == io_state_in_12 ? 8'h3e : _GEN_3249; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3251 = 8'hb3 == io_state_in_12 ? 8'h4b : _GEN_3250; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3252 = 8'hb4 == io_state_in_12 ? 8'hc6 : _GEN_3251; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3253 = 8'hb5 == io_state_in_12 ? 8'hd2 : _GEN_3252; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3254 = 8'hb6 == io_state_in_12 ? 8'h79 : _GEN_3253; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3255 = 8'hb7 == io_state_in_12 ? 8'h20 : _GEN_3254; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3256 = 8'hb8 == io_state_in_12 ? 8'h9a : _GEN_3255; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3257 = 8'hb9 == io_state_in_12 ? 8'hdb : _GEN_3256; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3258 = 8'hba == io_state_in_12 ? 8'hc0 : _GEN_3257; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3259 = 8'hbb == io_state_in_12 ? 8'hfe : _GEN_3258; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3260 = 8'hbc == io_state_in_12 ? 8'h78 : _GEN_3259; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3261 = 8'hbd == io_state_in_12 ? 8'hcd : _GEN_3260; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3262 = 8'hbe == io_state_in_12 ? 8'h5a : _GEN_3261; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3263 = 8'hbf == io_state_in_12 ? 8'hf4 : _GEN_3262; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3264 = 8'hc0 == io_state_in_12 ? 8'h1f : _GEN_3263; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3265 = 8'hc1 == io_state_in_12 ? 8'hdd : _GEN_3264; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3266 = 8'hc2 == io_state_in_12 ? 8'ha8 : _GEN_3265; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3267 = 8'hc3 == io_state_in_12 ? 8'h33 : _GEN_3266; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3268 = 8'hc4 == io_state_in_12 ? 8'h88 : _GEN_3267; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3269 = 8'hc5 == io_state_in_12 ? 8'h7 : _GEN_3268; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3270 = 8'hc6 == io_state_in_12 ? 8'hc7 : _GEN_3269; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3271 = 8'hc7 == io_state_in_12 ? 8'h31 : _GEN_3270; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3272 = 8'hc8 == io_state_in_12 ? 8'hb1 : _GEN_3271; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3273 = 8'hc9 == io_state_in_12 ? 8'h12 : _GEN_3272; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3274 = 8'hca == io_state_in_12 ? 8'h10 : _GEN_3273; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3275 = 8'hcb == io_state_in_12 ? 8'h59 : _GEN_3274; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3276 = 8'hcc == io_state_in_12 ? 8'h27 : _GEN_3275; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3277 = 8'hcd == io_state_in_12 ? 8'h80 : _GEN_3276; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3278 = 8'hce == io_state_in_12 ? 8'hec : _GEN_3277; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3279 = 8'hcf == io_state_in_12 ? 8'h5f : _GEN_3278; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3280 = 8'hd0 == io_state_in_12 ? 8'h60 : _GEN_3279; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3281 = 8'hd1 == io_state_in_12 ? 8'h51 : _GEN_3280; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3282 = 8'hd2 == io_state_in_12 ? 8'h7f : _GEN_3281; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3283 = 8'hd3 == io_state_in_12 ? 8'ha9 : _GEN_3282; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3284 = 8'hd4 == io_state_in_12 ? 8'h19 : _GEN_3283; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3285 = 8'hd5 == io_state_in_12 ? 8'hb5 : _GEN_3284; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3286 = 8'hd6 == io_state_in_12 ? 8'h4a : _GEN_3285; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3287 = 8'hd7 == io_state_in_12 ? 8'hd : _GEN_3286; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3288 = 8'hd8 == io_state_in_12 ? 8'h2d : _GEN_3287; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3289 = 8'hd9 == io_state_in_12 ? 8'he5 : _GEN_3288; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3290 = 8'hda == io_state_in_12 ? 8'h7a : _GEN_3289; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3291 = 8'hdb == io_state_in_12 ? 8'h9f : _GEN_3290; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3292 = 8'hdc == io_state_in_12 ? 8'h93 : _GEN_3291; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3293 = 8'hdd == io_state_in_12 ? 8'hc9 : _GEN_3292; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3294 = 8'hde == io_state_in_12 ? 8'h9c : _GEN_3293; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3295 = 8'hdf == io_state_in_12 ? 8'hef : _GEN_3294; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3296 = 8'he0 == io_state_in_12 ? 8'ha0 : _GEN_3295; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3297 = 8'he1 == io_state_in_12 ? 8'he0 : _GEN_3296; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3298 = 8'he2 == io_state_in_12 ? 8'h3b : _GEN_3297; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3299 = 8'he3 == io_state_in_12 ? 8'h4d : _GEN_3298; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3300 = 8'he4 == io_state_in_12 ? 8'hae : _GEN_3299; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3301 = 8'he5 == io_state_in_12 ? 8'h2a : _GEN_3300; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3302 = 8'he6 == io_state_in_12 ? 8'hf5 : _GEN_3301; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3303 = 8'he7 == io_state_in_12 ? 8'hb0 : _GEN_3302; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3304 = 8'he8 == io_state_in_12 ? 8'hc8 : _GEN_3303; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3305 = 8'he9 == io_state_in_12 ? 8'heb : _GEN_3304; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3306 = 8'hea == io_state_in_12 ? 8'hbb : _GEN_3305; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3307 = 8'heb == io_state_in_12 ? 8'h3c : _GEN_3306; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3308 = 8'hec == io_state_in_12 ? 8'h83 : _GEN_3307; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3309 = 8'hed == io_state_in_12 ? 8'h53 : _GEN_3308; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3310 = 8'hee == io_state_in_12 ? 8'h99 : _GEN_3309; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3311 = 8'hef == io_state_in_12 ? 8'h61 : _GEN_3310; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3312 = 8'hf0 == io_state_in_12 ? 8'h17 : _GEN_3311; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3313 = 8'hf1 == io_state_in_12 ? 8'h2b : _GEN_3312; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3314 = 8'hf2 == io_state_in_12 ? 8'h4 : _GEN_3313; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3315 = 8'hf3 == io_state_in_12 ? 8'h7e : _GEN_3314; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3316 = 8'hf4 == io_state_in_12 ? 8'hba : _GEN_3315; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3317 = 8'hf5 == io_state_in_12 ? 8'h77 : _GEN_3316; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3318 = 8'hf6 == io_state_in_12 ? 8'hd6 : _GEN_3317; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3319 = 8'hf7 == io_state_in_12 ? 8'h26 : _GEN_3318; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3320 = 8'hf8 == io_state_in_12 ? 8'he1 : _GEN_3319; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3321 = 8'hf9 == io_state_in_12 ? 8'h69 : _GEN_3320; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3322 = 8'hfa == io_state_in_12 ? 8'h14 : _GEN_3321; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3323 = 8'hfb == io_state_in_12 ? 8'h63 : _GEN_3322; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3324 = 8'hfc == io_state_in_12 ? 8'h55 : _GEN_3323; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3325 = 8'hfd == io_state_in_12 ? 8'h21 : _GEN_3324; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3326 = 8'hfe == io_state_in_12 ? 8'hc : _GEN_3325; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3329 = 8'h1 == io_state_in_13 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3330 = 8'h2 == io_state_in_13 ? 8'h6a : _GEN_3329; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3331 = 8'h3 == io_state_in_13 ? 8'hd5 : _GEN_3330; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3332 = 8'h4 == io_state_in_13 ? 8'h30 : _GEN_3331; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3333 = 8'h5 == io_state_in_13 ? 8'h36 : _GEN_3332; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3334 = 8'h6 == io_state_in_13 ? 8'ha5 : _GEN_3333; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3335 = 8'h7 == io_state_in_13 ? 8'h38 : _GEN_3334; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3336 = 8'h8 == io_state_in_13 ? 8'hbf : _GEN_3335; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3337 = 8'h9 == io_state_in_13 ? 8'h40 : _GEN_3336; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3338 = 8'ha == io_state_in_13 ? 8'ha3 : _GEN_3337; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3339 = 8'hb == io_state_in_13 ? 8'h9e : _GEN_3338; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3340 = 8'hc == io_state_in_13 ? 8'h81 : _GEN_3339; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3341 = 8'hd == io_state_in_13 ? 8'hf3 : _GEN_3340; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3342 = 8'he == io_state_in_13 ? 8'hd7 : _GEN_3341; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3343 = 8'hf == io_state_in_13 ? 8'hfb : _GEN_3342; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3344 = 8'h10 == io_state_in_13 ? 8'h7c : _GEN_3343; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3345 = 8'h11 == io_state_in_13 ? 8'he3 : _GEN_3344; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3346 = 8'h12 == io_state_in_13 ? 8'h39 : _GEN_3345; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3347 = 8'h13 == io_state_in_13 ? 8'h82 : _GEN_3346; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3348 = 8'h14 == io_state_in_13 ? 8'h9b : _GEN_3347; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3349 = 8'h15 == io_state_in_13 ? 8'h2f : _GEN_3348; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3350 = 8'h16 == io_state_in_13 ? 8'hff : _GEN_3349; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3351 = 8'h17 == io_state_in_13 ? 8'h87 : _GEN_3350; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3352 = 8'h18 == io_state_in_13 ? 8'h34 : _GEN_3351; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3353 = 8'h19 == io_state_in_13 ? 8'h8e : _GEN_3352; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3354 = 8'h1a == io_state_in_13 ? 8'h43 : _GEN_3353; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3355 = 8'h1b == io_state_in_13 ? 8'h44 : _GEN_3354; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3356 = 8'h1c == io_state_in_13 ? 8'hc4 : _GEN_3355; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3357 = 8'h1d == io_state_in_13 ? 8'hde : _GEN_3356; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3358 = 8'h1e == io_state_in_13 ? 8'he9 : _GEN_3357; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3359 = 8'h1f == io_state_in_13 ? 8'hcb : _GEN_3358; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3360 = 8'h20 == io_state_in_13 ? 8'h54 : _GEN_3359; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3361 = 8'h21 == io_state_in_13 ? 8'h7b : _GEN_3360; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3362 = 8'h22 == io_state_in_13 ? 8'h94 : _GEN_3361; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3363 = 8'h23 == io_state_in_13 ? 8'h32 : _GEN_3362; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3364 = 8'h24 == io_state_in_13 ? 8'ha6 : _GEN_3363; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3365 = 8'h25 == io_state_in_13 ? 8'hc2 : _GEN_3364; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3366 = 8'h26 == io_state_in_13 ? 8'h23 : _GEN_3365; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3367 = 8'h27 == io_state_in_13 ? 8'h3d : _GEN_3366; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3368 = 8'h28 == io_state_in_13 ? 8'hee : _GEN_3367; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3369 = 8'h29 == io_state_in_13 ? 8'h4c : _GEN_3368; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3370 = 8'h2a == io_state_in_13 ? 8'h95 : _GEN_3369; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3371 = 8'h2b == io_state_in_13 ? 8'hb : _GEN_3370; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3372 = 8'h2c == io_state_in_13 ? 8'h42 : _GEN_3371; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3373 = 8'h2d == io_state_in_13 ? 8'hfa : _GEN_3372; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3374 = 8'h2e == io_state_in_13 ? 8'hc3 : _GEN_3373; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3375 = 8'h2f == io_state_in_13 ? 8'h4e : _GEN_3374; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3376 = 8'h30 == io_state_in_13 ? 8'h8 : _GEN_3375; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3377 = 8'h31 == io_state_in_13 ? 8'h2e : _GEN_3376; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3378 = 8'h32 == io_state_in_13 ? 8'ha1 : _GEN_3377; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3379 = 8'h33 == io_state_in_13 ? 8'h66 : _GEN_3378; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3380 = 8'h34 == io_state_in_13 ? 8'h28 : _GEN_3379; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3381 = 8'h35 == io_state_in_13 ? 8'hd9 : _GEN_3380; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3382 = 8'h36 == io_state_in_13 ? 8'h24 : _GEN_3381; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3383 = 8'h37 == io_state_in_13 ? 8'hb2 : _GEN_3382; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3384 = 8'h38 == io_state_in_13 ? 8'h76 : _GEN_3383; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3385 = 8'h39 == io_state_in_13 ? 8'h5b : _GEN_3384; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3386 = 8'h3a == io_state_in_13 ? 8'ha2 : _GEN_3385; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3387 = 8'h3b == io_state_in_13 ? 8'h49 : _GEN_3386; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3388 = 8'h3c == io_state_in_13 ? 8'h6d : _GEN_3387; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3389 = 8'h3d == io_state_in_13 ? 8'h8b : _GEN_3388; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3390 = 8'h3e == io_state_in_13 ? 8'hd1 : _GEN_3389; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3391 = 8'h3f == io_state_in_13 ? 8'h25 : _GEN_3390; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3392 = 8'h40 == io_state_in_13 ? 8'h72 : _GEN_3391; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3393 = 8'h41 == io_state_in_13 ? 8'hf8 : _GEN_3392; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3394 = 8'h42 == io_state_in_13 ? 8'hf6 : _GEN_3393; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3395 = 8'h43 == io_state_in_13 ? 8'h64 : _GEN_3394; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3396 = 8'h44 == io_state_in_13 ? 8'h86 : _GEN_3395; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3397 = 8'h45 == io_state_in_13 ? 8'h68 : _GEN_3396; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3398 = 8'h46 == io_state_in_13 ? 8'h98 : _GEN_3397; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3399 = 8'h47 == io_state_in_13 ? 8'h16 : _GEN_3398; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3400 = 8'h48 == io_state_in_13 ? 8'hd4 : _GEN_3399; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3401 = 8'h49 == io_state_in_13 ? 8'ha4 : _GEN_3400; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3402 = 8'h4a == io_state_in_13 ? 8'h5c : _GEN_3401; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3403 = 8'h4b == io_state_in_13 ? 8'hcc : _GEN_3402; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3404 = 8'h4c == io_state_in_13 ? 8'h5d : _GEN_3403; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3405 = 8'h4d == io_state_in_13 ? 8'h65 : _GEN_3404; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3406 = 8'h4e == io_state_in_13 ? 8'hb6 : _GEN_3405; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3407 = 8'h4f == io_state_in_13 ? 8'h92 : _GEN_3406; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3408 = 8'h50 == io_state_in_13 ? 8'h6c : _GEN_3407; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3409 = 8'h51 == io_state_in_13 ? 8'h70 : _GEN_3408; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3410 = 8'h52 == io_state_in_13 ? 8'h48 : _GEN_3409; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3411 = 8'h53 == io_state_in_13 ? 8'h50 : _GEN_3410; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3412 = 8'h54 == io_state_in_13 ? 8'hfd : _GEN_3411; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3413 = 8'h55 == io_state_in_13 ? 8'hed : _GEN_3412; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3414 = 8'h56 == io_state_in_13 ? 8'hb9 : _GEN_3413; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3415 = 8'h57 == io_state_in_13 ? 8'hda : _GEN_3414; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3416 = 8'h58 == io_state_in_13 ? 8'h5e : _GEN_3415; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3417 = 8'h59 == io_state_in_13 ? 8'h15 : _GEN_3416; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3418 = 8'h5a == io_state_in_13 ? 8'h46 : _GEN_3417; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3419 = 8'h5b == io_state_in_13 ? 8'h57 : _GEN_3418; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3420 = 8'h5c == io_state_in_13 ? 8'ha7 : _GEN_3419; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3421 = 8'h5d == io_state_in_13 ? 8'h8d : _GEN_3420; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3422 = 8'h5e == io_state_in_13 ? 8'h9d : _GEN_3421; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3423 = 8'h5f == io_state_in_13 ? 8'h84 : _GEN_3422; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3424 = 8'h60 == io_state_in_13 ? 8'h90 : _GEN_3423; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3425 = 8'h61 == io_state_in_13 ? 8'hd8 : _GEN_3424; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3426 = 8'h62 == io_state_in_13 ? 8'hab : _GEN_3425; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3427 = 8'h63 == io_state_in_13 ? 8'h0 : _GEN_3426; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3428 = 8'h64 == io_state_in_13 ? 8'h8c : _GEN_3427; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3429 = 8'h65 == io_state_in_13 ? 8'hbc : _GEN_3428; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3430 = 8'h66 == io_state_in_13 ? 8'hd3 : _GEN_3429; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3431 = 8'h67 == io_state_in_13 ? 8'ha : _GEN_3430; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3432 = 8'h68 == io_state_in_13 ? 8'hf7 : _GEN_3431; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3433 = 8'h69 == io_state_in_13 ? 8'he4 : _GEN_3432; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3434 = 8'h6a == io_state_in_13 ? 8'h58 : _GEN_3433; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3435 = 8'h6b == io_state_in_13 ? 8'h5 : _GEN_3434; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3436 = 8'h6c == io_state_in_13 ? 8'hb8 : _GEN_3435; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3437 = 8'h6d == io_state_in_13 ? 8'hb3 : _GEN_3436; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3438 = 8'h6e == io_state_in_13 ? 8'h45 : _GEN_3437; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3439 = 8'h6f == io_state_in_13 ? 8'h6 : _GEN_3438; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3440 = 8'h70 == io_state_in_13 ? 8'hd0 : _GEN_3439; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3441 = 8'h71 == io_state_in_13 ? 8'h2c : _GEN_3440; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3442 = 8'h72 == io_state_in_13 ? 8'h1e : _GEN_3441; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3443 = 8'h73 == io_state_in_13 ? 8'h8f : _GEN_3442; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3444 = 8'h74 == io_state_in_13 ? 8'hca : _GEN_3443; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3445 = 8'h75 == io_state_in_13 ? 8'h3f : _GEN_3444; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3446 = 8'h76 == io_state_in_13 ? 8'hf : _GEN_3445; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3447 = 8'h77 == io_state_in_13 ? 8'h2 : _GEN_3446; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3448 = 8'h78 == io_state_in_13 ? 8'hc1 : _GEN_3447; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3449 = 8'h79 == io_state_in_13 ? 8'haf : _GEN_3448; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3450 = 8'h7a == io_state_in_13 ? 8'hbd : _GEN_3449; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3451 = 8'h7b == io_state_in_13 ? 8'h3 : _GEN_3450; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3452 = 8'h7c == io_state_in_13 ? 8'h1 : _GEN_3451; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3453 = 8'h7d == io_state_in_13 ? 8'h13 : _GEN_3452; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3454 = 8'h7e == io_state_in_13 ? 8'h8a : _GEN_3453; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3455 = 8'h7f == io_state_in_13 ? 8'h6b : _GEN_3454; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3456 = 8'h80 == io_state_in_13 ? 8'h3a : _GEN_3455; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3457 = 8'h81 == io_state_in_13 ? 8'h91 : _GEN_3456; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3458 = 8'h82 == io_state_in_13 ? 8'h11 : _GEN_3457; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3459 = 8'h83 == io_state_in_13 ? 8'h41 : _GEN_3458; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3460 = 8'h84 == io_state_in_13 ? 8'h4f : _GEN_3459; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3461 = 8'h85 == io_state_in_13 ? 8'h67 : _GEN_3460; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3462 = 8'h86 == io_state_in_13 ? 8'hdc : _GEN_3461; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3463 = 8'h87 == io_state_in_13 ? 8'hea : _GEN_3462; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3464 = 8'h88 == io_state_in_13 ? 8'h97 : _GEN_3463; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3465 = 8'h89 == io_state_in_13 ? 8'hf2 : _GEN_3464; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3466 = 8'h8a == io_state_in_13 ? 8'hcf : _GEN_3465; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3467 = 8'h8b == io_state_in_13 ? 8'hce : _GEN_3466; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3468 = 8'h8c == io_state_in_13 ? 8'hf0 : _GEN_3467; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3469 = 8'h8d == io_state_in_13 ? 8'hb4 : _GEN_3468; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3470 = 8'h8e == io_state_in_13 ? 8'he6 : _GEN_3469; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3471 = 8'h8f == io_state_in_13 ? 8'h73 : _GEN_3470; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3472 = 8'h90 == io_state_in_13 ? 8'h96 : _GEN_3471; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3473 = 8'h91 == io_state_in_13 ? 8'hac : _GEN_3472; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3474 = 8'h92 == io_state_in_13 ? 8'h74 : _GEN_3473; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3475 = 8'h93 == io_state_in_13 ? 8'h22 : _GEN_3474; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3476 = 8'h94 == io_state_in_13 ? 8'he7 : _GEN_3475; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3477 = 8'h95 == io_state_in_13 ? 8'had : _GEN_3476; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3478 = 8'h96 == io_state_in_13 ? 8'h35 : _GEN_3477; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3479 = 8'h97 == io_state_in_13 ? 8'h85 : _GEN_3478; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3480 = 8'h98 == io_state_in_13 ? 8'he2 : _GEN_3479; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3481 = 8'h99 == io_state_in_13 ? 8'hf9 : _GEN_3480; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3482 = 8'h9a == io_state_in_13 ? 8'h37 : _GEN_3481; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3483 = 8'h9b == io_state_in_13 ? 8'he8 : _GEN_3482; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3484 = 8'h9c == io_state_in_13 ? 8'h1c : _GEN_3483; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3485 = 8'h9d == io_state_in_13 ? 8'h75 : _GEN_3484; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3486 = 8'h9e == io_state_in_13 ? 8'hdf : _GEN_3485; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3487 = 8'h9f == io_state_in_13 ? 8'h6e : _GEN_3486; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3488 = 8'ha0 == io_state_in_13 ? 8'h47 : _GEN_3487; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3489 = 8'ha1 == io_state_in_13 ? 8'hf1 : _GEN_3488; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3490 = 8'ha2 == io_state_in_13 ? 8'h1a : _GEN_3489; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3491 = 8'ha3 == io_state_in_13 ? 8'h71 : _GEN_3490; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3492 = 8'ha4 == io_state_in_13 ? 8'h1d : _GEN_3491; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3493 = 8'ha5 == io_state_in_13 ? 8'h29 : _GEN_3492; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3494 = 8'ha6 == io_state_in_13 ? 8'hc5 : _GEN_3493; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3495 = 8'ha7 == io_state_in_13 ? 8'h89 : _GEN_3494; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3496 = 8'ha8 == io_state_in_13 ? 8'h6f : _GEN_3495; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3497 = 8'ha9 == io_state_in_13 ? 8'hb7 : _GEN_3496; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3498 = 8'haa == io_state_in_13 ? 8'h62 : _GEN_3497; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3499 = 8'hab == io_state_in_13 ? 8'he : _GEN_3498; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3500 = 8'hac == io_state_in_13 ? 8'haa : _GEN_3499; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3501 = 8'had == io_state_in_13 ? 8'h18 : _GEN_3500; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3502 = 8'hae == io_state_in_13 ? 8'hbe : _GEN_3501; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3503 = 8'haf == io_state_in_13 ? 8'h1b : _GEN_3502; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3504 = 8'hb0 == io_state_in_13 ? 8'hfc : _GEN_3503; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3505 = 8'hb1 == io_state_in_13 ? 8'h56 : _GEN_3504; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3506 = 8'hb2 == io_state_in_13 ? 8'h3e : _GEN_3505; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3507 = 8'hb3 == io_state_in_13 ? 8'h4b : _GEN_3506; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3508 = 8'hb4 == io_state_in_13 ? 8'hc6 : _GEN_3507; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3509 = 8'hb5 == io_state_in_13 ? 8'hd2 : _GEN_3508; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3510 = 8'hb6 == io_state_in_13 ? 8'h79 : _GEN_3509; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3511 = 8'hb7 == io_state_in_13 ? 8'h20 : _GEN_3510; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3512 = 8'hb8 == io_state_in_13 ? 8'h9a : _GEN_3511; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3513 = 8'hb9 == io_state_in_13 ? 8'hdb : _GEN_3512; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3514 = 8'hba == io_state_in_13 ? 8'hc0 : _GEN_3513; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3515 = 8'hbb == io_state_in_13 ? 8'hfe : _GEN_3514; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3516 = 8'hbc == io_state_in_13 ? 8'h78 : _GEN_3515; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3517 = 8'hbd == io_state_in_13 ? 8'hcd : _GEN_3516; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3518 = 8'hbe == io_state_in_13 ? 8'h5a : _GEN_3517; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3519 = 8'hbf == io_state_in_13 ? 8'hf4 : _GEN_3518; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3520 = 8'hc0 == io_state_in_13 ? 8'h1f : _GEN_3519; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3521 = 8'hc1 == io_state_in_13 ? 8'hdd : _GEN_3520; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3522 = 8'hc2 == io_state_in_13 ? 8'ha8 : _GEN_3521; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3523 = 8'hc3 == io_state_in_13 ? 8'h33 : _GEN_3522; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3524 = 8'hc4 == io_state_in_13 ? 8'h88 : _GEN_3523; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3525 = 8'hc5 == io_state_in_13 ? 8'h7 : _GEN_3524; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3526 = 8'hc6 == io_state_in_13 ? 8'hc7 : _GEN_3525; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3527 = 8'hc7 == io_state_in_13 ? 8'h31 : _GEN_3526; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3528 = 8'hc8 == io_state_in_13 ? 8'hb1 : _GEN_3527; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3529 = 8'hc9 == io_state_in_13 ? 8'h12 : _GEN_3528; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3530 = 8'hca == io_state_in_13 ? 8'h10 : _GEN_3529; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3531 = 8'hcb == io_state_in_13 ? 8'h59 : _GEN_3530; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3532 = 8'hcc == io_state_in_13 ? 8'h27 : _GEN_3531; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3533 = 8'hcd == io_state_in_13 ? 8'h80 : _GEN_3532; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3534 = 8'hce == io_state_in_13 ? 8'hec : _GEN_3533; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3535 = 8'hcf == io_state_in_13 ? 8'h5f : _GEN_3534; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3536 = 8'hd0 == io_state_in_13 ? 8'h60 : _GEN_3535; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3537 = 8'hd1 == io_state_in_13 ? 8'h51 : _GEN_3536; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3538 = 8'hd2 == io_state_in_13 ? 8'h7f : _GEN_3537; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3539 = 8'hd3 == io_state_in_13 ? 8'ha9 : _GEN_3538; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3540 = 8'hd4 == io_state_in_13 ? 8'h19 : _GEN_3539; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3541 = 8'hd5 == io_state_in_13 ? 8'hb5 : _GEN_3540; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3542 = 8'hd6 == io_state_in_13 ? 8'h4a : _GEN_3541; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3543 = 8'hd7 == io_state_in_13 ? 8'hd : _GEN_3542; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3544 = 8'hd8 == io_state_in_13 ? 8'h2d : _GEN_3543; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3545 = 8'hd9 == io_state_in_13 ? 8'he5 : _GEN_3544; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3546 = 8'hda == io_state_in_13 ? 8'h7a : _GEN_3545; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3547 = 8'hdb == io_state_in_13 ? 8'h9f : _GEN_3546; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3548 = 8'hdc == io_state_in_13 ? 8'h93 : _GEN_3547; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3549 = 8'hdd == io_state_in_13 ? 8'hc9 : _GEN_3548; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3550 = 8'hde == io_state_in_13 ? 8'h9c : _GEN_3549; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3551 = 8'hdf == io_state_in_13 ? 8'hef : _GEN_3550; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3552 = 8'he0 == io_state_in_13 ? 8'ha0 : _GEN_3551; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3553 = 8'he1 == io_state_in_13 ? 8'he0 : _GEN_3552; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3554 = 8'he2 == io_state_in_13 ? 8'h3b : _GEN_3553; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3555 = 8'he3 == io_state_in_13 ? 8'h4d : _GEN_3554; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3556 = 8'he4 == io_state_in_13 ? 8'hae : _GEN_3555; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3557 = 8'he5 == io_state_in_13 ? 8'h2a : _GEN_3556; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3558 = 8'he6 == io_state_in_13 ? 8'hf5 : _GEN_3557; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3559 = 8'he7 == io_state_in_13 ? 8'hb0 : _GEN_3558; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3560 = 8'he8 == io_state_in_13 ? 8'hc8 : _GEN_3559; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3561 = 8'he9 == io_state_in_13 ? 8'heb : _GEN_3560; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3562 = 8'hea == io_state_in_13 ? 8'hbb : _GEN_3561; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3563 = 8'heb == io_state_in_13 ? 8'h3c : _GEN_3562; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3564 = 8'hec == io_state_in_13 ? 8'h83 : _GEN_3563; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3565 = 8'hed == io_state_in_13 ? 8'h53 : _GEN_3564; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3566 = 8'hee == io_state_in_13 ? 8'h99 : _GEN_3565; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3567 = 8'hef == io_state_in_13 ? 8'h61 : _GEN_3566; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3568 = 8'hf0 == io_state_in_13 ? 8'h17 : _GEN_3567; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3569 = 8'hf1 == io_state_in_13 ? 8'h2b : _GEN_3568; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3570 = 8'hf2 == io_state_in_13 ? 8'h4 : _GEN_3569; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3571 = 8'hf3 == io_state_in_13 ? 8'h7e : _GEN_3570; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3572 = 8'hf4 == io_state_in_13 ? 8'hba : _GEN_3571; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3573 = 8'hf5 == io_state_in_13 ? 8'h77 : _GEN_3572; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3574 = 8'hf6 == io_state_in_13 ? 8'hd6 : _GEN_3573; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3575 = 8'hf7 == io_state_in_13 ? 8'h26 : _GEN_3574; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3576 = 8'hf8 == io_state_in_13 ? 8'he1 : _GEN_3575; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3577 = 8'hf9 == io_state_in_13 ? 8'h69 : _GEN_3576; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3578 = 8'hfa == io_state_in_13 ? 8'h14 : _GEN_3577; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3579 = 8'hfb == io_state_in_13 ? 8'h63 : _GEN_3578; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3580 = 8'hfc == io_state_in_13 ? 8'h55 : _GEN_3579; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3581 = 8'hfd == io_state_in_13 ? 8'h21 : _GEN_3580; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3582 = 8'hfe == io_state_in_13 ? 8'hc : _GEN_3581; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3585 = 8'h1 == io_state_in_14 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3586 = 8'h2 == io_state_in_14 ? 8'h6a : _GEN_3585; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3587 = 8'h3 == io_state_in_14 ? 8'hd5 : _GEN_3586; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3588 = 8'h4 == io_state_in_14 ? 8'h30 : _GEN_3587; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3589 = 8'h5 == io_state_in_14 ? 8'h36 : _GEN_3588; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3590 = 8'h6 == io_state_in_14 ? 8'ha5 : _GEN_3589; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3591 = 8'h7 == io_state_in_14 ? 8'h38 : _GEN_3590; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3592 = 8'h8 == io_state_in_14 ? 8'hbf : _GEN_3591; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3593 = 8'h9 == io_state_in_14 ? 8'h40 : _GEN_3592; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3594 = 8'ha == io_state_in_14 ? 8'ha3 : _GEN_3593; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3595 = 8'hb == io_state_in_14 ? 8'h9e : _GEN_3594; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3596 = 8'hc == io_state_in_14 ? 8'h81 : _GEN_3595; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3597 = 8'hd == io_state_in_14 ? 8'hf3 : _GEN_3596; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3598 = 8'he == io_state_in_14 ? 8'hd7 : _GEN_3597; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3599 = 8'hf == io_state_in_14 ? 8'hfb : _GEN_3598; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3600 = 8'h10 == io_state_in_14 ? 8'h7c : _GEN_3599; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3601 = 8'h11 == io_state_in_14 ? 8'he3 : _GEN_3600; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3602 = 8'h12 == io_state_in_14 ? 8'h39 : _GEN_3601; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3603 = 8'h13 == io_state_in_14 ? 8'h82 : _GEN_3602; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3604 = 8'h14 == io_state_in_14 ? 8'h9b : _GEN_3603; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3605 = 8'h15 == io_state_in_14 ? 8'h2f : _GEN_3604; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3606 = 8'h16 == io_state_in_14 ? 8'hff : _GEN_3605; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3607 = 8'h17 == io_state_in_14 ? 8'h87 : _GEN_3606; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3608 = 8'h18 == io_state_in_14 ? 8'h34 : _GEN_3607; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3609 = 8'h19 == io_state_in_14 ? 8'h8e : _GEN_3608; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3610 = 8'h1a == io_state_in_14 ? 8'h43 : _GEN_3609; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3611 = 8'h1b == io_state_in_14 ? 8'h44 : _GEN_3610; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3612 = 8'h1c == io_state_in_14 ? 8'hc4 : _GEN_3611; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3613 = 8'h1d == io_state_in_14 ? 8'hde : _GEN_3612; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3614 = 8'h1e == io_state_in_14 ? 8'he9 : _GEN_3613; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3615 = 8'h1f == io_state_in_14 ? 8'hcb : _GEN_3614; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3616 = 8'h20 == io_state_in_14 ? 8'h54 : _GEN_3615; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3617 = 8'h21 == io_state_in_14 ? 8'h7b : _GEN_3616; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3618 = 8'h22 == io_state_in_14 ? 8'h94 : _GEN_3617; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3619 = 8'h23 == io_state_in_14 ? 8'h32 : _GEN_3618; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3620 = 8'h24 == io_state_in_14 ? 8'ha6 : _GEN_3619; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3621 = 8'h25 == io_state_in_14 ? 8'hc2 : _GEN_3620; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3622 = 8'h26 == io_state_in_14 ? 8'h23 : _GEN_3621; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3623 = 8'h27 == io_state_in_14 ? 8'h3d : _GEN_3622; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3624 = 8'h28 == io_state_in_14 ? 8'hee : _GEN_3623; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3625 = 8'h29 == io_state_in_14 ? 8'h4c : _GEN_3624; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3626 = 8'h2a == io_state_in_14 ? 8'h95 : _GEN_3625; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3627 = 8'h2b == io_state_in_14 ? 8'hb : _GEN_3626; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3628 = 8'h2c == io_state_in_14 ? 8'h42 : _GEN_3627; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3629 = 8'h2d == io_state_in_14 ? 8'hfa : _GEN_3628; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3630 = 8'h2e == io_state_in_14 ? 8'hc3 : _GEN_3629; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3631 = 8'h2f == io_state_in_14 ? 8'h4e : _GEN_3630; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3632 = 8'h30 == io_state_in_14 ? 8'h8 : _GEN_3631; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3633 = 8'h31 == io_state_in_14 ? 8'h2e : _GEN_3632; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3634 = 8'h32 == io_state_in_14 ? 8'ha1 : _GEN_3633; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3635 = 8'h33 == io_state_in_14 ? 8'h66 : _GEN_3634; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3636 = 8'h34 == io_state_in_14 ? 8'h28 : _GEN_3635; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3637 = 8'h35 == io_state_in_14 ? 8'hd9 : _GEN_3636; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3638 = 8'h36 == io_state_in_14 ? 8'h24 : _GEN_3637; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3639 = 8'h37 == io_state_in_14 ? 8'hb2 : _GEN_3638; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3640 = 8'h38 == io_state_in_14 ? 8'h76 : _GEN_3639; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3641 = 8'h39 == io_state_in_14 ? 8'h5b : _GEN_3640; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3642 = 8'h3a == io_state_in_14 ? 8'ha2 : _GEN_3641; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3643 = 8'h3b == io_state_in_14 ? 8'h49 : _GEN_3642; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3644 = 8'h3c == io_state_in_14 ? 8'h6d : _GEN_3643; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3645 = 8'h3d == io_state_in_14 ? 8'h8b : _GEN_3644; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3646 = 8'h3e == io_state_in_14 ? 8'hd1 : _GEN_3645; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3647 = 8'h3f == io_state_in_14 ? 8'h25 : _GEN_3646; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3648 = 8'h40 == io_state_in_14 ? 8'h72 : _GEN_3647; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3649 = 8'h41 == io_state_in_14 ? 8'hf8 : _GEN_3648; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3650 = 8'h42 == io_state_in_14 ? 8'hf6 : _GEN_3649; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3651 = 8'h43 == io_state_in_14 ? 8'h64 : _GEN_3650; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3652 = 8'h44 == io_state_in_14 ? 8'h86 : _GEN_3651; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3653 = 8'h45 == io_state_in_14 ? 8'h68 : _GEN_3652; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3654 = 8'h46 == io_state_in_14 ? 8'h98 : _GEN_3653; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3655 = 8'h47 == io_state_in_14 ? 8'h16 : _GEN_3654; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3656 = 8'h48 == io_state_in_14 ? 8'hd4 : _GEN_3655; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3657 = 8'h49 == io_state_in_14 ? 8'ha4 : _GEN_3656; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3658 = 8'h4a == io_state_in_14 ? 8'h5c : _GEN_3657; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3659 = 8'h4b == io_state_in_14 ? 8'hcc : _GEN_3658; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3660 = 8'h4c == io_state_in_14 ? 8'h5d : _GEN_3659; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3661 = 8'h4d == io_state_in_14 ? 8'h65 : _GEN_3660; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3662 = 8'h4e == io_state_in_14 ? 8'hb6 : _GEN_3661; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3663 = 8'h4f == io_state_in_14 ? 8'h92 : _GEN_3662; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3664 = 8'h50 == io_state_in_14 ? 8'h6c : _GEN_3663; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3665 = 8'h51 == io_state_in_14 ? 8'h70 : _GEN_3664; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3666 = 8'h52 == io_state_in_14 ? 8'h48 : _GEN_3665; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3667 = 8'h53 == io_state_in_14 ? 8'h50 : _GEN_3666; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3668 = 8'h54 == io_state_in_14 ? 8'hfd : _GEN_3667; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3669 = 8'h55 == io_state_in_14 ? 8'hed : _GEN_3668; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3670 = 8'h56 == io_state_in_14 ? 8'hb9 : _GEN_3669; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3671 = 8'h57 == io_state_in_14 ? 8'hda : _GEN_3670; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3672 = 8'h58 == io_state_in_14 ? 8'h5e : _GEN_3671; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3673 = 8'h59 == io_state_in_14 ? 8'h15 : _GEN_3672; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3674 = 8'h5a == io_state_in_14 ? 8'h46 : _GEN_3673; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3675 = 8'h5b == io_state_in_14 ? 8'h57 : _GEN_3674; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3676 = 8'h5c == io_state_in_14 ? 8'ha7 : _GEN_3675; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3677 = 8'h5d == io_state_in_14 ? 8'h8d : _GEN_3676; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3678 = 8'h5e == io_state_in_14 ? 8'h9d : _GEN_3677; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3679 = 8'h5f == io_state_in_14 ? 8'h84 : _GEN_3678; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3680 = 8'h60 == io_state_in_14 ? 8'h90 : _GEN_3679; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3681 = 8'h61 == io_state_in_14 ? 8'hd8 : _GEN_3680; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3682 = 8'h62 == io_state_in_14 ? 8'hab : _GEN_3681; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3683 = 8'h63 == io_state_in_14 ? 8'h0 : _GEN_3682; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3684 = 8'h64 == io_state_in_14 ? 8'h8c : _GEN_3683; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3685 = 8'h65 == io_state_in_14 ? 8'hbc : _GEN_3684; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3686 = 8'h66 == io_state_in_14 ? 8'hd3 : _GEN_3685; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3687 = 8'h67 == io_state_in_14 ? 8'ha : _GEN_3686; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3688 = 8'h68 == io_state_in_14 ? 8'hf7 : _GEN_3687; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3689 = 8'h69 == io_state_in_14 ? 8'he4 : _GEN_3688; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3690 = 8'h6a == io_state_in_14 ? 8'h58 : _GEN_3689; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3691 = 8'h6b == io_state_in_14 ? 8'h5 : _GEN_3690; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3692 = 8'h6c == io_state_in_14 ? 8'hb8 : _GEN_3691; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3693 = 8'h6d == io_state_in_14 ? 8'hb3 : _GEN_3692; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3694 = 8'h6e == io_state_in_14 ? 8'h45 : _GEN_3693; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3695 = 8'h6f == io_state_in_14 ? 8'h6 : _GEN_3694; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3696 = 8'h70 == io_state_in_14 ? 8'hd0 : _GEN_3695; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3697 = 8'h71 == io_state_in_14 ? 8'h2c : _GEN_3696; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3698 = 8'h72 == io_state_in_14 ? 8'h1e : _GEN_3697; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3699 = 8'h73 == io_state_in_14 ? 8'h8f : _GEN_3698; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3700 = 8'h74 == io_state_in_14 ? 8'hca : _GEN_3699; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3701 = 8'h75 == io_state_in_14 ? 8'h3f : _GEN_3700; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3702 = 8'h76 == io_state_in_14 ? 8'hf : _GEN_3701; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3703 = 8'h77 == io_state_in_14 ? 8'h2 : _GEN_3702; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3704 = 8'h78 == io_state_in_14 ? 8'hc1 : _GEN_3703; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3705 = 8'h79 == io_state_in_14 ? 8'haf : _GEN_3704; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3706 = 8'h7a == io_state_in_14 ? 8'hbd : _GEN_3705; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3707 = 8'h7b == io_state_in_14 ? 8'h3 : _GEN_3706; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3708 = 8'h7c == io_state_in_14 ? 8'h1 : _GEN_3707; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3709 = 8'h7d == io_state_in_14 ? 8'h13 : _GEN_3708; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3710 = 8'h7e == io_state_in_14 ? 8'h8a : _GEN_3709; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3711 = 8'h7f == io_state_in_14 ? 8'h6b : _GEN_3710; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3712 = 8'h80 == io_state_in_14 ? 8'h3a : _GEN_3711; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3713 = 8'h81 == io_state_in_14 ? 8'h91 : _GEN_3712; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3714 = 8'h82 == io_state_in_14 ? 8'h11 : _GEN_3713; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3715 = 8'h83 == io_state_in_14 ? 8'h41 : _GEN_3714; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3716 = 8'h84 == io_state_in_14 ? 8'h4f : _GEN_3715; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3717 = 8'h85 == io_state_in_14 ? 8'h67 : _GEN_3716; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3718 = 8'h86 == io_state_in_14 ? 8'hdc : _GEN_3717; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3719 = 8'h87 == io_state_in_14 ? 8'hea : _GEN_3718; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3720 = 8'h88 == io_state_in_14 ? 8'h97 : _GEN_3719; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3721 = 8'h89 == io_state_in_14 ? 8'hf2 : _GEN_3720; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3722 = 8'h8a == io_state_in_14 ? 8'hcf : _GEN_3721; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3723 = 8'h8b == io_state_in_14 ? 8'hce : _GEN_3722; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3724 = 8'h8c == io_state_in_14 ? 8'hf0 : _GEN_3723; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3725 = 8'h8d == io_state_in_14 ? 8'hb4 : _GEN_3724; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3726 = 8'h8e == io_state_in_14 ? 8'he6 : _GEN_3725; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3727 = 8'h8f == io_state_in_14 ? 8'h73 : _GEN_3726; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3728 = 8'h90 == io_state_in_14 ? 8'h96 : _GEN_3727; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3729 = 8'h91 == io_state_in_14 ? 8'hac : _GEN_3728; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3730 = 8'h92 == io_state_in_14 ? 8'h74 : _GEN_3729; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3731 = 8'h93 == io_state_in_14 ? 8'h22 : _GEN_3730; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3732 = 8'h94 == io_state_in_14 ? 8'he7 : _GEN_3731; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3733 = 8'h95 == io_state_in_14 ? 8'had : _GEN_3732; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3734 = 8'h96 == io_state_in_14 ? 8'h35 : _GEN_3733; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3735 = 8'h97 == io_state_in_14 ? 8'h85 : _GEN_3734; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3736 = 8'h98 == io_state_in_14 ? 8'he2 : _GEN_3735; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3737 = 8'h99 == io_state_in_14 ? 8'hf9 : _GEN_3736; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3738 = 8'h9a == io_state_in_14 ? 8'h37 : _GEN_3737; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3739 = 8'h9b == io_state_in_14 ? 8'he8 : _GEN_3738; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3740 = 8'h9c == io_state_in_14 ? 8'h1c : _GEN_3739; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3741 = 8'h9d == io_state_in_14 ? 8'h75 : _GEN_3740; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3742 = 8'h9e == io_state_in_14 ? 8'hdf : _GEN_3741; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3743 = 8'h9f == io_state_in_14 ? 8'h6e : _GEN_3742; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3744 = 8'ha0 == io_state_in_14 ? 8'h47 : _GEN_3743; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3745 = 8'ha1 == io_state_in_14 ? 8'hf1 : _GEN_3744; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3746 = 8'ha2 == io_state_in_14 ? 8'h1a : _GEN_3745; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3747 = 8'ha3 == io_state_in_14 ? 8'h71 : _GEN_3746; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3748 = 8'ha4 == io_state_in_14 ? 8'h1d : _GEN_3747; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3749 = 8'ha5 == io_state_in_14 ? 8'h29 : _GEN_3748; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3750 = 8'ha6 == io_state_in_14 ? 8'hc5 : _GEN_3749; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3751 = 8'ha7 == io_state_in_14 ? 8'h89 : _GEN_3750; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3752 = 8'ha8 == io_state_in_14 ? 8'h6f : _GEN_3751; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3753 = 8'ha9 == io_state_in_14 ? 8'hb7 : _GEN_3752; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3754 = 8'haa == io_state_in_14 ? 8'h62 : _GEN_3753; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3755 = 8'hab == io_state_in_14 ? 8'he : _GEN_3754; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3756 = 8'hac == io_state_in_14 ? 8'haa : _GEN_3755; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3757 = 8'had == io_state_in_14 ? 8'h18 : _GEN_3756; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3758 = 8'hae == io_state_in_14 ? 8'hbe : _GEN_3757; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3759 = 8'haf == io_state_in_14 ? 8'h1b : _GEN_3758; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3760 = 8'hb0 == io_state_in_14 ? 8'hfc : _GEN_3759; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3761 = 8'hb1 == io_state_in_14 ? 8'h56 : _GEN_3760; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3762 = 8'hb2 == io_state_in_14 ? 8'h3e : _GEN_3761; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3763 = 8'hb3 == io_state_in_14 ? 8'h4b : _GEN_3762; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3764 = 8'hb4 == io_state_in_14 ? 8'hc6 : _GEN_3763; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3765 = 8'hb5 == io_state_in_14 ? 8'hd2 : _GEN_3764; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3766 = 8'hb6 == io_state_in_14 ? 8'h79 : _GEN_3765; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3767 = 8'hb7 == io_state_in_14 ? 8'h20 : _GEN_3766; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3768 = 8'hb8 == io_state_in_14 ? 8'h9a : _GEN_3767; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3769 = 8'hb9 == io_state_in_14 ? 8'hdb : _GEN_3768; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3770 = 8'hba == io_state_in_14 ? 8'hc0 : _GEN_3769; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3771 = 8'hbb == io_state_in_14 ? 8'hfe : _GEN_3770; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3772 = 8'hbc == io_state_in_14 ? 8'h78 : _GEN_3771; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3773 = 8'hbd == io_state_in_14 ? 8'hcd : _GEN_3772; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3774 = 8'hbe == io_state_in_14 ? 8'h5a : _GEN_3773; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3775 = 8'hbf == io_state_in_14 ? 8'hf4 : _GEN_3774; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3776 = 8'hc0 == io_state_in_14 ? 8'h1f : _GEN_3775; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3777 = 8'hc1 == io_state_in_14 ? 8'hdd : _GEN_3776; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3778 = 8'hc2 == io_state_in_14 ? 8'ha8 : _GEN_3777; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3779 = 8'hc3 == io_state_in_14 ? 8'h33 : _GEN_3778; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3780 = 8'hc4 == io_state_in_14 ? 8'h88 : _GEN_3779; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3781 = 8'hc5 == io_state_in_14 ? 8'h7 : _GEN_3780; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3782 = 8'hc6 == io_state_in_14 ? 8'hc7 : _GEN_3781; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3783 = 8'hc7 == io_state_in_14 ? 8'h31 : _GEN_3782; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3784 = 8'hc8 == io_state_in_14 ? 8'hb1 : _GEN_3783; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3785 = 8'hc9 == io_state_in_14 ? 8'h12 : _GEN_3784; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3786 = 8'hca == io_state_in_14 ? 8'h10 : _GEN_3785; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3787 = 8'hcb == io_state_in_14 ? 8'h59 : _GEN_3786; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3788 = 8'hcc == io_state_in_14 ? 8'h27 : _GEN_3787; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3789 = 8'hcd == io_state_in_14 ? 8'h80 : _GEN_3788; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3790 = 8'hce == io_state_in_14 ? 8'hec : _GEN_3789; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3791 = 8'hcf == io_state_in_14 ? 8'h5f : _GEN_3790; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3792 = 8'hd0 == io_state_in_14 ? 8'h60 : _GEN_3791; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3793 = 8'hd1 == io_state_in_14 ? 8'h51 : _GEN_3792; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3794 = 8'hd2 == io_state_in_14 ? 8'h7f : _GEN_3793; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3795 = 8'hd3 == io_state_in_14 ? 8'ha9 : _GEN_3794; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3796 = 8'hd4 == io_state_in_14 ? 8'h19 : _GEN_3795; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3797 = 8'hd5 == io_state_in_14 ? 8'hb5 : _GEN_3796; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3798 = 8'hd6 == io_state_in_14 ? 8'h4a : _GEN_3797; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3799 = 8'hd7 == io_state_in_14 ? 8'hd : _GEN_3798; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3800 = 8'hd8 == io_state_in_14 ? 8'h2d : _GEN_3799; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3801 = 8'hd9 == io_state_in_14 ? 8'he5 : _GEN_3800; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3802 = 8'hda == io_state_in_14 ? 8'h7a : _GEN_3801; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3803 = 8'hdb == io_state_in_14 ? 8'h9f : _GEN_3802; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3804 = 8'hdc == io_state_in_14 ? 8'h93 : _GEN_3803; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3805 = 8'hdd == io_state_in_14 ? 8'hc9 : _GEN_3804; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3806 = 8'hde == io_state_in_14 ? 8'h9c : _GEN_3805; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3807 = 8'hdf == io_state_in_14 ? 8'hef : _GEN_3806; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3808 = 8'he0 == io_state_in_14 ? 8'ha0 : _GEN_3807; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3809 = 8'he1 == io_state_in_14 ? 8'he0 : _GEN_3808; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3810 = 8'he2 == io_state_in_14 ? 8'h3b : _GEN_3809; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3811 = 8'he3 == io_state_in_14 ? 8'h4d : _GEN_3810; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3812 = 8'he4 == io_state_in_14 ? 8'hae : _GEN_3811; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3813 = 8'he5 == io_state_in_14 ? 8'h2a : _GEN_3812; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3814 = 8'he6 == io_state_in_14 ? 8'hf5 : _GEN_3813; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3815 = 8'he7 == io_state_in_14 ? 8'hb0 : _GEN_3814; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3816 = 8'he8 == io_state_in_14 ? 8'hc8 : _GEN_3815; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3817 = 8'he9 == io_state_in_14 ? 8'heb : _GEN_3816; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3818 = 8'hea == io_state_in_14 ? 8'hbb : _GEN_3817; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3819 = 8'heb == io_state_in_14 ? 8'h3c : _GEN_3818; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3820 = 8'hec == io_state_in_14 ? 8'h83 : _GEN_3819; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3821 = 8'hed == io_state_in_14 ? 8'h53 : _GEN_3820; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3822 = 8'hee == io_state_in_14 ? 8'h99 : _GEN_3821; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3823 = 8'hef == io_state_in_14 ? 8'h61 : _GEN_3822; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3824 = 8'hf0 == io_state_in_14 ? 8'h17 : _GEN_3823; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3825 = 8'hf1 == io_state_in_14 ? 8'h2b : _GEN_3824; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3826 = 8'hf2 == io_state_in_14 ? 8'h4 : _GEN_3825; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3827 = 8'hf3 == io_state_in_14 ? 8'h7e : _GEN_3826; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3828 = 8'hf4 == io_state_in_14 ? 8'hba : _GEN_3827; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3829 = 8'hf5 == io_state_in_14 ? 8'h77 : _GEN_3828; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3830 = 8'hf6 == io_state_in_14 ? 8'hd6 : _GEN_3829; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3831 = 8'hf7 == io_state_in_14 ? 8'h26 : _GEN_3830; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3832 = 8'hf8 == io_state_in_14 ? 8'he1 : _GEN_3831; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3833 = 8'hf9 == io_state_in_14 ? 8'h69 : _GEN_3832; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3834 = 8'hfa == io_state_in_14 ? 8'h14 : _GEN_3833; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3835 = 8'hfb == io_state_in_14 ? 8'h63 : _GEN_3834; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3836 = 8'hfc == io_state_in_14 ? 8'h55 : _GEN_3835; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3837 = 8'hfd == io_state_in_14 ? 8'h21 : _GEN_3836; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3838 = 8'hfe == io_state_in_14 ? 8'hc : _GEN_3837; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3841 = 8'h1 == io_state_in_15 ? 8'h9 : 8'h52; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3842 = 8'h2 == io_state_in_15 ? 8'h6a : _GEN_3841; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3843 = 8'h3 == io_state_in_15 ? 8'hd5 : _GEN_3842; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3844 = 8'h4 == io_state_in_15 ? 8'h30 : _GEN_3843; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3845 = 8'h5 == io_state_in_15 ? 8'h36 : _GEN_3844; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3846 = 8'h6 == io_state_in_15 ? 8'ha5 : _GEN_3845; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3847 = 8'h7 == io_state_in_15 ? 8'h38 : _GEN_3846; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3848 = 8'h8 == io_state_in_15 ? 8'hbf : _GEN_3847; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3849 = 8'h9 == io_state_in_15 ? 8'h40 : _GEN_3848; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3850 = 8'ha == io_state_in_15 ? 8'ha3 : _GEN_3849; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3851 = 8'hb == io_state_in_15 ? 8'h9e : _GEN_3850; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3852 = 8'hc == io_state_in_15 ? 8'h81 : _GEN_3851; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3853 = 8'hd == io_state_in_15 ? 8'hf3 : _GEN_3852; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3854 = 8'he == io_state_in_15 ? 8'hd7 : _GEN_3853; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3855 = 8'hf == io_state_in_15 ? 8'hfb : _GEN_3854; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3856 = 8'h10 == io_state_in_15 ? 8'h7c : _GEN_3855; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3857 = 8'h11 == io_state_in_15 ? 8'he3 : _GEN_3856; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3858 = 8'h12 == io_state_in_15 ? 8'h39 : _GEN_3857; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3859 = 8'h13 == io_state_in_15 ? 8'h82 : _GEN_3858; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3860 = 8'h14 == io_state_in_15 ? 8'h9b : _GEN_3859; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3861 = 8'h15 == io_state_in_15 ? 8'h2f : _GEN_3860; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3862 = 8'h16 == io_state_in_15 ? 8'hff : _GEN_3861; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3863 = 8'h17 == io_state_in_15 ? 8'h87 : _GEN_3862; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3864 = 8'h18 == io_state_in_15 ? 8'h34 : _GEN_3863; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3865 = 8'h19 == io_state_in_15 ? 8'h8e : _GEN_3864; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3866 = 8'h1a == io_state_in_15 ? 8'h43 : _GEN_3865; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3867 = 8'h1b == io_state_in_15 ? 8'h44 : _GEN_3866; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3868 = 8'h1c == io_state_in_15 ? 8'hc4 : _GEN_3867; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3869 = 8'h1d == io_state_in_15 ? 8'hde : _GEN_3868; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3870 = 8'h1e == io_state_in_15 ? 8'he9 : _GEN_3869; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3871 = 8'h1f == io_state_in_15 ? 8'hcb : _GEN_3870; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3872 = 8'h20 == io_state_in_15 ? 8'h54 : _GEN_3871; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3873 = 8'h21 == io_state_in_15 ? 8'h7b : _GEN_3872; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3874 = 8'h22 == io_state_in_15 ? 8'h94 : _GEN_3873; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3875 = 8'h23 == io_state_in_15 ? 8'h32 : _GEN_3874; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3876 = 8'h24 == io_state_in_15 ? 8'ha6 : _GEN_3875; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3877 = 8'h25 == io_state_in_15 ? 8'hc2 : _GEN_3876; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3878 = 8'h26 == io_state_in_15 ? 8'h23 : _GEN_3877; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3879 = 8'h27 == io_state_in_15 ? 8'h3d : _GEN_3878; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3880 = 8'h28 == io_state_in_15 ? 8'hee : _GEN_3879; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3881 = 8'h29 == io_state_in_15 ? 8'h4c : _GEN_3880; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3882 = 8'h2a == io_state_in_15 ? 8'h95 : _GEN_3881; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3883 = 8'h2b == io_state_in_15 ? 8'hb : _GEN_3882; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3884 = 8'h2c == io_state_in_15 ? 8'h42 : _GEN_3883; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3885 = 8'h2d == io_state_in_15 ? 8'hfa : _GEN_3884; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3886 = 8'h2e == io_state_in_15 ? 8'hc3 : _GEN_3885; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3887 = 8'h2f == io_state_in_15 ? 8'h4e : _GEN_3886; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3888 = 8'h30 == io_state_in_15 ? 8'h8 : _GEN_3887; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3889 = 8'h31 == io_state_in_15 ? 8'h2e : _GEN_3888; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3890 = 8'h32 == io_state_in_15 ? 8'ha1 : _GEN_3889; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3891 = 8'h33 == io_state_in_15 ? 8'h66 : _GEN_3890; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3892 = 8'h34 == io_state_in_15 ? 8'h28 : _GEN_3891; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3893 = 8'h35 == io_state_in_15 ? 8'hd9 : _GEN_3892; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3894 = 8'h36 == io_state_in_15 ? 8'h24 : _GEN_3893; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3895 = 8'h37 == io_state_in_15 ? 8'hb2 : _GEN_3894; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3896 = 8'h38 == io_state_in_15 ? 8'h76 : _GEN_3895; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3897 = 8'h39 == io_state_in_15 ? 8'h5b : _GEN_3896; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3898 = 8'h3a == io_state_in_15 ? 8'ha2 : _GEN_3897; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3899 = 8'h3b == io_state_in_15 ? 8'h49 : _GEN_3898; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3900 = 8'h3c == io_state_in_15 ? 8'h6d : _GEN_3899; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3901 = 8'h3d == io_state_in_15 ? 8'h8b : _GEN_3900; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3902 = 8'h3e == io_state_in_15 ? 8'hd1 : _GEN_3901; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3903 = 8'h3f == io_state_in_15 ? 8'h25 : _GEN_3902; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3904 = 8'h40 == io_state_in_15 ? 8'h72 : _GEN_3903; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3905 = 8'h41 == io_state_in_15 ? 8'hf8 : _GEN_3904; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3906 = 8'h42 == io_state_in_15 ? 8'hf6 : _GEN_3905; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3907 = 8'h43 == io_state_in_15 ? 8'h64 : _GEN_3906; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3908 = 8'h44 == io_state_in_15 ? 8'h86 : _GEN_3907; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3909 = 8'h45 == io_state_in_15 ? 8'h68 : _GEN_3908; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3910 = 8'h46 == io_state_in_15 ? 8'h98 : _GEN_3909; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3911 = 8'h47 == io_state_in_15 ? 8'h16 : _GEN_3910; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3912 = 8'h48 == io_state_in_15 ? 8'hd4 : _GEN_3911; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3913 = 8'h49 == io_state_in_15 ? 8'ha4 : _GEN_3912; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3914 = 8'h4a == io_state_in_15 ? 8'h5c : _GEN_3913; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3915 = 8'h4b == io_state_in_15 ? 8'hcc : _GEN_3914; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3916 = 8'h4c == io_state_in_15 ? 8'h5d : _GEN_3915; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3917 = 8'h4d == io_state_in_15 ? 8'h65 : _GEN_3916; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3918 = 8'h4e == io_state_in_15 ? 8'hb6 : _GEN_3917; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3919 = 8'h4f == io_state_in_15 ? 8'h92 : _GEN_3918; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3920 = 8'h50 == io_state_in_15 ? 8'h6c : _GEN_3919; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3921 = 8'h51 == io_state_in_15 ? 8'h70 : _GEN_3920; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3922 = 8'h52 == io_state_in_15 ? 8'h48 : _GEN_3921; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3923 = 8'h53 == io_state_in_15 ? 8'h50 : _GEN_3922; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3924 = 8'h54 == io_state_in_15 ? 8'hfd : _GEN_3923; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3925 = 8'h55 == io_state_in_15 ? 8'hed : _GEN_3924; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3926 = 8'h56 == io_state_in_15 ? 8'hb9 : _GEN_3925; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3927 = 8'h57 == io_state_in_15 ? 8'hda : _GEN_3926; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3928 = 8'h58 == io_state_in_15 ? 8'h5e : _GEN_3927; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3929 = 8'h59 == io_state_in_15 ? 8'h15 : _GEN_3928; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3930 = 8'h5a == io_state_in_15 ? 8'h46 : _GEN_3929; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3931 = 8'h5b == io_state_in_15 ? 8'h57 : _GEN_3930; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3932 = 8'h5c == io_state_in_15 ? 8'ha7 : _GEN_3931; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3933 = 8'h5d == io_state_in_15 ? 8'h8d : _GEN_3932; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3934 = 8'h5e == io_state_in_15 ? 8'h9d : _GEN_3933; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3935 = 8'h5f == io_state_in_15 ? 8'h84 : _GEN_3934; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3936 = 8'h60 == io_state_in_15 ? 8'h90 : _GEN_3935; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3937 = 8'h61 == io_state_in_15 ? 8'hd8 : _GEN_3936; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3938 = 8'h62 == io_state_in_15 ? 8'hab : _GEN_3937; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3939 = 8'h63 == io_state_in_15 ? 8'h0 : _GEN_3938; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3940 = 8'h64 == io_state_in_15 ? 8'h8c : _GEN_3939; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3941 = 8'h65 == io_state_in_15 ? 8'hbc : _GEN_3940; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3942 = 8'h66 == io_state_in_15 ? 8'hd3 : _GEN_3941; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3943 = 8'h67 == io_state_in_15 ? 8'ha : _GEN_3942; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3944 = 8'h68 == io_state_in_15 ? 8'hf7 : _GEN_3943; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3945 = 8'h69 == io_state_in_15 ? 8'he4 : _GEN_3944; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3946 = 8'h6a == io_state_in_15 ? 8'h58 : _GEN_3945; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3947 = 8'h6b == io_state_in_15 ? 8'h5 : _GEN_3946; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3948 = 8'h6c == io_state_in_15 ? 8'hb8 : _GEN_3947; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3949 = 8'h6d == io_state_in_15 ? 8'hb3 : _GEN_3948; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3950 = 8'h6e == io_state_in_15 ? 8'h45 : _GEN_3949; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3951 = 8'h6f == io_state_in_15 ? 8'h6 : _GEN_3950; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3952 = 8'h70 == io_state_in_15 ? 8'hd0 : _GEN_3951; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3953 = 8'h71 == io_state_in_15 ? 8'h2c : _GEN_3952; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3954 = 8'h72 == io_state_in_15 ? 8'h1e : _GEN_3953; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3955 = 8'h73 == io_state_in_15 ? 8'h8f : _GEN_3954; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3956 = 8'h74 == io_state_in_15 ? 8'hca : _GEN_3955; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3957 = 8'h75 == io_state_in_15 ? 8'h3f : _GEN_3956; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3958 = 8'h76 == io_state_in_15 ? 8'hf : _GEN_3957; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3959 = 8'h77 == io_state_in_15 ? 8'h2 : _GEN_3958; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3960 = 8'h78 == io_state_in_15 ? 8'hc1 : _GEN_3959; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3961 = 8'h79 == io_state_in_15 ? 8'haf : _GEN_3960; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3962 = 8'h7a == io_state_in_15 ? 8'hbd : _GEN_3961; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3963 = 8'h7b == io_state_in_15 ? 8'h3 : _GEN_3962; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3964 = 8'h7c == io_state_in_15 ? 8'h1 : _GEN_3963; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3965 = 8'h7d == io_state_in_15 ? 8'h13 : _GEN_3964; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3966 = 8'h7e == io_state_in_15 ? 8'h8a : _GEN_3965; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3967 = 8'h7f == io_state_in_15 ? 8'h6b : _GEN_3966; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3968 = 8'h80 == io_state_in_15 ? 8'h3a : _GEN_3967; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3969 = 8'h81 == io_state_in_15 ? 8'h91 : _GEN_3968; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3970 = 8'h82 == io_state_in_15 ? 8'h11 : _GEN_3969; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3971 = 8'h83 == io_state_in_15 ? 8'h41 : _GEN_3970; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3972 = 8'h84 == io_state_in_15 ? 8'h4f : _GEN_3971; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3973 = 8'h85 == io_state_in_15 ? 8'h67 : _GEN_3972; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3974 = 8'h86 == io_state_in_15 ? 8'hdc : _GEN_3973; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3975 = 8'h87 == io_state_in_15 ? 8'hea : _GEN_3974; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3976 = 8'h88 == io_state_in_15 ? 8'h97 : _GEN_3975; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3977 = 8'h89 == io_state_in_15 ? 8'hf2 : _GEN_3976; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3978 = 8'h8a == io_state_in_15 ? 8'hcf : _GEN_3977; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3979 = 8'h8b == io_state_in_15 ? 8'hce : _GEN_3978; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3980 = 8'h8c == io_state_in_15 ? 8'hf0 : _GEN_3979; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3981 = 8'h8d == io_state_in_15 ? 8'hb4 : _GEN_3980; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3982 = 8'h8e == io_state_in_15 ? 8'he6 : _GEN_3981; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3983 = 8'h8f == io_state_in_15 ? 8'h73 : _GEN_3982; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3984 = 8'h90 == io_state_in_15 ? 8'h96 : _GEN_3983; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3985 = 8'h91 == io_state_in_15 ? 8'hac : _GEN_3984; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3986 = 8'h92 == io_state_in_15 ? 8'h74 : _GEN_3985; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3987 = 8'h93 == io_state_in_15 ? 8'h22 : _GEN_3986; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3988 = 8'h94 == io_state_in_15 ? 8'he7 : _GEN_3987; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3989 = 8'h95 == io_state_in_15 ? 8'had : _GEN_3988; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3990 = 8'h96 == io_state_in_15 ? 8'h35 : _GEN_3989; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3991 = 8'h97 == io_state_in_15 ? 8'h85 : _GEN_3990; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3992 = 8'h98 == io_state_in_15 ? 8'he2 : _GEN_3991; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3993 = 8'h99 == io_state_in_15 ? 8'hf9 : _GEN_3992; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3994 = 8'h9a == io_state_in_15 ? 8'h37 : _GEN_3993; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3995 = 8'h9b == io_state_in_15 ? 8'he8 : _GEN_3994; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3996 = 8'h9c == io_state_in_15 ? 8'h1c : _GEN_3995; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3997 = 8'h9d == io_state_in_15 ? 8'h75 : _GEN_3996; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3998 = 8'h9e == io_state_in_15 ? 8'hdf : _GEN_3997; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_3999 = 8'h9f == io_state_in_15 ? 8'h6e : _GEN_3998; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4000 = 8'ha0 == io_state_in_15 ? 8'h47 : _GEN_3999; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4001 = 8'ha1 == io_state_in_15 ? 8'hf1 : _GEN_4000; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4002 = 8'ha2 == io_state_in_15 ? 8'h1a : _GEN_4001; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4003 = 8'ha3 == io_state_in_15 ? 8'h71 : _GEN_4002; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4004 = 8'ha4 == io_state_in_15 ? 8'h1d : _GEN_4003; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4005 = 8'ha5 == io_state_in_15 ? 8'h29 : _GEN_4004; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4006 = 8'ha6 == io_state_in_15 ? 8'hc5 : _GEN_4005; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4007 = 8'ha7 == io_state_in_15 ? 8'h89 : _GEN_4006; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4008 = 8'ha8 == io_state_in_15 ? 8'h6f : _GEN_4007; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4009 = 8'ha9 == io_state_in_15 ? 8'hb7 : _GEN_4008; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4010 = 8'haa == io_state_in_15 ? 8'h62 : _GEN_4009; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4011 = 8'hab == io_state_in_15 ? 8'he : _GEN_4010; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4012 = 8'hac == io_state_in_15 ? 8'haa : _GEN_4011; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4013 = 8'had == io_state_in_15 ? 8'h18 : _GEN_4012; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4014 = 8'hae == io_state_in_15 ? 8'hbe : _GEN_4013; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4015 = 8'haf == io_state_in_15 ? 8'h1b : _GEN_4014; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4016 = 8'hb0 == io_state_in_15 ? 8'hfc : _GEN_4015; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4017 = 8'hb1 == io_state_in_15 ? 8'h56 : _GEN_4016; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4018 = 8'hb2 == io_state_in_15 ? 8'h3e : _GEN_4017; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4019 = 8'hb3 == io_state_in_15 ? 8'h4b : _GEN_4018; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4020 = 8'hb4 == io_state_in_15 ? 8'hc6 : _GEN_4019; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4021 = 8'hb5 == io_state_in_15 ? 8'hd2 : _GEN_4020; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4022 = 8'hb6 == io_state_in_15 ? 8'h79 : _GEN_4021; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4023 = 8'hb7 == io_state_in_15 ? 8'h20 : _GEN_4022; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4024 = 8'hb8 == io_state_in_15 ? 8'h9a : _GEN_4023; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4025 = 8'hb9 == io_state_in_15 ? 8'hdb : _GEN_4024; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4026 = 8'hba == io_state_in_15 ? 8'hc0 : _GEN_4025; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4027 = 8'hbb == io_state_in_15 ? 8'hfe : _GEN_4026; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4028 = 8'hbc == io_state_in_15 ? 8'h78 : _GEN_4027; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4029 = 8'hbd == io_state_in_15 ? 8'hcd : _GEN_4028; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4030 = 8'hbe == io_state_in_15 ? 8'h5a : _GEN_4029; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4031 = 8'hbf == io_state_in_15 ? 8'hf4 : _GEN_4030; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4032 = 8'hc0 == io_state_in_15 ? 8'h1f : _GEN_4031; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4033 = 8'hc1 == io_state_in_15 ? 8'hdd : _GEN_4032; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4034 = 8'hc2 == io_state_in_15 ? 8'ha8 : _GEN_4033; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4035 = 8'hc3 == io_state_in_15 ? 8'h33 : _GEN_4034; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4036 = 8'hc4 == io_state_in_15 ? 8'h88 : _GEN_4035; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4037 = 8'hc5 == io_state_in_15 ? 8'h7 : _GEN_4036; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4038 = 8'hc6 == io_state_in_15 ? 8'hc7 : _GEN_4037; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4039 = 8'hc7 == io_state_in_15 ? 8'h31 : _GEN_4038; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4040 = 8'hc8 == io_state_in_15 ? 8'hb1 : _GEN_4039; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4041 = 8'hc9 == io_state_in_15 ? 8'h12 : _GEN_4040; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4042 = 8'hca == io_state_in_15 ? 8'h10 : _GEN_4041; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4043 = 8'hcb == io_state_in_15 ? 8'h59 : _GEN_4042; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4044 = 8'hcc == io_state_in_15 ? 8'h27 : _GEN_4043; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4045 = 8'hcd == io_state_in_15 ? 8'h80 : _GEN_4044; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4046 = 8'hce == io_state_in_15 ? 8'hec : _GEN_4045; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4047 = 8'hcf == io_state_in_15 ? 8'h5f : _GEN_4046; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4048 = 8'hd0 == io_state_in_15 ? 8'h60 : _GEN_4047; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4049 = 8'hd1 == io_state_in_15 ? 8'h51 : _GEN_4048; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4050 = 8'hd2 == io_state_in_15 ? 8'h7f : _GEN_4049; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4051 = 8'hd3 == io_state_in_15 ? 8'ha9 : _GEN_4050; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4052 = 8'hd4 == io_state_in_15 ? 8'h19 : _GEN_4051; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4053 = 8'hd5 == io_state_in_15 ? 8'hb5 : _GEN_4052; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4054 = 8'hd6 == io_state_in_15 ? 8'h4a : _GEN_4053; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4055 = 8'hd7 == io_state_in_15 ? 8'hd : _GEN_4054; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4056 = 8'hd8 == io_state_in_15 ? 8'h2d : _GEN_4055; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4057 = 8'hd9 == io_state_in_15 ? 8'he5 : _GEN_4056; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4058 = 8'hda == io_state_in_15 ? 8'h7a : _GEN_4057; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4059 = 8'hdb == io_state_in_15 ? 8'h9f : _GEN_4058; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4060 = 8'hdc == io_state_in_15 ? 8'h93 : _GEN_4059; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4061 = 8'hdd == io_state_in_15 ? 8'hc9 : _GEN_4060; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4062 = 8'hde == io_state_in_15 ? 8'h9c : _GEN_4061; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4063 = 8'hdf == io_state_in_15 ? 8'hef : _GEN_4062; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4064 = 8'he0 == io_state_in_15 ? 8'ha0 : _GEN_4063; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4065 = 8'he1 == io_state_in_15 ? 8'he0 : _GEN_4064; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4066 = 8'he2 == io_state_in_15 ? 8'h3b : _GEN_4065; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4067 = 8'he3 == io_state_in_15 ? 8'h4d : _GEN_4066; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4068 = 8'he4 == io_state_in_15 ? 8'hae : _GEN_4067; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4069 = 8'he5 == io_state_in_15 ? 8'h2a : _GEN_4068; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4070 = 8'he6 == io_state_in_15 ? 8'hf5 : _GEN_4069; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4071 = 8'he7 == io_state_in_15 ? 8'hb0 : _GEN_4070; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4072 = 8'he8 == io_state_in_15 ? 8'hc8 : _GEN_4071; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4073 = 8'he9 == io_state_in_15 ? 8'heb : _GEN_4072; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4074 = 8'hea == io_state_in_15 ? 8'hbb : _GEN_4073; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4075 = 8'heb == io_state_in_15 ? 8'h3c : _GEN_4074; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4076 = 8'hec == io_state_in_15 ? 8'h83 : _GEN_4075; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4077 = 8'hed == io_state_in_15 ? 8'h53 : _GEN_4076; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4078 = 8'hee == io_state_in_15 ? 8'h99 : _GEN_4077; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4079 = 8'hef == io_state_in_15 ? 8'h61 : _GEN_4078; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4080 = 8'hf0 == io_state_in_15 ? 8'h17 : _GEN_4079; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4081 = 8'hf1 == io_state_in_15 ? 8'h2b : _GEN_4080; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4082 = 8'hf2 == io_state_in_15 ? 8'h4 : _GEN_4081; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4083 = 8'hf3 == io_state_in_15 ? 8'h7e : _GEN_4082; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4084 = 8'hf4 == io_state_in_15 ? 8'hba : _GEN_4083; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4085 = 8'hf5 == io_state_in_15 ? 8'h77 : _GEN_4084; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4086 = 8'hf6 == io_state_in_15 ? 8'hd6 : _GEN_4085; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4087 = 8'hf7 == io_state_in_15 ? 8'h26 : _GEN_4086; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4088 = 8'hf8 == io_state_in_15 ? 8'he1 : _GEN_4087; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4089 = 8'hf9 == io_state_in_15 ? 8'h69 : _GEN_4088; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4090 = 8'hfa == io_state_in_15 ? 8'h14 : _GEN_4089; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4091 = 8'hfb == io_state_in_15 ? 8'h63 : _GEN_4090; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4092 = 8'hfc == io_state_in_15 ? 8'h55 : _GEN_4091; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4093 = 8'hfd == io_state_in_15 ? 8'h21 : _GEN_4092; // @[InvSubBytes.scala 36:{23,23}]
  wire [7:0] _GEN_4094 = 8'hfe == io_state_in_15 ? 8'hc : _GEN_4093; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_0 = 8'hff == io_state_in_0 ? 8'h7d : _GEN_254; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_1 = 8'hff == io_state_in_1 ? 8'h7d : _GEN_510; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_2 = 8'hff == io_state_in_2 ? 8'h7d : _GEN_766; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_3 = 8'hff == io_state_in_3 ? 8'h7d : _GEN_1022; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_4 = 8'hff == io_state_in_4 ? 8'h7d : _GEN_1278; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_5 = 8'hff == io_state_in_5 ? 8'h7d : _GEN_1534; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_6 = 8'hff == io_state_in_6 ? 8'h7d : _GEN_1790; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_7 = 8'hff == io_state_in_7 ? 8'h7d : _GEN_2046; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_8 = 8'hff == io_state_in_8 ? 8'h7d : _GEN_2302; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_9 = 8'hff == io_state_in_9 ? 8'h7d : _GEN_2558; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_10 = 8'hff == io_state_in_10 ? 8'h7d : _GEN_2814; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_11 = 8'hff == io_state_in_11 ? 8'h7d : _GEN_3070; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_12 = 8'hff == io_state_in_12 ? 8'h7d : _GEN_3326; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_13 = 8'hff == io_state_in_13 ? 8'h7d : _GEN_3582; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_14 = 8'hff == io_state_in_14 ? 8'h7d : _GEN_3838; // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_15 = 8'hff == io_state_in_15 ? 8'h7d : _GEN_4094; // @[InvSubBytes.scala 36:{23,23}]
endmodule
module InvShiftRows(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  assign io_state_out_0 = io_state_in_0; // @[InvShiftRows.scala 13:19]
  assign io_state_out_1 = io_state_in_13; // @[InvShiftRows.scala 14:19]
  assign io_state_out_2 = io_state_in_10; // @[InvShiftRows.scala 15:19]
  assign io_state_out_3 = io_state_in_7; // @[InvShiftRows.scala 16:19]
  assign io_state_out_4 = io_state_in_4; // @[InvShiftRows.scala 18:19]
  assign io_state_out_5 = io_state_in_1; // @[InvShiftRows.scala 19:19]
  assign io_state_out_6 = io_state_in_14; // @[InvShiftRows.scala 20:19]
  assign io_state_out_7 = io_state_in_11; // @[InvShiftRows.scala 21:19]
  assign io_state_out_8 = io_state_in_8; // @[InvShiftRows.scala 23:19]
  assign io_state_out_9 = io_state_in_5; // @[InvShiftRows.scala 24:19]
  assign io_state_out_10 = io_state_in_2; // @[InvShiftRows.scala 25:20]
  assign io_state_out_11 = io_state_in_15; // @[InvShiftRows.scala 26:20]
  assign io_state_out_12 = io_state_in_12; // @[InvShiftRows.scala 28:20]
  assign io_state_out_13 = io_state_in_9; // @[InvShiftRows.scala 29:20]
  assign io_state_out_14 = io_state_in_6; // @[InvShiftRows.scala 30:20]
  assign io_state_out_15 = io_state_in_3; // @[InvShiftRows.scala 31:20]
endmodule
module InvMixColumns(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  wire [7:0] _GEN_1 = 8'h1 == io_state_in_0 ? 8'he : 8'h0; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_2 = 8'h2 == io_state_in_0 ? 8'h1c : _GEN_1; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_3 = 8'h3 == io_state_in_0 ? 8'h12 : _GEN_2; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_4 = 8'h4 == io_state_in_0 ? 8'h38 : _GEN_3; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_5 = 8'h5 == io_state_in_0 ? 8'h36 : _GEN_4; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_6 = 8'h6 == io_state_in_0 ? 8'h24 : _GEN_5; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_7 = 8'h7 == io_state_in_0 ? 8'h2a : _GEN_6; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_8 = 8'h8 == io_state_in_0 ? 8'h70 : _GEN_7; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_9 = 8'h9 == io_state_in_0 ? 8'h7e : _GEN_8; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_10 = 8'ha == io_state_in_0 ? 8'h6c : _GEN_9; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_11 = 8'hb == io_state_in_0 ? 8'h62 : _GEN_10; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_12 = 8'hc == io_state_in_0 ? 8'h48 : _GEN_11; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_13 = 8'hd == io_state_in_0 ? 8'h46 : _GEN_12; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_14 = 8'he == io_state_in_0 ? 8'h54 : _GEN_13; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_15 = 8'hf == io_state_in_0 ? 8'h5a : _GEN_14; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_16 = 8'h10 == io_state_in_0 ? 8'he0 : _GEN_15; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_17 = 8'h11 == io_state_in_0 ? 8'hee : _GEN_16; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_18 = 8'h12 == io_state_in_0 ? 8'hfc : _GEN_17; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_19 = 8'h13 == io_state_in_0 ? 8'hf2 : _GEN_18; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_20 = 8'h14 == io_state_in_0 ? 8'hd8 : _GEN_19; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_21 = 8'h15 == io_state_in_0 ? 8'hd6 : _GEN_20; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_22 = 8'h16 == io_state_in_0 ? 8'hc4 : _GEN_21; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_23 = 8'h17 == io_state_in_0 ? 8'hca : _GEN_22; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_24 = 8'h18 == io_state_in_0 ? 8'h90 : _GEN_23; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_25 = 8'h19 == io_state_in_0 ? 8'h9e : _GEN_24; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_26 = 8'h1a == io_state_in_0 ? 8'h8c : _GEN_25; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_27 = 8'h1b == io_state_in_0 ? 8'h82 : _GEN_26; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_28 = 8'h1c == io_state_in_0 ? 8'ha8 : _GEN_27; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_29 = 8'h1d == io_state_in_0 ? 8'ha6 : _GEN_28; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_30 = 8'h1e == io_state_in_0 ? 8'hb4 : _GEN_29; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_31 = 8'h1f == io_state_in_0 ? 8'hba : _GEN_30; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_32 = 8'h20 == io_state_in_0 ? 8'hdb : _GEN_31; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_33 = 8'h21 == io_state_in_0 ? 8'hd5 : _GEN_32; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_34 = 8'h22 == io_state_in_0 ? 8'hc7 : _GEN_33; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_35 = 8'h23 == io_state_in_0 ? 8'hc9 : _GEN_34; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_36 = 8'h24 == io_state_in_0 ? 8'he3 : _GEN_35; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_37 = 8'h25 == io_state_in_0 ? 8'hed : _GEN_36; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_38 = 8'h26 == io_state_in_0 ? 8'hff : _GEN_37; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_39 = 8'h27 == io_state_in_0 ? 8'hf1 : _GEN_38; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_40 = 8'h28 == io_state_in_0 ? 8'hab : _GEN_39; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_41 = 8'h29 == io_state_in_0 ? 8'ha5 : _GEN_40; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_42 = 8'h2a == io_state_in_0 ? 8'hb7 : _GEN_41; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_43 = 8'h2b == io_state_in_0 ? 8'hb9 : _GEN_42; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_44 = 8'h2c == io_state_in_0 ? 8'h93 : _GEN_43; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_45 = 8'h2d == io_state_in_0 ? 8'h9d : _GEN_44; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_46 = 8'h2e == io_state_in_0 ? 8'h8f : _GEN_45; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_47 = 8'h2f == io_state_in_0 ? 8'h81 : _GEN_46; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_48 = 8'h30 == io_state_in_0 ? 8'h3b : _GEN_47; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_49 = 8'h31 == io_state_in_0 ? 8'h35 : _GEN_48; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_50 = 8'h32 == io_state_in_0 ? 8'h27 : _GEN_49; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_51 = 8'h33 == io_state_in_0 ? 8'h29 : _GEN_50; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_52 = 8'h34 == io_state_in_0 ? 8'h3 : _GEN_51; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_53 = 8'h35 == io_state_in_0 ? 8'hd : _GEN_52; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_54 = 8'h36 == io_state_in_0 ? 8'h1f : _GEN_53; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_55 = 8'h37 == io_state_in_0 ? 8'h11 : _GEN_54; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_56 = 8'h38 == io_state_in_0 ? 8'h4b : _GEN_55; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_57 = 8'h39 == io_state_in_0 ? 8'h45 : _GEN_56; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_58 = 8'h3a == io_state_in_0 ? 8'h57 : _GEN_57; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_59 = 8'h3b == io_state_in_0 ? 8'h59 : _GEN_58; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_60 = 8'h3c == io_state_in_0 ? 8'h73 : _GEN_59; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_61 = 8'h3d == io_state_in_0 ? 8'h7d : _GEN_60; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_62 = 8'h3e == io_state_in_0 ? 8'h6f : _GEN_61; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_63 = 8'h3f == io_state_in_0 ? 8'h61 : _GEN_62; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_64 = 8'h40 == io_state_in_0 ? 8'had : _GEN_63; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_65 = 8'h41 == io_state_in_0 ? 8'ha3 : _GEN_64; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_66 = 8'h42 == io_state_in_0 ? 8'hb1 : _GEN_65; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_67 = 8'h43 == io_state_in_0 ? 8'hbf : _GEN_66; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_68 = 8'h44 == io_state_in_0 ? 8'h95 : _GEN_67; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_69 = 8'h45 == io_state_in_0 ? 8'h9b : _GEN_68; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_70 = 8'h46 == io_state_in_0 ? 8'h89 : _GEN_69; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_71 = 8'h47 == io_state_in_0 ? 8'h87 : _GEN_70; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_72 = 8'h48 == io_state_in_0 ? 8'hdd : _GEN_71; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_73 = 8'h49 == io_state_in_0 ? 8'hd3 : _GEN_72; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_74 = 8'h4a == io_state_in_0 ? 8'hc1 : _GEN_73; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_75 = 8'h4b == io_state_in_0 ? 8'hcf : _GEN_74; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_76 = 8'h4c == io_state_in_0 ? 8'he5 : _GEN_75; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_77 = 8'h4d == io_state_in_0 ? 8'heb : _GEN_76; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_78 = 8'h4e == io_state_in_0 ? 8'hf9 : _GEN_77; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_79 = 8'h4f == io_state_in_0 ? 8'hf7 : _GEN_78; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_80 = 8'h50 == io_state_in_0 ? 8'h4d : _GEN_79; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_81 = 8'h51 == io_state_in_0 ? 8'h43 : _GEN_80; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_82 = 8'h52 == io_state_in_0 ? 8'h51 : _GEN_81; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_83 = 8'h53 == io_state_in_0 ? 8'h5f : _GEN_82; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_84 = 8'h54 == io_state_in_0 ? 8'h75 : _GEN_83; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_85 = 8'h55 == io_state_in_0 ? 8'h7b : _GEN_84; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_86 = 8'h56 == io_state_in_0 ? 8'h69 : _GEN_85; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_87 = 8'h57 == io_state_in_0 ? 8'h67 : _GEN_86; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_88 = 8'h58 == io_state_in_0 ? 8'h3d : _GEN_87; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_89 = 8'h59 == io_state_in_0 ? 8'h33 : _GEN_88; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_90 = 8'h5a == io_state_in_0 ? 8'h21 : _GEN_89; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_91 = 8'h5b == io_state_in_0 ? 8'h2f : _GEN_90; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_92 = 8'h5c == io_state_in_0 ? 8'h5 : _GEN_91; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_93 = 8'h5d == io_state_in_0 ? 8'hb : _GEN_92; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_94 = 8'h5e == io_state_in_0 ? 8'h19 : _GEN_93; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_95 = 8'h5f == io_state_in_0 ? 8'h17 : _GEN_94; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_96 = 8'h60 == io_state_in_0 ? 8'h76 : _GEN_95; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_97 = 8'h61 == io_state_in_0 ? 8'h78 : _GEN_96; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_98 = 8'h62 == io_state_in_0 ? 8'h6a : _GEN_97; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_99 = 8'h63 == io_state_in_0 ? 8'h64 : _GEN_98; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_100 = 8'h64 == io_state_in_0 ? 8'h4e : _GEN_99; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_101 = 8'h65 == io_state_in_0 ? 8'h40 : _GEN_100; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_102 = 8'h66 == io_state_in_0 ? 8'h52 : _GEN_101; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_103 = 8'h67 == io_state_in_0 ? 8'h5c : _GEN_102; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_104 = 8'h68 == io_state_in_0 ? 8'h6 : _GEN_103; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_105 = 8'h69 == io_state_in_0 ? 8'h8 : _GEN_104; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_106 = 8'h6a == io_state_in_0 ? 8'h1a : _GEN_105; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_107 = 8'h6b == io_state_in_0 ? 8'h14 : _GEN_106; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_108 = 8'h6c == io_state_in_0 ? 8'h3e : _GEN_107; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_109 = 8'h6d == io_state_in_0 ? 8'h30 : _GEN_108; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_110 = 8'h6e == io_state_in_0 ? 8'h22 : _GEN_109; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_111 = 8'h6f == io_state_in_0 ? 8'h2c : _GEN_110; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_112 = 8'h70 == io_state_in_0 ? 8'h96 : _GEN_111; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_113 = 8'h71 == io_state_in_0 ? 8'h98 : _GEN_112; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_114 = 8'h72 == io_state_in_0 ? 8'h8a : _GEN_113; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_115 = 8'h73 == io_state_in_0 ? 8'h84 : _GEN_114; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_116 = 8'h74 == io_state_in_0 ? 8'hae : _GEN_115; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_117 = 8'h75 == io_state_in_0 ? 8'ha0 : _GEN_116; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_118 = 8'h76 == io_state_in_0 ? 8'hb2 : _GEN_117; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_119 = 8'h77 == io_state_in_0 ? 8'hbc : _GEN_118; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_120 = 8'h78 == io_state_in_0 ? 8'he6 : _GEN_119; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_121 = 8'h79 == io_state_in_0 ? 8'he8 : _GEN_120; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_122 = 8'h7a == io_state_in_0 ? 8'hfa : _GEN_121; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_123 = 8'h7b == io_state_in_0 ? 8'hf4 : _GEN_122; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_124 = 8'h7c == io_state_in_0 ? 8'hde : _GEN_123; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_125 = 8'h7d == io_state_in_0 ? 8'hd0 : _GEN_124; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_126 = 8'h7e == io_state_in_0 ? 8'hc2 : _GEN_125; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_127 = 8'h7f == io_state_in_0 ? 8'hcc : _GEN_126; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_128 = 8'h80 == io_state_in_0 ? 8'h41 : _GEN_127; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_129 = 8'h81 == io_state_in_0 ? 8'h4f : _GEN_128; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_130 = 8'h82 == io_state_in_0 ? 8'h5d : _GEN_129; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_131 = 8'h83 == io_state_in_0 ? 8'h53 : _GEN_130; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_132 = 8'h84 == io_state_in_0 ? 8'h79 : _GEN_131; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_133 = 8'h85 == io_state_in_0 ? 8'h77 : _GEN_132; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_134 = 8'h86 == io_state_in_0 ? 8'h65 : _GEN_133; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_135 = 8'h87 == io_state_in_0 ? 8'h6b : _GEN_134; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_136 = 8'h88 == io_state_in_0 ? 8'h31 : _GEN_135; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_137 = 8'h89 == io_state_in_0 ? 8'h3f : _GEN_136; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_138 = 8'h8a == io_state_in_0 ? 8'h2d : _GEN_137; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_139 = 8'h8b == io_state_in_0 ? 8'h23 : _GEN_138; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_140 = 8'h8c == io_state_in_0 ? 8'h9 : _GEN_139; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_141 = 8'h8d == io_state_in_0 ? 8'h7 : _GEN_140; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_142 = 8'h8e == io_state_in_0 ? 8'h15 : _GEN_141; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_143 = 8'h8f == io_state_in_0 ? 8'h1b : _GEN_142; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_144 = 8'h90 == io_state_in_0 ? 8'ha1 : _GEN_143; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_145 = 8'h91 == io_state_in_0 ? 8'haf : _GEN_144; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_146 = 8'h92 == io_state_in_0 ? 8'hbd : _GEN_145; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_147 = 8'h93 == io_state_in_0 ? 8'hb3 : _GEN_146; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_148 = 8'h94 == io_state_in_0 ? 8'h99 : _GEN_147; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_149 = 8'h95 == io_state_in_0 ? 8'h97 : _GEN_148; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_150 = 8'h96 == io_state_in_0 ? 8'h85 : _GEN_149; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_151 = 8'h97 == io_state_in_0 ? 8'h8b : _GEN_150; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_152 = 8'h98 == io_state_in_0 ? 8'hd1 : _GEN_151; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_153 = 8'h99 == io_state_in_0 ? 8'hdf : _GEN_152; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_154 = 8'h9a == io_state_in_0 ? 8'hcd : _GEN_153; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_155 = 8'h9b == io_state_in_0 ? 8'hc3 : _GEN_154; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_156 = 8'h9c == io_state_in_0 ? 8'he9 : _GEN_155; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_157 = 8'h9d == io_state_in_0 ? 8'he7 : _GEN_156; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_158 = 8'h9e == io_state_in_0 ? 8'hf5 : _GEN_157; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_159 = 8'h9f == io_state_in_0 ? 8'hfb : _GEN_158; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_160 = 8'ha0 == io_state_in_0 ? 8'h9a : _GEN_159; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_161 = 8'ha1 == io_state_in_0 ? 8'h94 : _GEN_160; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_162 = 8'ha2 == io_state_in_0 ? 8'h86 : _GEN_161; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_163 = 8'ha3 == io_state_in_0 ? 8'h88 : _GEN_162; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_164 = 8'ha4 == io_state_in_0 ? 8'ha2 : _GEN_163; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_165 = 8'ha5 == io_state_in_0 ? 8'hac : _GEN_164; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_166 = 8'ha6 == io_state_in_0 ? 8'hbe : _GEN_165; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_167 = 8'ha7 == io_state_in_0 ? 8'hb0 : _GEN_166; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_168 = 8'ha8 == io_state_in_0 ? 8'hea : _GEN_167; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_169 = 8'ha9 == io_state_in_0 ? 8'he4 : _GEN_168; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_170 = 8'haa == io_state_in_0 ? 8'hf6 : _GEN_169; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_171 = 8'hab == io_state_in_0 ? 8'hf8 : _GEN_170; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_172 = 8'hac == io_state_in_0 ? 8'hd2 : _GEN_171; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_173 = 8'had == io_state_in_0 ? 8'hdc : _GEN_172; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_174 = 8'hae == io_state_in_0 ? 8'hce : _GEN_173; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_175 = 8'haf == io_state_in_0 ? 8'hc0 : _GEN_174; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_176 = 8'hb0 == io_state_in_0 ? 8'h7a : _GEN_175; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_177 = 8'hb1 == io_state_in_0 ? 8'h74 : _GEN_176; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_178 = 8'hb2 == io_state_in_0 ? 8'h66 : _GEN_177; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_179 = 8'hb3 == io_state_in_0 ? 8'h68 : _GEN_178; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_180 = 8'hb4 == io_state_in_0 ? 8'h42 : _GEN_179; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_181 = 8'hb5 == io_state_in_0 ? 8'h4c : _GEN_180; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_182 = 8'hb6 == io_state_in_0 ? 8'h5e : _GEN_181; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_183 = 8'hb7 == io_state_in_0 ? 8'h50 : _GEN_182; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_184 = 8'hb8 == io_state_in_0 ? 8'ha : _GEN_183; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_185 = 8'hb9 == io_state_in_0 ? 8'h4 : _GEN_184; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_186 = 8'hba == io_state_in_0 ? 8'h16 : _GEN_185; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_187 = 8'hbb == io_state_in_0 ? 8'h18 : _GEN_186; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_188 = 8'hbc == io_state_in_0 ? 8'h32 : _GEN_187; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_189 = 8'hbd == io_state_in_0 ? 8'h3c : _GEN_188; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_190 = 8'hbe == io_state_in_0 ? 8'h2e : _GEN_189; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_191 = 8'hbf == io_state_in_0 ? 8'h20 : _GEN_190; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_192 = 8'hc0 == io_state_in_0 ? 8'hec : _GEN_191; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_193 = 8'hc1 == io_state_in_0 ? 8'he2 : _GEN_192; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_194 = 8'hc2 == io_state_in_0 ? 8'hf0 : _GEN_193; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_195 = 8'hc3 == io_state_in_0 ? 8'hfe : _GEN_194; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_196 = 8'hc4 == io_state_in_0 ? 8'hd4 : _GEN_195; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_197 = 8'hc5 == io_state_in_0 ? 8'hda : _GEN_196; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_198 = 8'hc6 == io_state_in_0 ? 8'hc8 : _GEN_197; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_199 = 8'hc7 == io_state_in_0 ? 8'hc6 : _GEN_198; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_200 = 8'hc8 == io_state_in_0 ? 8'h9c : _GEN_199; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_201 = 8'hc9 == io_state_in_0 ? 8'h92 : _GEN_200; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_202 = 8'hca == io_state_in_0 ? 8'h80 : _GEN_201; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_203 = 8'hcb == io_state_in_0 ? 8'h8e : _GEN_202; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_204 = 8'hcc == io_state_in_0 ? 8'ha4 : _GEN_203; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_205 = 8'hcd == io_state_in_0 ? 8'haa : _GEN_204; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_206 = 8'hce == io_state_in_0 ? 8'hb8 : _GEN_205; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_207 = 8'hcf == io_state_in_0 ? 8'hb6 : _GEN_206; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_208 = 8'hd0 == io_state_in_0 ? 8'hc : _GEN_207; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_209 = 8'hd1 == io_state_in_0 ? 8'h2 : _GEN_208; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_210 = 8'hd2 == io_state_in_0 ? 8'h10 : _GEN_209; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_211 = 8'hd3 == io_state_in_0 ? 8'h1e : _GEN_210; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_212 = 8'hd4 == io_state_in_0 ? 8'h34 : _GEN_211; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_213 = 8'hd5 == io_state_in_0 ? 8'h3a : _GEN_212; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_214 = 8'hd6 == io_state_in_0 ? 8'h28 : _GEN_213; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_215 = 8'hd7 == io_state_in_0 ? 8'h26 : _GEN_214; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_216 = 8'hd8 == io_state_in_0 ? 8'h7c : _GEN_215; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_217 = 8'hd9 == io_state_in_0 ? 8'h72 : _GEN_216; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_218 = 8'hda == io_state_in_0 ? 8'h60 : _GEN_217; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_219 = 8'hdb == io_state_in_0 ? 8'h6e : _GEN_218; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_220 = 8'hdc == io_state_in_0 ? 8'h44 : _GEN_219; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_221 = 8'hdd == io_state_in_0 ? 8'h4a : _GEN_220; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_222 = 8'hde == io_state_in_0 ? 8'h58 : _GEN_221; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_223 = 8'hdf == io_state_in_0 ? 8'h56 : _GEN_222; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_224 = 8'he0 == io_state_in_0 ? 8'h37 : _GEN_223; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_225 = 8'he1 == io_state_in_0 ? 8'h39 : _GEN_224; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_226 = 8'he2 == io_state_in_0 ? 8'h2b : _GEN_225; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_227 = 8'he3 == io_state_in_0 ? 8'h25 : _GEN_226; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_228 = 8'he4 == io_state_in_0 ? 8'hf : _GEN_227; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_229 = 8'he5 == io_state_in_0 ? 8'h1 : _GEN_228; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_230 = 8'he6 == io_state_in_0 ? 8'h13 : _GEN_229; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_231 = 8'he7 == io_state_in_0 ? 8'h1d : _GEN_230; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_232 = 8'he8 == io_state_in_0 ? 8'h47 : _GEN_231; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_233 = 8'he9 == io_state_in_0 ? 8'h49 : _GEN_232; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_234 = 8'hea == io_state_in_0 ? 8'h5b : _GEN_233; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_235 = 8'heb == io_state_in_0 ? 8'h55 : _GEN_234; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_236 = 8'hec == io_state_in_0 ? 8'h7f : _GEN_235; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_237 = 8'hed == io_state_in_0 ? 8'h71 : _GEN_236; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_238 = 8'hee == io_state_in_0 ? 8'h63 : _GEN_237; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_239 = 8'hef == io_state_in_0 ? 8'h6d : _GEN_238; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_240 = 8'hf0 == io_state_in_0 ? 8'hd7 : _GEN_239; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_241 = 8'hf1 == io_state_in_0 ? 8'hd9 : _GEN_240; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_242 = 8'hf2 == io_state_in_0 ? 8'hcb : _GEN_241; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_243 = 8'hf3 == io_state_in_0 ? 8'hc5 : _GEN_242; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_244 = 8'hf4 == io_state_in_0 ? 8'hef : _GEN_243; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_245 = 8'hf5 == io_state_in_0 ? 8'he1 : _GEN_244; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_246 = 8'hf6 == io_state_in_0 ? 8'hf3 : _GEN_245; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_247 = 8'hf7 == io_state_in_0 ? 8'hfd : _GEN_246; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_248 = 8'hf8 == io_state_in_0 ? 8'ha7 : _GEN_247; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_249 = 8'hf9 == io_state_in_0 ? 8'ha9 : _GEN_248; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_250 = 8'hfa == io_state_in_0 ? 8'hbb : _GEN_249; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_251 = 8'hfb == io_state_in_0 ? 8'hb5 : _GEN_250; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_252 = 8'hfc == io_state_in_0 ? 8'h9f : _GEN_251; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_253 = 8'hfd == io_state_in_0 ? 8'h91 : _GEN_252; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_254 = 8'hfe == io_state_in_0 ? 8'h83 : _GEN_253; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_255 = 8'hff == io_state_in_0 ? 8'h8d : _GEN_254; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_257 = 8'h1 == io_state_in_1 ? 8'hb : 8'h0; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_258 = 8'h2 == io_state_in_1 ? 8'h16 : _GEN_257; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_259 = 8'h3 == io_state_in_1 ? 8'h1d : _GEN_258; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_260 = 8'h4 == io_state_in_1 ? 8'h2c : _GEN_259; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_261 = 8'h5 == io_state_in_1 ? 8'h27 : _GEN_260; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_262 = 8'h6 == io_state_in_1 ? 8'h3a : _GEN_261; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_263 = 8'h7 == io_state_in_1 ? 8'h31 : _GEN_262; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_264 = 8'h8 == io_state_in_1 ? 8'h58 : _GEN_263; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_265 = 8'h9 == io_state_in_1 ? 8'h53 : _GEN_264; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_266 = 8'ha == io_state_in_1 ? 8'h4e : _GEN_265; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_267 = 8'hb == io_state_in_1 ? 8'h45 : _GEN_266; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_268 = 8'hc == io_state_in_1 ? 8'h74 : _GEN_267; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_269 = 8'hd == io_state_in_1 ? 8'h7f : _GEN_268; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_270 = 8'he == io_state_in_1 ? 8'h62 : _GEN_269; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_271 = 8'hf == io_state_in_1 ? 8'h69 : _GEN_270; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_272 = 8'h10 == io_state_in_1 ? 8'hb0 : _GEN_271; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_273 = 8'h11 == io_state_in_1 ? 8'hbb : _GEN_272; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_274 = 8'h12 == io_state_in_1 ? 8'ha6 : _GEN_273; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_275 = 8'h13 == io_state_in_1 ? 8'had : _GEN_274; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_276 = 8'h14 == io_state_in_1 ? 8'h9c : _GEN_275; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_277 = 8'h15 == io_state_in_1 ? 8'h97 : _GEN_276; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_278 = 8'h16 == io_state_in_1 ? 8'h8a : _GEN_277; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_279 = 8'h17 == io_state_in_1 ? 8'h81 : _GEN_278; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_280 = 8'h18 == io_state_in_1 ? 8'he8 : _GEN_279; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_281 = 8'h19 == io_state_in_1 ? 8'he3 : _GEN_280; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_282 = 8'h1a == io_state_in_1 ? 8'hfe : _GEN_281; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_283 = 8'h1b == io_state_in_1 ? 8'hf5 : _GEN_282; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_284 = 8'h1c == io_state_in_1 ? 8'hc4 : _GEN_283; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_285 = 8'h1d == io_state_in_1 ? 8'hcf : _GEN_284; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_286 = 8'h1e == io_state_in_1 ? 8'hd2 : _GEN_285; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_287 = 8'h1f == io_state_in_1 ? 8'hd9 : _GEN_286; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_288 = 8'h20 == io_state_in_1 ? 8'h7b : _GEN_287; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_289 = 8'h21 == io_state_in_1 ? 8'h70 : _GEN_288; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_290 = 8'h22 == io_state_in_1 ? 8'h6d : _GEN_289; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_291 = 8'h23 == io_state_in_1 ? 8'h66 : _GEN_290; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_292 = 8'h24 == io_state_in_1 ? 8'h57 : _GEN_291; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_293 = 8'h25 == io_state_in_1 ? 8'h5c : _GEN_292; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_294 = 8'h26 == io_state_in_1 ? 8'h41 : _GEN_293; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_295 = 8'h27 == io_state_in_1 ? 8'h4a : _GEN_294; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_296 = 8'h28 == io_state_in_1 ? 8'h23 : _GEN_295; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_297 = 8'h29 == io_state_in_1 ? 8'h28 : _GEN_296; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_298 = 8'h2a == io_state_in_1 ? 8'h35 : _GEN_297; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_299 = 8'h2b == io_state_in_1 ? 8'h3e : _GEN_298; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_300 = 8'h2c == io_state_in_1 ? 8'hf : _GEN_299; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_301 = 8'h2d == io_state_in_1 ? 8'h4 : _GEN_300; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_302 = 8'h2e == io_state_in_1 ? 8'h19 : _GEN_301; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_303 = 8'h2f == io_state_in_1 ? 8'h12 : _GEN_302; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_304 = 8'h30 == io_state_in_1 ? 8'hcb : _GEN_303; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_305 = 8'h31 == io_state_in_1 ? 8'hc0 : _GEN_304; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_306 = 8'h32 == io_state_in_1 ? 8'hdd : _GEN_305; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_307 = 8'h33 == io_state_in_1 ? 8'hd6 : _GEN_306; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_308 = 8'h34 == io_state_in_1 ? 8'he7 : _GEN_307; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_309 = 8'h35 == io_state_in_1 ? 8'hec : _GEN_308; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_310 = 8'h36 == io_state_in_1 ? 8'hf1 : _GEN_309; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_311 = 8'h37 == io_state_in_1 ? 8'hfa : _GEN_310; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_312 = 8'h38 == io_state_in_1 ? 8'h93 : _GEN_311; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_313 = 8'h39 == io_state_in_1 ? 8'h98 : _GEN_312; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_314 = 8'h3a == io_state_in_1 ? 8'h85 : _GEN_313; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_315 = 8'h3b == io_state_in_1 ? 8'h8e : _GEN_314; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_316 = 8'h3c == io_state_in_1 ? 8'hbf : _GEN_315; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_317 = 8'h3d == io_state_in_1 ? 8'hb4 : _GEN_316; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_318 = 8'h3e == io_state_in_1 ? 8'ha9 : _GEN_317; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_319 = 8'h3f == io_state_in_1 ? 8'ha2 : _GEN_318; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_320 = 8'h40 == io_state_in_1 ? 8'hf6 : _GEN_319; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_321 = 8'h41 == io_state_in_1 ? 8'hfd : _GEN_320; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_322 = 8'h42 == io_state_in_1 ? 8'he0 : _GEN_321; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_323 = 8'h43 == io_state_in_1 ? 8'heb : _GEN_322; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_324 = 8'h44 == io_state_in_1 ? 8'hda : _GEN_323; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_325 = 8'h45 == io_state_in_1 ? 8'hd1 : _GEN_324; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_326 = 8'h46 == io_state_in_1 ? 8'hcc : _GEN_325; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_327 = 8'h47 == io_state_in_1 ? 8'hc7 : _GEN_326; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_328 = 8'h48 == io_state_in_1 ? 8'hae : _GEN_327; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_329 = 8'h49 == io_state_in_1 ? 8'ha5 : _GEN_328; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_330 = 8'h4a == io_state_in_1 ? 8'hb8 : _GEN_329; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_331 = 8'h4b == io_state_in_1 ? 8'hb3 : _GEN_330; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_332 = 8'h4c == io_state_in_1 ? 8'h82 : _GEN_331; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_333 = 8'h4d == io_state_in_1 ? 8'h89 : _GEN_332; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_334 = 8'h4e == io_state_in_1 ? 8'h94 : _GEN_333; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_335 = 8'h4f == io_state_in_1 ? 8'h9f : _GEN_334; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_336 = 8'h50 == io_state_in_1 ? 8'h46 : _GEN_335; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_337 = 8'h51 == io_state_in_1 ? 8'h4d : _GEN_336; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_338 = 8'h52 == io_state_in_1 ? 8'h50 : _GEN_337; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_339 = 8'h53 == io_state_in_1 ? 8'h5b : _GEN_338; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_340 = 8'h54 == io_state_in_1 ? 8'h6a : _GEN_339; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_341 = 8'h55 == io_state_in_1 ? 8'h61 : _GEN_340; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_342 = 8'h56 == io_state_in_1 ? 8'h7c : _GEN_341; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_343 = 8'h57 == io_state_in_1 ? 8'h77 : _GEN_342; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_344 = 8'h58 == io_state_in_1 ? 8'h1e : _GEN_343; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_345 = 8'h59 == io_state_in_1 ? 8'h15 : _GEN_344; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_346 = 8'h5a == io_state_in_1 ? 8'h8 : _GEN_345; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_347 = 8'h5b == io_state_in_1 ? 8'h3 : _GEN_346; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_348 = 8'h5c == io_state_in_1 ? 8'h32 : _GEN_347; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_349 = 8'h5d == io_state_in_1 ? 8'h39 : _GEN_348; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_350 = 8'h5e == io_state_in_1 ? 8'h24 : _GEN_349; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_351 = 8'h5f == io_state_in_1 ? 8'h2f : _GEN_350; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_352 = 8'h60 == io_state_in_1 ? 8'h8d : _GEN_351; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_353 = 8'h61 == io_state_in_1 ? 8'h86 : _GEN_352; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_354 = 8'h62 == io_state_in_1 ? 8'h9b : _GEN_353; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_355 = 8'h63 == io_state_in_1 ? 8'h90 : _GEN_354; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_356 = 8'h64 == io_state_in_1 ? 8'ha1 : _GEN_355; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_357 = 8'h65 == io_state_in_1 ? 8'haa : _GEN_356; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_358 = 8'h66 == io_state_in_1 ? 8'hb7 : _GEN_357; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_359 = 8'h67 == io_state_in_1 ? 8'hbc : _GEN_358; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_360 = 8'h68 == io_state_in_1 ? 8'hd5 : _GEN_359; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_361 = 8'h69 == io_state_in_1 ? 8'hde : _GEN_360; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_362 = 8'h6a == io_state_in_1 ? 8'hc3 : _GEN_361; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_363 = 8'h6b == io_state_in_1 ? 8'hc8 : _GEN_362; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_364 = 8'h6c == io_state_in_1 ? 8'hf9 : _GEN_363; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_365 = 8'h6d == io_state_in_1 ? 8'hf2 : _GEN_364; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_366 = 8'h6e == io_state_in_1 ? 8'hef : _GEN_365; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_367 = 8'h6f == io_state_in_1 ? 8'he4 : _GEN_366; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_368 = 8'h70 == io_state_in_1 ? 8'h3d : _GEN_367; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_369 = 8'h71 == io_state_in_1 ? 8'h36 : _GEN_368; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_370 = 8'h72 == io_state_in_1 ? 8'h2b : _GEN_369; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_371 = 8'h73 == io_state_in_1 ? 8'h20 : _GEN_370; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_372 = 8'h74 == io_state_in_1 ? 8'h11 : _GEN_371; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_373 = 8'h75 == io_state_in_1 ? 8'h1a : _GEN_372; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_374 = 8'h76 == io_state_in_1 ? 8'h7 : _GEN_373; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_375 = 8'h77 == io_state_in_1 ? 8'hc : _GEN_374; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_376 = 8'h78 == io_state_in_1 ? 8'h65 : _GEN_375; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_377 = 8'h79 == io_state_in_1 ? 8'h6e : _GEN_376; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_378 = 8'h7a == io_state_in_1 ? 8'h73 : _GEN_377; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_379 = 8'h7b == io_state_in_1 ? 8'h78 : _GEN_378; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_380 = 8'h7c == io_state_in_1 ? 8'h49 : _GEN_379; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_381 = 8'h7d == io_state_in_1 ? 8'h42 : _GEN_380; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_382 = 8'h7e == io_state_in_1 ? 8'h5f : _GEN_381; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_383 = 8'h7f == io_state_in_1 ? 8'h54 : _GEN_382; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_384 = 8'h80 == io_state_in_1 ? 8'hf7 : _GEN_383; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_385 = 8'h81 == io_state_in_1 ? 8'hfc : _GEN_384; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_386 = 8'h82 == io_state_in_1 ? 8'he1 : _GEN_385; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_387 = 8'h83 == io_state_in_1 ? 8'hea : _GEN_386; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_388 = 8'h84 == io_state_in_1 ? 8'hdb : _GEN_387; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_389 = 8'h85 == io_state_in_1 ? 8'hd0 : _GEN_388; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_390 = 8'h86 == io_state_in_1 ? 8'hcd : _GEN_389; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_391 = 8'h87 == io_state_in_1 ? 8'hc6 : _GEN_390; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_392 = 8'h88 == io_state_in_1 ? 8'haf : _GEN_391; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_393 = 8'h89 == io_state_in_1 ? 8'ha4 : _GEN_392; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_394 = 8'h8a == io_state_in_1 ? 8'hb9 : _GEN_393; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_395 = 8'h8b == io_state_in_1 ? 8'hb2 : _GEN_394; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_396 = 8'h8c == io_state_in_1 ? 8'h83 : _GEN_395; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_397 = 8'h8d == io_state_in_1 ? 8'h88 : _GEN_396; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_398 = 8'h8e == io_state_in_1 ? 8'h95 : _GEN_397; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_399 = 8'h8f == io_state_in_1 ? 8'h9e : _GEN_398; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_400 = 8'h90 == io_state_in_1 ? 8'h47 : _GEN_399; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_401 = 8'h91 == io_state_in_1 ? 8'h4c : _GEN_400; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_402 = 8'h92 == io_state_in_1 ? 8'h51 : _GEN_401; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_403 = 8'h93 == io_state_in_1 ? 8'h5a : _GEN_402; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_404 = 8'h94 == io_state_in_1 ? 8'h6b : _GEN_403; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_405 = 8'h95 == io_state_in_1 ? 8'h60 : _GEN_404; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_406 = 8'h96 == io_state_in_1 ? 8'h7d : _GEN_405; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_407 = 8'h97 == io_state_in_1 ? 8'h76 : _GEN_406; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_408 = 8'h98 == io_state_in_1 ? 8'h1f : _GEN_407; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_409 = 8'h99 == io_state_in_1 ? 8'h14 : _GEN_408; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_410 = 8'h9a == io_state_in_1 ? 8'h9 : _GEN_409; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_411 = 8'h9b == io_state_in_1 ? 8'h2 : _GEN_410; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_412 = 8'h9c == io_state_in_1 ? 8'h33 : _GEN_411; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_413 = 8'h9d == io_state_in_1 ? 8'h38 : _GEN_412; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_414 = 8'h9e == io_state_in_1 ? 8'h25 : _GEN_413; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_415 = 8'h9f == io_state_in_1 ? 8'h2e : _GEN_414; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_416 = 8'ha0 == io_state_in_1 ? 8'h8c : _GEN_415; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_417 = 8'ha1 == io_state_in_1 ? 8'h87 : _GEN_416; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_418 = 8'ha2 == io_state_in_1 ? 8'h9a : _GEN_417; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_419 = 8'ha3 == io_state_in_1 ? 8'h91 : _GEN_418; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_420 = 8'ha4 == io_state_in_1 ? 8'ha0 : _GEN_419; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_421 = 8'ha5 == io_state_in_1 ? 8'hab : _GEN_420; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_422 = 8'ha6 == io_state_in_1 ? 8'hb6 : _GEN_421; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_423 = 8'ha7 == io_state_in_1 ? 8'hbd : _GEN_422; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_424 = 8'ha8 == io_state_in_1 ? 8'hd4 : _GEN_423; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_425 = 8'ha9 == io_state_in_1 ? 8'hdf : _GEN_424; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_426 = 8'haa == io_state_in_1 ? 8'hc2 : _GEN_425; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_427 = 8'hab == io_state_in_1 ? 8'hc9 : _GEN_426; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_428 = 8'hac == io_state_in_1 ? 8'hf8 : _GEN_427; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_429 = 8'had == io_state_in_1 ? 8'hf3 : _GEN_428; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_430 = 8'hae == io_state_in_1 ? 8'hee : _GEN_429; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_431 = 8'haf == io_state_in_1 ? 8'he5 : _GEN_430; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_432 = 8'hb0 == io_state_in_1 ? 8'h3c : _GEN_431; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_433 = 8'hb1 == io_state_in_1 ? 8'h37 : _GEN_432; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_434 = 8'hb2 == io_state_in_1 ? 8'h2a : _GEN_433; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_435 = 8'hb3 == io_state_in_1 ? 8'h21 : _GEN_434; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_436 = 8'hb4 == io_state_in_1 ? 8'h10 : _GEN_435; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_437 = 8'hb5 == io_state_in_1 ? 8'h1b : _GEN_436; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_438 = 8'hb6 == io_state_in_1 ? 8'h6 : _GEN_437; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_439 = 8'hb7 == io_state_in_1 ? 8'hd : _GEN_438; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_440 = 8'hb8 == io_state_in_1 ? 8'h64 : _GEN_439; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_441 = 8'hb9 == io_state_in_1 ? 8'h6f : _GEN_440; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_442 = 8'hba == io_state_in_1 ? 8'h72 : _GEN_441; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_443 = 8'hbb == io_state_in_1 ? 8'h79 : _GEN_442; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_444 = 8'hbc == io_state_in_1 ? 8'h48 : _GEN_443; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_445 = 8'hbd == io_state_in_1 ? 8'h43 : _GEN_444; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_446 = 8'hbe == io_state_in_1 ? 8'h5e : _GEN_445; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_447 = 8'hbf == io_state_in_1 ? 8'h55 : _GEN_446; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_448 = 8'hc0 == io_state_in_1 ? 8'h1 : _GEN_447; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_449 = 8'hc1 == io_state_in_1 ? 8'ha : _GEN_448; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_450 = 8'hc2 == io_state_in_1 ? 8'h17 : _GEN_449; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_451 = 8'hc3 == io_state_in_1 ? 8'h1c : _GEN_450; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_452 = 8'hc4 == io_state_in_1 ? 8'h2d : _GEN_451; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_453 = 8'hc5 == io_state_in_1 ? 8'h26 : _GEN_452; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_454 = 8'hc6 == io_state_in_1 ? 8'h3b : _GEN_453; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_455 = 8'hc7 == io_state_in_1 ? 8'h30 : _GEN_454; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_456 = 8'hc8 == io_state_in_1 ? 8'h59 : _GEN_455; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_457 = 8'hc9 == io_state_in_1 ? 8'h52 : _GEN_456; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_458 = 8'hca == io_state_in_1 ? 8'h4f : _GEN_457; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_459 = 8'hcb == io_state_in_1 ? 8'h44 : _GEN_458; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_460 = 8'hcc == io_state_in_1 ? 8'h75 : _GEN_459; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_461 = 8'hcd == io_state_in_1 ? 8'h7e : _GEN_460; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_462 = 8'hce == io_state_in_1 ? 8'h63 : _GEN_461; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_463 = 8'hcf == io_state_in_1 ? 8'h68 : _GEN_462; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_464 = 8'hd0 == io_state_in_1 ? 8'hb1 : _GEN_463; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_465 = 8'hd1 == io_state_in_1 ? 8'hba : _GEN_464; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_466 = 8'hd2 == io_state_in_1 ? 8'ha7 : _GEN_465; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_467 = 8'hd3 == io_state_in_1 ? 8'hac : _GEN_466; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_468 = 8'hd4 == io_state_in_1 ? 8'h9d : _GEN_467; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_469 = 8'hd5 == io_state_in_1 ? 8'h96 : _GEN_468; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_470 = 8'hd6 == io_state_in_1 ? 8'h8b : _GEN_469; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_471 = 8'hd7 == io_state_in_1 ? 8'h80 : _GEN_470; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_472 = 8'hd8 == io_state_in_1 ? 8'he9 : _GEN_471; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_473 = 8'hd9 == io_state_in_1 ? 8'he2 : _GEN_472; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_474 = 8'hda == io_state_in_1 ? 8'hff : _GEN_473; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_475 = 8'hdb == io_state_in_1 ? 8'hf4 : _GEN_474; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_476 = 8'hdc == io_state_in_1 ? 8'hc5 : _GEN_475; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_477 = 8'hdd == io_state_in_1 ? 8'hce : _GEN_476; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_478 = 8'hde == io_state_in_1 ? 8'hd3 : _GEN_477; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_479 = 8'hdf == io_state_in_1 ? 8'hd8 : _GEN_478; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_480 = 8'he0 == io_state_in_1 ? 8'h7a : _GEN_479; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_481 = 8'he1 == io_state_in_1 ? 8'h71 : _GEN_480; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_482 = 8'he2 == io_state_in_1 ? 8'h6c : _GEN_481; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_483 = 8'he3 == io_state_in_1 ? 8'h67 : _GEN_482; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_484 = 8'he4 == io_state_in_1 ? 8'h56 : _GEN_483; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_485 = 8'he5 == io_state_in_1 ? 8'h5d : _GEN_484; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_486 = 8'he6 == io_state_in_1 ? 8'h40 : _GEN_485; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_487 = 8'he7 == io_state_in_1 ? 8'h4b : _GEN_486; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_488 = 8'he8 == io_state_in_1 ? 8'h22 : _GEN_487; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_489 = 8'he9 == io_state_in_1 ? 8'h29 : _GEN_488; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_490 = 8'hea == io_state_in_1 ? 8'h34 : _GEN_489; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_491 = 8'heb == io_state_in_1 ? 8'h3f : _GEN_490; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_492 = 8'hec == io_state_in_1 ? 8'he : _GEN_491; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_493 = 8'hed == io_state_in_1 ? 8'h5 : _GEN_492; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_494 = 8'hee == io_state_in_1 ? 8'h18 : _GEN_493; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_495 = 8'hef == io_state_in_1 ? 8'h13 : _GEN_494; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_496 = 8'hf0 == io_state_in_1 ? 8'hca : _GEN_495; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_497 = 8'hf1 == io_state_in_1 ? 8'hc1 : _GEN_496; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_498 = 8'hf2 == io_state_in_1 ? 8'hdc : _GEN_497; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_499 = 8'hf3 == io_state_in_1 ? 8'hd7 : _GEN_498; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_500 = 8'hf4 == io_state_in_1 ? 8'he6 : _GEN_499; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_501 = 8'hf5 == io_state_in_1 ? 8'hed : _GEN_500; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_502 = 8'hf6 == io_state_in_1 ? 8'hf0 : _GEN_501; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_503 = 8'hf7 == io_state_in_1 ? 8'hfb : _GEN_502; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_504 = 8'hf8 == io_state_in_1 ? 8'h92 : _GEN_503; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_505 = 8'hf9 == io_state_in_1 ? 8'h99 : _GEN_504; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_506 = 8'hfa == io_state_in_1 ? 8'h84 : _GEN_505; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_507 = 8'hfb == io_state_in_1 ? 8'h8f : _GEN_506; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_508 = 8'hfc == io_state_in_1 ? 8'hbe : _GEN_507; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_509 = 8'hfd == io_state_in_1 ? 8'hb5 : _GEN_508; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_510 = 8'hfe == io_state_in_1 ? 8'ha8 : _GEN_509; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _GEN_511 = 8'hff == io_state_in_1 ? 8'ha3 : _GEN_510; // @[InvMixColumns.scala 126:{41,41}]
  wire [7:0] _tmp_state_0_T = _GEN_255 ^ _GEN_511; // @[InvMixColumns.scala 126:41]
  wire [7:0] _GEN_513 = 8'h1 == io_state_in_2 ? 8'hd : 8'h0; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_514 = 8'h2 == io_state_in_2 ? 8'h1a : _GEN_513; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_515 = 8'h3 == io_state_in_2 ? 8'h17 : _GEN_514; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_516 = 8'h4 == io_state_in_2 ? 8'h34 : _GEN_515; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_517 = 8'h5 == io_state_in_2 ? 8'h39 : _GEN_516; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_518 = 8'h6 == io_state_in_2 ? 8'h2e : _GEN_517; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_519 = 8'h7 == io_state_in_2 ? 8'h23 : _GEN_518; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_520 = 8'h8 == io_state_in_2 ? 8'h68 : _GEN_519; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_521 = 8'h9 == io_state_in_2 ? 8'h65 : _GEN_520; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_522 = 8'ha == io_state_in_2 ? 8'h72 : _GEN_521; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_523 = 8'hb == io_state_in_2 ? 8'h7f : _GEN_522; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_524 = 8'hc == io_state_in_2 ? 8'h5c : _GEN_523; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_525 = 8'hd == io_state_in_2 ? 8'h51 : _GEN_524; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_526 = 8'he == io_state_in_2 ? 8'h46 : _GEN_525; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_527 = 8'hf == io_state_in_2 ? 8'h4b : _GEN_526; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_528 = 8'h10 == io_state_in_2 ? 8'hd0 : _GEN_527; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_529 = 8'h11 == io_state_in_2 ? 8'hdd : _GEN_528; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_530 = 8'h12 == io_state_in_2 ? 8'hca : _GEN_529; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_531 = 8'h13 == io_state_in_2 ? 8'hc7 : _GEN_530; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_532 = 8'h14 == io_state_in_2 ? 8'he4 : _GEN_531; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_533 = 8'h15 == io_state_in_2 ? 8'he9 : _GEN_532; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_534 = 8'h16 == io_state_in_2 ? 8'hfe : _GEN_533; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_535 = 8'h17 == io_state_in_2 ? 8'hf3 : _GEN_534; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_536 = 8'h18 == io_state_in_2 ? 8'hb8 : _GEN_535; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_537 = 8'h19 == io_state_in_2 ? 8'hb5 : _GEN_536; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_538 = 8'h1a == io_state_in_2 ? 8'ha2 : _GEN_537; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_539 = 8'h1b == io_state_in_2 ? 8'haf : _GEN_538; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_540 = 8'h1c == io_state_in_2 ? 8'h8c : _GEN_539; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_541 = 8'h1d == io_state_in_2 ? 8'h81 : _GEN_540; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_542 = 8'h1e == io_state_in_2 ? 8'h96 : _GEN_541; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_543 = 8'h1f == io_state_in_2 ? 8'h9b : _GEN_542; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_544 = 8'h20 == io_state_in_2 ? 8'hbb : _GEN_543; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_545 = 8'h21 == io_state_in_2 ? 8'hb6 : _GEN_544; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_546 = 8'h22 == io_state_in_2 ? 8'ha1 : _GEN_545; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_547 = 8'h23 == io_state_in_2 ? 8'hac : _GEN_546; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_548 = 8'h24 == io_state_in_2 ? 8'h8f : _GEN_547; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_549 = 8'h25 == io_state_in_2 ? 8'h82 : _GEN_548; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_550 = 8'h26 == io_state_in_2 ? 8'h95 : _GEN_549; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_551 = 8'h27 == io_state_in_2 ? 8'h98 : _GEN_550; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_552 = 8'h28 == io_state_in_2 ? 8'hd3 : _GEN_551; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_553 = 8'h29 == io_state_in_2 ? 8'hde : _GEN_552; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_554 = 8'h2a == io_state_in_2 ? 8'hc9 : _GEN_553; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_555 = 8'h2b == io_state_in_2 ? 8'hc4 : _GEN_554; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_556 = 8'h2c == io_state_in_2 ? 8'he7 : _GEN_555; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_557 = 8'h2d == io_state_in_2 ? 8'hea : _GEN_556; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_558 = 8'h2e == io_state_in_2 ? 8'hfd : _GEN_557; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_559 = 8'h2f == io_state_in_2 ? 8'hf0 : _GEN_558; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_560 = 8'h30 == io_state_in_2 ? 8'h6b : _GEN_559; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_561 = 8'h31 == io_state_in_2 ? 8'h66 : _GEN_560; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_562 = 8'h32 == io_state_in_2 ? 8'h71 : _GEN_561; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_563 = 8'h33 == io_state_in_2 ? 8'h7c : _GEN_562; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_564 = 8'h34 == io_state_in_2 ? 8'h5f : _GEN_563; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_565 = 8'h35 == io_state_in_2 ? 8'h52 : _GEN_564; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_566 = 8'h36 == io_state_in_2 ? 8'h45 : _GEN_565; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_567 = 8'h37 == io_state_in_2 ? 8'h48 : _GEN_566; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_568 = 8'h38 == io_state_in_2 ? 8'h3 : _GEN_567; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_569 = 8'h39 == io_state_in_2 ? 8'he : _GEN_568; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_570 = 8'h3a == io_state_in_2 ? 8'h19 : _GEN_569; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_571 = 8'h3b == io_state_in_2 ? 8'h14 : _GEN_570; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_572 = 8'h3c == io_state_in_2 ? 8'h37 : _GEN_571; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_573 = 8'h3d == io_state_in_2 ? 8'h3a : _GEN_572; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_574 = 8'h3e == io_state_in_2 ? 8'h2d : _GEN_573; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_575 = 8'h3f == io_state_in_2 ? 8'h20 : _GEN_574; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_576 = 8'h40 == io_state_in_2 ? 8'h6d : _GEN_575; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_577 = 8'h41 == io_state_in_2 ? 8'h60 : _GEN_576; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_578 = 8'h42 == io_state_in_2 ? 8'h77 : _GEN_577; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_579 = 8'h43 == io_state_in_2 ? 8'h7a : _GEN_578; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_580 = 8'h44 == io_state_in_2 ? 8'h59 : _GEN_579; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_581 = 8'h45 == io_state_in_2 ? 8'h54 : _GEN_580; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_582 = 8'h46 == io_state_in_2 ? 8'h43 : _GEN_581; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_583 = 8'h47 == io_state_in_2 ? 8'h4e : _GEN_582; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_584 = 8'h48 == io_state_in_2 ? 8'h5 : _GEN_583; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_585 = 8'h49 == io_state_in_2 ? 8'h8 : _GEN_584; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_586 = 8'h4a == io_state_in_2 ? 8'h1f : _GEN_585; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_587 = 8'h4b == io_state_in_2 ? 8'h12 : _GEN_586; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_588 = 8'h4c == io_state_in_2 ? 8'h31 : _GEN_587; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_589 = 8'h4d == io_state_in_2 ? 8'h3c : _GEN_588; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_590 = 8'h4e == io_state_in_2 ? 8'h2b : _GEN_589; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_591 = 8'h4f == io_state_in_2 ? 8'h26 : _GEN_590; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_592 = 8'h50 == io_state_in_2 ? 8'hbd : _GEN_591; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_593 = 8'h51 == io_state_in_2 ? 8'hb0 : _GEN_592; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_594 = 8'h52 == io_state_in_2 ? 8'ha7 : _GEN_593; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_595 = 8'h53 == io_state_in_2 ? 8'haa : _GEN_594; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_596 = 8'h54 == io_state_in_2 ? 8'h89 : _GEN_595; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_597 = 8'h55 == io_state_in_2 ? 8'h84 : _GEN_596; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_598 = 8'h56 == io_state_in_2 ? 8'h93 : _GEN_597; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_599 = 8'h57 == io_state_in_2 ? 8'h9e : _GEN_598; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_600 = 8'h58 == io_state_in_2 ? 8'hd5 : _GEN_599; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_601 = 8'h59 == io_state_in_2 ? 8'hd8 : _GEN_600; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_602 = 8'h5a == io_state_in_2 ? 8'hcf : _GEN_601; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_603 = 8'h5b == io_state_in_2 ? 8'hc2 : _GEN_602; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_604 = 8'h5c == io_state_in_2 ? 8'he1 : _GEN_603; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_605 = 8'h5d == io_state_in_2 ? 8'hec : _GEN_604; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_606 = 8'h5e == io_state_in_2 ? 8'hfb : _GEN_605; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_607 = 8'h5f == io_state_in_2 ? 8'hf6 : _GEN_606; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_608 = 8'h60 == io_state_in_2 ? 8'hd6 : _GEN_607; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_609 = 8'h61 == io_state_in_2 ? 8'hdb : _GEN_608; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_610 = 8'h62 == io_state_in_2 ? 8'hcc : _GEN_609; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_611 = 8'h63 == io_state_in_2 ? 8'hc1 : _GEN_610; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_612 = 8'h64 == io_state_in_2 ? 8'he2 : _GEN_611; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_613 = 8'h65 == io_state_in_2 ? 8'hef : _GEN_612; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_614 = 8'h66 == io_state_in_2 ? 8'hf8 : _GEN_613; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_615 = 8'h67 == io_state_in_2 ? 8'hf5 : _GEN_614; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_616 = 8'h68 == io_state_in_2 ? 8'hbe : _GEN_615; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_617 = 8'h69 == io_state_in_2 ? 8'hb3 : _GEN_616; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_618 = 8'h6a == io_state_in_2 ? 8'ha4 : _GEN_617; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_619 = 8'h6b == io_state_in_2 ? 8'ha9 : _GEN_618; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_620 = 8'h6c == io_state_in_2 ? 8'h8a : _GEN_619; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_621 = 8'h6d == io_state_in_2 ? 8'h87 : _GEN_620; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_622 = 8'h6e == io_state_in_2 ? 8'h90 : _GEN_621; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_623 = 8'h6f == io_state_in_2 ? 8'h9d : _GEN_622; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_624 = 8'h70 == io_state_in_2 ? 8'h6 : _GEN_623; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_625 = 8'h71 == io_state_in_2 ? 8'hb : _GEN_624; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_626 = 8'h72 == io_state_in_2 ? 8'h1c : _GEN_625; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_627 = 8'h73 == io_state_in_2 ? 8'h11 : _GEN_626; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_628 = 8'h74 == io_state_in_2 ? 8'h32 : _GEN_627; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_629 = 8'h75 == io_state_in_2 ? 8'h3f : _GEN_628; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_630 = 8'h76 == io_state_in_2 ? 8'h28 : _GEN_629; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_631 = 8'h77 == io_state_in_2 ? 8'h25 : _GEN_630; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_632 = 8'h78 == io_state_in_2 ? 8'h6e : _GEN_631; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_633 = 8'h79 == io_state_in_2 ? 8'h63 : _GEN_632; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_634 = 8'h7a == io_state_in_2 ? 8'h74 : _GEN_633; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_635 = 8'h7b == io_state_in_2 ? 8'h79 : _GEN_634; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_636 = 8'h7c == io_state_in_2 ? 8'h5a : _GEN_635; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_637 = 8'h7d == io_state_in_2 ? 8'h57 : _GEN_636; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_638 = 8'h7e == io_state_in_2 ? 8'h40 : _GEN_637; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_639 = 8'h7f == io_state_in_2 ? 8'h4d : _GEN_638; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_640 = 8'h80 == io_state_in_2 ? 8'hda : _GEN_639; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_641 = 8'h81 == io_state_in_2 ? 8'hd7 : _GEN_640; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_642 = 8'h82 == io_state_in_2 ? 8'hc0 : _GEN_641; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_643 = 8'h83 == io_state_in_2 ? 8'hcd : _GEN_642; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_644 = 8'h84 == io_state_in_2 ? 8'hee : _GEN_643; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_645 = 8'h85 == io_state_in_2 ? 8'he3 : _GEN_644; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_646 = 8'h86 == io_state_in_2 ? 8'hf4 : _GEN_645; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_647 = 8'h87 == io_state_in_2 ? 8'hf9 : _GEN_646; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_648 = 8'h88 == io_state_in_2 ? 8'hb2 : _GEN_647; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_649 = 8'h89 == io_state_in_2 ? 8'hbf : _GEN_648; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_650 = 8'h8a == io_state_in_2 ? 8'ha8 : _GEN_649; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_651 = 8'h8b == io_state_in_2 ? 8'ha5 : _GEN_650; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_652 = 8'h8c == io_state_in_2 ? 8'h86 : _GEN_651; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_653 = 8'h8d == io_state_in_2 ? 8'h8b : _GEN_652; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_654 = 8'h8e == io_state_in_2 ? 8'h9c : _GEN_653; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_655 = 8'h8f == io_state_in_2 ? 8'h91 : _GEN_654; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_656 = 8'h90 == io_state_in_2 ? 8'ha : _GEN_655; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_657 = 8'h91 == io_state_in_2 ? 8'h7 : _GEN_656; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_658 = 8'h92 == io_state_in_2 ? 8'h10 : _GEN_657; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_659 = 8'h93 == io_state_in_2 ? 8'h1d : _GEN_658; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_660 = 8'h94 == io_state_in_2 ? 8'h3e : _GEN_659; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_661 = 8'h95 == io_state_in_2 ? 8'h33 : _GEN_660; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_662 = 8'h96 == io_state_in_2 ? 8'h24 : _GEN_661; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_663 = 8'h97 == io_state_in_2 ? 8'h29 : _GEN_662; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_664 = 8'h98 == io_state_in_2 ? 8'h62 : _GEN_663; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_665 = 8'h99 == io_state_in_2 ? 8'h6f : _GEN_664; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_666 = 8'h9a == io_state_in_2 ? 8'h78 : _GEN_665; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_667 = 8'h9b == io_state_in_2 ? 8'h75 : _GEN_666; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_668 = 8'h9c == io_state_in_2 ? 8'h56 : _GEN_667; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_669 = 8'h9d == io_state_in_2 ? 8'h5b : _GEN_668; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_670 = 8'h9e == io_state_in_2 ? 8'h4c : _GEN_669; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_671 = 8'h9f == io_state_in_2 ? 8'h41 : _GEN_670; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_672 = 8'ha0 == io_state_in_2 ? 8'h61 : _GEN_671; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_673 = 8'ha1 == io_state_in_2 ? 8'h6c : _GEN_672; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_674 = 8'ha2 == io_state_in_2 ? 8'h7b : _GEN_673; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_675 = 8'ha3 == io_state_in_2 ? 8'h76 : _GEN_674; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_676 = 8'ha4 == io_state_in_2 ? 8'h55 : _GEN_675; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_677 = 8'ha5 == io_state_in_2 ? 8'h58 : _GEN_676; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_678 = 8'ha6 == io_state_in_2 ? 8'h4f : _GEN_677; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_679 = 8'ha7 == io_state_in_2 ? 8'h42 : _GEN_678; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_680 = 8'ha8 == io_state_in_2 ? 8'h9 : _GEN_679; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_681 = 8'ha9 == io_state_in_2 ? 8'h4 : _GEN_680; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_682 = 8'haa == io_state_in_2 ? 8'h13 : _GEN_681; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_683 = 8'hab == io_state_in_2 ? 8'h1e : _GEN_682; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_684 = 8'hac == io_state_in_2 ? 8'h3d : _GEN_683; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_685 = 8'had == io_state_in_2 ? 8'h30 : _GEN_684; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_686 = 8'hae == io_state_in_2 ? 8'h27 : _GEN_685; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_687 = 8'haf == io_state_in_2 ? 8'h2a : _GEN_686; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_688 = 8'hb0 == io_state_in_2 ? 8'hb1 : _GEN_687; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_689 = 8'hb1 == io_state_in_2 ? 8'hbc : _GEN_688; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_690 = 8'hb2 == io_state_in_2 ? 8'hab : _GEN_689; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_691 = 8'hb3 == io_state_in_2 ? 8'ha6 : _GEN_690; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_692 = 8'hb4 == io_state_in_2 ? 8'h85 : _GEN_691; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_693 = 8'hb5 == io_state_in_2 ? 8'h88 : _GEN_692; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_694 = 8'hb6 == io_state_in_2 ? 8'h9f : _GEN_693; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_695 = 8'hb7 == io_state_in_2 ? 8'h92 : _GEN_694; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_696 = 8'hb8 == io_state_in_2 ? 8'hd9 : _GEN_695; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_697 = 8'hb9 == io_state_in_2 ? 8'hd4 : _GEN_696; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_698 = 8'hba == io_state_in_2 ? 8'hc3 : _GEN_697; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_699 = 8'hbb == io_state_in_2 ? 8'hce : _GEN_698; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_700 = 8'hbc == io_state_in_2 ? 8'hed : _GEN_699; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_701 = 8'hbd == io_state_in_2 ? 8'he0 : _GEN_700; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_702 = 8'hbe == io_state_in_2 ? 8'hf7 : _GEN_701; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_703 = 8'hbf == io_state_in_2 ? 8'hfa : _GEN_702; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_704 = 8'hc0 == io_state_in_2 ? 8'hb7 : _GEN_703; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_705 = 8'hc1 == io_state_in_2 ? 8'hba : _GEN_704; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_706 = 8'hc2 == io_state_in_2 ? 8'had : _GEN_705; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_707 = 8'hc3 == io_state_in_2 ? 8'ha0 : _GEN_706; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_708 = 8'hc4 == io_state_in_2 ? 8'h83 : _GEN_707; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_709 = 8'hc5 == io_state_in_2 ? 8'h8e : _GEN_708; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_710 = 8'hc6 == io_state_in_2 ? 8'h99 : _GEN_709; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_711 = 8'hc7 == io_state_in_2 ? 8'h94 : _GEN_710; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_712 = 8'hc8 == io_state_in_2 ? 8'hdf : _GEN_711; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_713 = 8'hc9 == io_state_in_2 ? 8'hd2 : _GEN_712; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_714 = 8'hca == io_state_in_2 ? 8'hc5 : _GEN_713; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_715 = 8'hcb == io_state_in_2 ? 8'hc8 : _GEN_714; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_716 = 8'hcc == io_state_in_2 ? 8'heb : _GEN_715; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_717 = 8'hcd == io_state_in_2 ? 8'he6 : _GEN_716; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_718 = 8'hce == io_state_in_2 ? 8'hf1 : _GEN_717; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_719 = 8'hcf == io_state_in_2 ? 8'hfc : _GEN_718; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_720 = 8'hd0 == io_state_in_2 ? 8'h67 : _GEN_719; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_721 = 8'hd1 == io_state_in_2 ? 8'h6a : _GEN_720; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_722 = 8'hd2 == io_state_in_2 ? 8'h7d : _GEN_721; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_723 = 8'hd3 == io_state_in_2 ? 8'h70 : _GEN_722; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_724 = 8'hd4 == io_state_in_2 ? 8'h53 : _GEN_723; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_725 = 8'hd5 == io_state_in_2 ? 8'h5e : _GEN_724; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_726 = 8'hd6 == io_state_in_2 ? 8'h49 : _GEN_725; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_727 = 8'hd7 == io_state_in_2 ? 8'h44 : _GEN_726; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_728 = 8'hd8 == io_state_in_2 ? 8'hf : _GEN_727; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_729 = 8'hd9 == io_state_in_2 ? 8'h2 : _GEN_728; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_730 = 8'hda == io_state_in_2 ? 8'h15 : _GEN_729; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_731 = 8'hdb == io_state_in_2 ? 8'h18 : _GEN_730; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_732 = 8'hdc == io_state_in_2 ? 8'h3b : _GEN_731; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_733 = 8'hdd == io_state_in_2 ? 8'h36 : _GEN_732; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_734 = 8'hde == io_state_in_2 ? 8'h21 : _GEN_733; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_735 = 8'hdf == io_state_in_2 ? 8'h2c : _GEN_734; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_736 = 8'he0 == io_state_in_2 ? 8'hc : _GEN_735; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_737 = 8'he1 == io_state_in_2 ? 8'h1 : _GEN_736; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_738 = 8'he2 == io_state_in_2 ? 8'h16 : _GEN_737; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_739 = 8'he3 == io_state_in_2 ? 8'h1b : _GEN_738; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_740 = 8'he4 == io_state_in_2 ? 8'h38 : _GEN_739; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_741 = 8'he5 == io_state_in_2 ? 8'h35 : _GEN_740; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_742 = 8'he6 == io_state_in_2 ? 8'h22 : _GEN_741; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_743 = 8'he7 == io_state_in_2 ? 8'h2f : _GEN_742; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_744 = 8'he8 == io_state_in_2 ? 8'h64 : _GEN_743; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_745 = 8'he9 == io_state_in_2 ? 8'h69 : _GEN_744; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_746 = 8'hea == io_state_in_2 ? 8'h7e : _GEN_745; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_747 = 8'heb == io_state_in_2 ? 8'h73 : _GEN_746; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_748 = 8'hec == io_state_in_2 ? 8'h50 : _GEN_747; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_749 = 8'hed == io_state_in_2 ? 8'h5d : _GEN_748; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_750 = 8'hee == io_state_in_2 ? 8'h4a : _GEN_749; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_751 = 8'hef == io_state_in_2 ? 8'h47 : _GEN_750; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_752 = 8'hf0 == io_state_in_2 ? 8'hdc : _GEN_751; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_753 = 8'hf1 == io_state_in_2 ? 8'hd1 : _GEN_752; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_754 = 8'hf2 == io_state_in_2 ? 8'hc6 : _GEN_753; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_755 = 8'hf3 == io_state_in_2 ? 8'hcb : _GEN_754; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_756 = 8'hf4 == io_state_in_2 ? 8'he8 : _GEN_755; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_757 = 8'hf5 == io_state_in_2 ? 8'he5 : _GEN_756; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_758 = 8'hf6 == io_state_in_2 ? 8'hf2 : _GEN_757; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_759 = 8'hf7 == io_state_in_2 ? 8'hff : _GEN_758; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_760 = 8'hf8 == io_state_in_2 ? 8'hb4 : _GEN_759; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_761 = 8'hf9 == io_state_in_2 ? 8'hb9 : _GEN_760; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_762 = 8'hfa == io_state_in_2 ? 8'hae : _GEN_761; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_763 = 8'hfb == io_state_in_2 ? 8'ha3 : _GEN_762; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_764 = 8'hfc == io_state_in_2 ? 8'h80 : _GEN_763; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_765 = 8'hfd == io_state_in_2 ? 8'h8d : _GEN_764; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_766 = 8'hfe == io_state_in_2 ? 8'h9a : _GEN_765; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _GEN_767 = 8'hff == io_state_in_2 ? 8'h97 : _GEN_766; // @[InvMixColumns.scala 126:{65,65}]
  wire [7:0] _tmp_state_0_T_1 = _tmp_state_0_T ^ _GEN_767; // @[InvMixColumns.scala 126:65]
  wire [7:0] _GEN_769 = 8'h1 == io_state_in_3 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_770 = 8'h2 == io_state_in_3 ? 8'h12 : _GEN_769; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_771 = 8'h3 == io_state_in_3 ? 8'h1b : _GEN_770; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_772 = 8'h4 == io_state_in_3 ? 8'h24 : _GEN_771; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_773 = 8'h5 == io_state_in_3 ? 8'h2d : _GEN_772; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_774 = 8'h6 == io_state_in_3 ? 8'h36 : _GEN_773; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_775 = 8'h7 == io_state_in_3 ? 8'h3f : _GEN_774; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_776 = 8'h8 == io_state_in_3 ? 8'h48 : _GEN_775; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_777 = 8'h9 == io_state_in_3 ? 8'h41 : _GEN_776; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_778 = 8'ha == io_state_in_3 ? 8'h5a : _GEN_777; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_779 = 8'hb == io_state_in_3 ? 8'h53 : _GEN_778; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_780 = 8'hc == io_state_in_3 ? 8'h6c : _GEN_779; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_781 = 8'hd == io_state_in_3 ? 8'h65 : _GEN_780; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_782 = 8'he == io_state_in_3 ? 8'h7e : _GEN_781; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_783 = 8'hf == io_state_in_3 ? 8'h77 : _GEN_782; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_784 = 8'h10 == io_state_in_3 ? 8'h90 : _GEN_783; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_785 = 8'h11 == io_state_in_3 ? 8'h99 : _GEN_784; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_786 = 8'h12 == io_state_in_3 ? 8'h82 : _GEN_785; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_787 = 8'h13 == io_state_in_3 ? 8'h8b : _GEN_786; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_788 = 8'h14 == io_state_in_3 ? 8'hb4 : _GEN_787; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_789 = 8'h15 == io_state_in_3 ? 8'hbd : _GEN_788; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_790 = 8'h16 == io_state_in_3 ? 8'ha6 : _GEN_789; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_791 = 8'h17 == io_state_in_3 ? 8'haf : _GEN_790; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_792 = 8'h18 == io_state_in_3 ? 8'hd8 : _GEN_791; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_793 = 8'h19 == io_state_in_3 ? 8'hd1 : _GEN_792; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_794 = 8'h1a == io_state_in_3 ? 8'hca : _GEN_793; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_795 = 8'h1b == io_state_in_3 ? 8'hc3 : _GEN_794; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_796 = 8'h1c == io_state_in_3 ? 8'hfc : _GEN_795; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_797 = 8'h1d == io_state_in_3 ? 8'hf5 : _GEN_796; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_798 = 8'h1e == io_state_in_3 ? 8'hee : _GEN_797; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_799 = 8'h1f == io_state_in_3 ? 8'he7 : _GEN_798; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_800 = 8'h20 == io_state_in_3 ? 8'h3b : _GEN_799; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_801 = 8'h21 == io_state_in_3 ? 8'h32 : _GEN_800; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_802 = 8'h22 == io_state_in_3 ? 8'h29 : _GEN_801; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_803 = 8'h23 == io_state_in_3 ? 8'h20 : _GEN_802; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_804 = 8'h24 == io_state_in_3 ? 8'h1f : _GEN_803; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_805 = 8'h25 == io_state_in_3 ? 8'h16 : _GEN_804; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_806 = 8'h26 == io_state_in_3 ? 8'hd : _GEN_805; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_807 = 8'h27 == io_state_in_3 ? 8'h4 : _GEN_806; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_808 = 8'h28 == io_state_in_3 ? 8'h73 : _GEN_807; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_809 = 8'h29 == io_state_in_3 ? 8'h7a : _GEN_808; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_810 = 8'h2a == io_state_in_3 ? 8'h61 : _GEN_809; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_811 = 8'h2b == io_state_in_3 ? 8'h68 : _GEN_810; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_812 = 8'h2c == io_state_in_3 ? 8'h57 : _GEN_811; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_813 = 8'h2d == io_state_in_3 ? 8'h5e : _GEN_812; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_814 = 8'h2e == io_state_in_3 ? 8'h45 : _GEN_813; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_815 = 8'h2f == io_state_in_3 ? 8'h4c : _GEN_814; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_816 = 8'h30 == io_state_in_3 ? 8'hab : _GEN_815; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_817 = 8'h31 == io_state_in_3 ? 8'ha2 : _GEN_816; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_818 = 8'h32 == io_state_in_3 ? 8'hb9 : _GEN_817; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_819 = 8'h33 == io_state_in_3 ? 8'hb0 : _GEN_818; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_820 = 8'h34 == io_state_in_3 ? 8'h8f : _GEN_819; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_821 = 8'h35 == io_state_in_3 ? 8'h86 : _GEN_820; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_822 = 8'h36 == io_state_in_3 ? 8'h9d : _GEN_821; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_823 = 8'h37 == io_state_in_3 ? 8'h94 : _GEN_822; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_824 = 8'h38 == io_state_in_3 ? 8'he3 : _GEN_823; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_825 = 8'h39 == io_state_in_3 ? 8'hea : _GEN_824; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_826 = 8'h3a == io_state_in_3 ? 8'hf1 : _GEN_825; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_827 = 8'h3b == io_state_in_3 ? 8'hf8 : _GEN_826; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_828 = 8'h3c == io_state_in_3 ? 8'hc7 : _GEN_827; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_829 = 8'h3d == io_state_in_3 ? 8'hce : _GEN_828; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_830 = 8'h3e == io_state_in_3 ? 8'hd5 : _GEN_829; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_831 = 8'h3f == io_state_in_3 ? 8'hdc : _GEN_830; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_832 = 8'h40 == io_state_in_3 ? 8'h76 : _GEN_831; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_833 = 8'h41 == io_state_in_3 ? 8'h7f : _GEN_832; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_834 = 8'h42 == io_state_in_3 ? 8'h64 : _GEN_833; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_835 = 8'h43 == io_state_in_3 ? 8'h6d : _GEN_834; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_836 = 8'h44 == io_state_in_3 ? 8'h52 : _GEN_835; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_837 = 8'h45 == io_state_in_3 ? 8'h5b : _GEN_836; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_838 = 8'h46 == io_state_in_3 ? 8'h40 : _GEN_837; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_839 = 8'h47 == io_state_in_3 ? 8'h49 : _GEN_838; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_840 = 8'h48 == io_state_in_3 ? 8'h3e : _GEN_839; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_841 = 8'h49 == io_state_in_3 ? 8'h37 : _GEN_840; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_842 = 8'h4a == io_state_in_3 ? 8'h2c : _GEN_841; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_843 = 8'h4b == io_state_in_3 ? 8'h25 : _GEN_842; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_844 = 8'h4c == io_state_in_3 ? 8'h1a : _GEN_843; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_845 = 8'h4d == io_state_in_3 ? 8'h13 : _GEN_844; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_846 = 8'h4e == io_state_in_3 ? 8'h8 : _GEN_845; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_847 = 8'h4f == io_state_in_3 ? 8'h1 : _GEN_846; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_848 = 8'h50 == io_state_in_3 ? 8'he6 : _GEN_847; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_849 = 8'h51 == io_state_in_3 ? 8'hef : _GEN_848; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_850 = 8'h52 == io_state_in_3 ? 8'hf4 : _GEN_849; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_851 = 8'h53 == io_state_in_3 ? 8'hfd : _GEN_850; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_852 = 8'h54 == io_state_in_3 ? 8'hc2 : _GEN_851; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_853 = 8'h55 == io_state_in_3 ? 8'hcb : _GEN_852; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_854 = 8'h56 == io_state_in_3 ? 8'hd0 : _GEN_853; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_855 = 8'h57 == io_state_in_3 ? 8'hd9 : _GEN_854; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_856 = 8'h58 == io_state_in_3 ? 8'hae : _GEN_855; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_857 = 8'h59 == io_state_in_3 ? 8'ha7 : _GEN_856; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_858 = 8'h5a == io_state_in_3 ? 8'hbc : _GEN_857; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_859 = 8'h5b == io_state_in_3 ? 8'hb5 : _GEN_858; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_860 = 8'h5c == io_state_in_3 ? 8'h8a : _GEN_859; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_861 = 8'h5d == io_state_in_3 ? 8'h83 : _GEN_860; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_862 = 8'h5e == io_state_in_3 ? 8'h98 : _GEN_861; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_863 = 8'h5f == io_state_in_3 ? 8'h91 : _GEN_862; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_864 = 8'h60 == io_state_in_3 ? 8'h4d : _GEN_863; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_865 = 8'h61 == io_state_in_3 ? 8'h44 : _GEN_864; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_866 = 8'h62 == io_state_in_3 ? 8'h5f : _GEN_865; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_867 = 8'h63 == io_state_in_3 ? 8'h56 : _GEN_866; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_868 = 8'h64 == io_state_in_3 ? 8'h69 : _GEN_867; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_869 = 8'h65 == io_state_in_3 ? 8'h60 : _GEN_868; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_870 = 8'h66 == io_state_in_3 ? 8'h7b : _GEN_869; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_871 = 8'h67 == io_state_in_3 ? 8'h72 : _GEN_870; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_872 = 8'h68 == io_state_in_3 ? 8'h5 : _GEN_871; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_873 = 8'h69 == io_state_in_3 ? 8'hc : _GEN_872; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_874 = 8'h6a == io_state_in_3 ? 8'h17 : _GEN_873; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_875 = 8'h6b == io_state_in_3 ? 8'h1e : _GEN_874; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_876 = 8'h6c == io_state_in_3 ? 8'h21 : _GEN_875; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_877 = 8'h6d == io_state_in_3 ? 8'h28 : _GEN_876; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_878 = 8'h6e == io_state_in_3 ? 8'h33 : _GEN_877; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_879 = 8'h6f == io_state_in_3 ? 8'h3a : _GEN_878; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_880 = 8'h70 == io_state_in_3 ? 8'hdd : _GEN_879; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_881 = 8'h71 == io_state_in_3 ? 8'hd4 : _GEN_880; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_882 = 8'h72 == io_state_in_3 ? 8'hcf : _GEN_881; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_883 = 8'h73 == io_state_in_3 ? 8'hc6 : _GEN_882; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_884 = 8'h74 == io_state_in_3 ? 8'hf9 : _GEN_883; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_885 = 8'h75 == io_state_in_3 ? 8'hf0 : _GEN_884; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_886 = 8'h76 == io_state_in_3 ? 8'heb : _GEN_885; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_887 = 8'h77 == io_state_in_3 ? 8'he2 : _GEN_886; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_888 = 8'h78 == io_state_in_3 ? 8'h95 : _GEN_887; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_889 = 8'h79 == io_state_in_3 ? 8'h9c : _GEN_888; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_890 = 8'h7a == io_state_in_3 ? 8'h87 : _GEN_889; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_891 = 8'h7b == io_state_in_3 ? 8'h8e : _GEN_890; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_892 = 8'h7c == io_state_in_3 ? 8'hb1 : _GEN_891; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_893 = 8'h7d == io_state_in_3 ? 8'hb8 : _GEN_892; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_894 = 8'h7e == io_state_in_3 ? 8'ha3 : _GEN_893; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_895 = 8'h7f == io_state_in_3 ? 8'haa : _GEN_894; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_896 = 8'h80 == io_state_in_3 ? 8'hec : _GEN_895; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_897 = 8'h81 == io_state_in_3 ? 8'he5 : _GEN_896; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_898 = 8'h82 == io_state_in_3 ? 8'hfe : _GEN_897; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_899 = 8'h83 == io_state_in_3 ? 8'hf7 : _GEN_898; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_900 = 8'h84 == io_state_in_3 ? 8'hc8 : _GEN_899; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_901 = 8'h85 == io_state_in_3 ? 8'hc1 : _GEN_900; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_902 = 8'h86 == io_state_in_3 ? 8'hda : _GEN_901; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_903 = 8'h87 == io_state_in_3 ? 8'hd3 : _GEN_902; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_904 = 8'h88 == io_state_in_3 ? 8'ha4 : _GEN_903; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_905 = 8'h89 == io_state_in_3 ? 8'had : _GEN_904; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_906 = 8'h8a == io_state_in_3 ? 8'hb6 : _GEN_905; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_907 = 8'h8b == io_state_in_3 ? 8'hbf : _GEN_906; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_908 = 8'h8c == io_state_in_3 ? 8'h80 : _GEN_907; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_909 = 8'h8d == io_state_in_3 ? 8'h89 : _GEN_908; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_910 = 8'h8e == io_state_in_3 ? 8'h92 : _GEN_909; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_911 = 8'h8f == io_state_in_3 ? 8'h9b : _GEN_910; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_912 = 8'h90 == io_state_in_3 ? 8'h7c : _GEN_911; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_913 = 8'h91 == io_state_in_3 ? 8'h75 : _GEN_912; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_914 = 8'h92 == io_state_in_3 ? 8'h6e : _GEN_913; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_915 = 8'h93 == io_state_in_3 ? 8'h67 : _GEN_914; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_916 = 8'h94 == io_state_in_3 ? 8'h58 : _GEN_915; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_917 = 8'h95 == io_state_in_3 ? 8'h51 : _GEN_916; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_918 = 8'h96 == io_state_in_3 ? 8'h4a : _GEN_917; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_919 = 8'h97 == io_state_in_3 ? 8'h43 : _GEN_918; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_920 = 8'h98 == io_state_in_3 ? 8'h34 : _GEN_919; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_921 = 8'h99 == io_state_in_3 ? 8'h3d : _GEN_920; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_922 = 8'h9a == io_state_in_3 ? 8'h26 : _GEN_921; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_923 = 8'h9b == io_state_in_3 ? 8'h2f : _GEN_922; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_924 = 8'h9c == io_state_in_3 ? 8'h10 : _GEN_923; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_925 = 8'h9d == io_state_in_3 ? 8'h19 : _GEN_924; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_926 = 8'h9e == io_state_in_3 ? 8'h2 : _GEN_925; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_927 = 8'h9f == io_state_in_3 ? 8'hb : _GEN_926; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_928 = 8'ha0 == io_state_in_3 ? 8'hd7 : _GEN_927; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_929 = 8'ha1 == io_state_in_3 ? 8'hde : _GEN_928; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_930 = 8'ha2 == io_state_in_3 ? 8'hc5 : _GEN_929; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_931 = 8'ha3 == io_state_in_3 ? 8'hcc : _GEN_930; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_932 = 8'ha4 == io_state_in_3 ? 8'hf3 : _GEN_931; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_933 = 8'ha5 == io_state_in_3 ? 8'hfa : _GEN_932; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_934 = 8'ha6 == io_state_in_3 ? 8'he1 : _GEN_933; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_935 = 8'ha7 == io_state_in_3 ? 8'he8 : _GEN_934; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_936 = 8'ha8 == io_state_in_3 ? 8'h9f : _GEN_935; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_937 = 8'ha9 == io_state_in_3 ? 8'h96 : _GEN_936; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_938 = 8'haa == io_state_in_3 ? 8'h8d : _GEN_937; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_939 = 8'hab == io_state_in_3 ? 8'h84 : _GEN_938; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_940 = 8'hac == io_state_in_3 ? 8'hbb : _GEN_939; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_941 = 8'had == io_state_in_3 ? 8'hb2 : _GEN_940; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_942 = 8'hae == io_state_in_3 ? 8'ha9 : _GEN_941; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_943 = 8'haf == io_state_in_3 ? 8'ha0 : _GEN_942; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_944 = 8'hb0 == io_state_in_3 ? 8'h47 : _GEN_943; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_945 = 8'hb1 == io_state_in_3 ? 8'h4e : _GEN_944; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_946 = 8'hb2 == io_state_in_3 ? 8'h55 : _GEN_945; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_947 = 8'hb3 == io_state_in_3 ? 8'h5c : _GEN_946; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_948 = 8'hb4 == io_state_in_3 ? 8'h63 : _GEN_947; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_949 = 8'hb5 == io_state_in_3 ? 8'h6a : _GEN_948; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_950 = 8'hb6 == io_state_in_3 ? 8'h71 : _GEN_949; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_951 = 8'hb7 == io_state_in_3 ? 8'h78 : _GEN_950; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_952 = 8'hb8 == io_state_in_3 ? 8'hf : _GEN_951; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_953 = 8'hb9 == io_state_in_3 ? 8'h6 : _GEN_952; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_954 = 8'hba == io_state_in_3 ? 8'h1d : _GEN_953; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_955 = 8'hbb == io_state_in_3 ? 8'h14 : _GEN_954; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_956 = 8'hbc == io_state_in_3 ? 8'h2b : _GEN_955; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_957 = 8'hbd == io_state_in_3 ? 8'h22 : _GEN_956; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_958 = 8'hbe == io_state_in_3 ? 8'h39 : _GEN_957; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_959 = 8'hbf == io_state_in_3 ? 8'h30 : _GEN_958; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_960 = 8'hc0 == io_state_in_3 ? 8'h9a : _GEN_959; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_961 = 8'hc1 == io_state_in_3 ? 8'h93 : _GEN_960; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_962 = 8'hc2 == io_state_in_3 ? 8'h88 : _GEN_961; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_963 = 8'hc3 == io_state_in_3 ? 8'h81 : _GEN_962; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_964 = 8'hc4 == io_state_in_3 ? 8'hbe : _GEN_963; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_965 = 8'hc5 == io_state_in_3 ? 8'hb7 : _GEN_964; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_966 = 8'hc6 == io_state_in_3 ? 8'hac : _GEN_965; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_967 = 8'hc7 == io_state_in_3 ? 8'ha5 : _GEN_966; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_968 = 8'hc8 == io_state_in_3 ? 8'hd2 : _GEN_967; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_969 = 8'hc9 == io_state_in_3 ? 8'hdb : _GEN_968; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_970 = 8'hca == io_state_in_3 ? 8'hc0 : _GEN_969; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_971 = 8'hcb == io_state_in_3 ? 8'hc9 : _GEN_970; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_972 = 8'hcc == io_state_in_3 ? 8'hf6 : _GEN_971; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_973 = 8'hcd == io_state_in_3 ? 8'hff : _GEN_972; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_974 = 8'hce == io_state_in_3 ? 8'he4 : _GEN_973; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_975 = 8'hcf == io_state_in_3 ? 8'hed : _GEN_974; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_976 = 8'hd0 == io_state_in_3 ? 8'ha : _GEN_975; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_977 = 8'hd1 == io_state_in_3 ? 8'h3 : _GEN_976; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_978 = 8'hd2 == io_state_in_3 ? 8'h18 : _GEN_977; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_979 = 8'hd3 == io_state_in_3 ? 8'h11 : _GEN_978; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_980 = 8'hd4 == io_state_in_3 ? 8'h2e : _GEN_979; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_981 = 8'hd5 == io_state_in_3 ? 8'h27 : _GEN_980; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_982 = 8'hd6 == io_state_in_3 ? 8'h3c : _GEN_981; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_983 = 8'hd7 == io_state_in_3 ? 8'h35 : _GEN_982; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_984 = 8'hd8 == io_state_in_3 ? 8'h42 : _GEN_983; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_985 = 8'hd9 == io_state_in_3 ? 8'h4b : _GEN_984; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_986 = 8'hda == io_state_in_3 ? 8'h50 : _GEN_985; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_987 = 8'hdb == io_state_in_3 ? 8'h59 : _GEN_986; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_988 = 8'hdc == io_state_in_3 ? 8'h66 : _GEN_987; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_989 = 8'hdd == io_state_in_3 ? 8'h6f : _GEN_988; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_990 = 8'hde == io_state_in_3 ? 8'h74 : _GEN_989; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_991 = 8'hdf == io_state_in_3 ? 8'h7d : _GEN_990; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_992 = 8'he0 == io_state_in_3 ? 8'ha1 : _GEN_991; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_993 = 8'he1 == io_state_in_3 ? 8'ha8 : _GEN_992; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_994 = 8'he2 == io_state_in_3 ? 8'hb3 : _GEN_993; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_995 = 8'he3 == io_state_in_3 ? 8'hba : _GEN_994; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_996 = 8'he4 == io_state_in_3 ? 8'h85 : _GEN_995; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_997 = 8'he5 == io_state_in_3 ? 8'h8c : _GEN_996; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_998 = 8'he6 == io_state_in_3 ? 8'h97 : _GEN_997; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_999 = 8'he7 == io_state_in_3 ? 8'h9e : _GEN_998; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1000 = 8'he8 == io_state_in_3 ? 8'he9 : _GEN_999; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1001 = 8'he9 == io_state_in_3 ? 8'he0 : _GEN_1000; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1002 = 8'hea == io_state_in_3 ? 8'hfb : _GEN_1001; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1003 = 8'heb == io_state_in_3 ? 8'hf2 : _GEN_1002; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1004 = 8'hec == io_state_in_3 ? 8'hcd : _GEN_1003; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1005 = 8'hed == io_state_in_3 ? 8'hc4 : _GEN_1004; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1006 = 8'hee == io_state_in_3 ? 8'hdf : _GEN_1005; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1007 = 8'hef == io_state_in_3 ? 8'hd6 : _GEN_1006; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1008 = 8'hf0 == io_state_in_3 ? 8'h31 : _GEN_1007; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1009 = 8'hf1 == io_state_in_3 ? 8'h38 : _GEN_1008; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1010 = 8'hf2 == io_state_in_3 ? 8'h23 : _GEN_1009; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1011 = 8'hf3 == io_state_in_3 ? 8'h2a : _GEN_1010; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1012 = 8'hf4 == io_state_in_3 ? 8'h15 : _GEN_1011; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1013 = 8'hf5 == io_state_in_3 ? 8'h1c : _GEN_1012; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1014 = 8'hf6 == io_state_in_3 ? 8'h7 : _GEN_1013; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1015 = 8'hf7 == io_state_in_3 ? 8'he : _GEN_1014; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1016 = 8'hf8 == io_state_in_3 ? 8'h79 : _GEN_1015; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1017 = 8'hf9 == io_state_in_3 ? 8'h70 : _GEN_1016; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1018 = 8'hfa == io_state_in_3 ? 8'h6b : _GEN_1017; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1019 = 8'hfb == io_state_in_3 ? 8'h62 : _GEN_1018; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1020 = 8'hfc == io_state_in_3 ? 8'h5d : _GEN_1019; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1021 = 8'hfd == io_state_in_3 ? 8'h54 : _GEN_1020; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1022 = 8'hfe == io_state_in_3 ? 8'h4f : _GEN_1021; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1023 = 8'hff == io_state_in_3 ? 8'h46 : _GEN_1022; // @[InvMixColumns.scala 126:{89,89}]
  wire [7:0] _GEN_1025 = 8'h1 == io_state_in_0 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1026 = 8'h2 == io_state_in_0 ? 8'h12 : _GEN_1025; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1027 = 8'h3 == io_state_in_0 ? 8'h1b : _GEN_1026; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1028 = 8'h4 == io_state_in_0 ? 8'h24 : _GEN_1027; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1029 = 8'h5 == io_state_in_0 ? 8'h2d : _GEN_1028; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1030 = 8'h6 == io_state_in_0 ? 8'h36 : _GEN_1029; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1031 = 8'h7 == io_state_in_0 ? 8'h3f : _GEN_1030; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1032 = 8'h8 == io_state_in_0 ? 8'h48 : _GEN_1031; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1033 = 8'h9 == io_state_in_0 ? 8'h41 : _GEN_1032; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1034 = 8'ha == io_state_in_0 ? 8'h5a : _GEN_1033; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1035 = 8'hb == io_state_in_0 ? 8'h53 : _GEN_1034; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1036 = 8'hc == io_state_in_0 ? 8'h6c : _GEN_1035; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1037 = 8'hd == io_state_in_0 ? 8'h65 : _GEN_1036; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1038 = 8'he == io_state_in_0 ? 8'h7e : _GEN_1037; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1039 = 8'hf == io_state_in_0 ? 8'h77 : _GEN_1038; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1040 = 8'h10 == io_state_in_0 ? 8'h90 : _GEN_1039; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1041 = 8'h11 == io_state_in_0 ? 8'h99 : _GEN_1040; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1042 = 8'h12 == io_state_in_0 ? 8'h82 : _GEN_1041; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1043 = 8'h13 == io_state_in_0 ? 8'h8b : _GEN_1042; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1044 = 8'h14 == io_state_in_0 ? 8'hb4 : _GEN_1043; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1045 = 8'h15 == io_state_in_0 ? 8'hbd : _GEN_1044; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1046 = 8'h16 == io_state_in_0 ? 8'ha6 : _GEN_1045; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1047 = 8'h17 == io_state_in_0 ? 8'haf : _GEN_1046; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1048 = 8'h18 == io_state_in_0 ? 8'hd8 : _GEN_1047; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1049 = 8'h19 == io_state_in_0 ? 8'hd1 : _GEN_1048; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1050 = 8'h1a == io_state_in_0 ? 8'hca : _GEN_1049; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1051 = 8'h1b == io_state_in_0 ? 8'hc3 : _GEN_1050; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1052 = 8'h1c == io_state_in_0 ? 8'hfc : _GEN_1051; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1053 = 8'h1d == io_state_in_0 ? 8'hf5 : _GEN_1052; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1054 = 8'h1e == io_state_in_0 ? 8'hee : _GEN_1053; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1055 = 8'h1f == io_state_in_0 ? 8'he7 : _GEN_1054; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1056 = 8'h20 == io_state_in_0 ? 8'h3b : _GEN_1055; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1057 = 8'h21 == io_state_in_0 ? 8'h32 : _GEN_1056; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1058 = 8'h22 == io_state_in_0 ? 8'h29 : _GEN_1057; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1059 = 8'h23 == io_state_in_0 ? 8'h20 : _GEN_1058; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1060 = 8'h24 == io_state_in_0 ? 8'h1f : _GEN_1059; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1061 = 8'h25 == io_state_in_0 ? 8'h16 : _GEN_1060; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1062 = 8'h26 == io_state_in_0 ? 8'hd : _GEN_1061; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1063 = 8'h27 == io_state_in_0 ? 8'h4 : _GEN_1062; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1064 = 8'h28 == io_state_in_0 ? 8'h73 : _GEN_1063; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1065 = 8'h29 == io_state_in_0 ? 8'h7a : _GEN_1064; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1066 = 8'h2a == io_state_in_0 ? 8'h61 : _GEN_1065; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1067 = 8'h2b == io_state_in_0 ? 8'h68 : _GEN_1066; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1068 = 8'h2c == io_state_in_0 ? 8'h57 : _GEN_1067; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1069 = 8'h2d == io_state_in_0 ? 8'h5e : _GEN_1068; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1070 = 8'h2e == io_state_in_0 ? 8'h45 : _GEN_1069; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1071 = 8'h2f == io_state_in_0 ? 8'h4c : _GEN_1070; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1072 = 8'h30 == io_state_in_0 ? 8'hab : _GEN_1071; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1073 = 8'h31 == io_state_in_0 ? 8'ha2 : _GEN_1072; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1074 = 8'h32 == io_state_in_0 ? 8'hb9 : _GEN_1073; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1075 = 8'h33 == io_state_in_0 ? 8'hb0 : _GEN_1074; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1076 = 8'h34 == io_state_in_0 ? 8'h8f : _GEN_1075; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1077 = 8'h35 == io_state_in_0 ? 8'h86 : _GEN_1076; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1078 = 8'h36 == io_state_in_0 ? 8'h9d : _GEN_1077; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1079 = 8'h37 == io_state_in_0 ? 8'h94 : _GEN_1078; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1080 = 8'h38 == io_state_in_0 ? 8'he3 : _GEN_1079; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1081 = 8'h39 == io_state_in_0 ? 8'hea : _GEN_1080; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1082 = 8'h3a == io_state_in_0 ? 8'hf1 : _GEN_1081; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1083 = 8'h3b == io_state_in_0 ? 8'hf8 : _GEN_1082; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1084 = 8'h3c == io_state_in_0 ? 8'hc7 : _GEN_1083; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1085 = 8'h3d == io_state_in_0 ? 8'hce : _GEN_1084; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1086 = 8'h3e == io_state_in_0 ? 8'hd5 : _GEN_1085; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1087 = 8'h3f == io_state_in_0 ? 8'hdc : _GEN_1086; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1088 = 8'h40 == io_state_in_0 ? 8'h76 : _GEN_1087; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1089 = 8'h41 == io_state_in_0 ? 8'h7f : _GEN_1088; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1090 = 8'h42 == io_state_in_0 ? 8'h64 : _GEN_1089; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1091 = 8'h43 == io_state_in_0 ? 8'h6d : _GEN_1090; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1092 = 8'h44 == io_state_in_0 ? 8'h52 : _GEN_1091; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1093 = 8'h45 == io_state_in_0 ? 8'h5b : _GEN_1092; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1094 = 8'h46 == io_state_in_0 ? 8'h40 : _GEN_1093; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1095 = 8'h47 == io_state_in_0 ? 8'h49 : _GEN_1094; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1096 = 8'h48 == io_state_in_0 ? 8'h3e : _GEN_1095; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1097 = 8'h49 == io_state_in_0 ? 8'h37 : _GEN_1096; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1098 = 8'h4a == io_state_in_0 ? 8'h2c : _GEN_1097; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1099 = 8'h4b == io_state_in_0 ? 8'h25 : _GEN_1098; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1100 = 8'h4c == io_state_in_0 ? 8'h1a : _GEN_1099; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1101 = 8'h4d == io_state_in_0 ? 8'h13 : _GEN_1100; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1102 = 8'h4e == io_state_in_0 ? 8'h8 : _GEN_1101; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1103 = 8'h4f == io_state_in_0 ? 8'h1 : _GEN_1102; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1104 = 8'h50 == io_state_in_0 ? 8'he6 : _GEN_1103; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1105 = 8'h51 == io_state_in_0 ? 8'hef : _GEN_1104; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1106 = 8'h52 == io_state_in_0 ? 8'hf4 : _GEN_1105; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1107 = 8'h53 == io_state_in_0 ? 8'hfd : _GEN_1106; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1108 = 8'h54 == io_state_in_0 ? 8'hc2 : _GEN_1107; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1109 = 8'h55 == io_state_in_0 ? 8'hcb : _GEN_1108; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1110 = 8'h56 == io_state_in_0 ? 8'hd0 : _GEN_1109; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1111 = 8'h57 == io_state_in_0 ? 8'hd9 : _GEN_1110; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1112 = 8'h58 == io_state_in_0 ? 8'hae : _GEN_1111; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1113 = 8'h59 == io_state_in_0 ? 8'ha7 : _GEN_1112; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1114 = 8'h5a == io_state_in_0 ? 8'hbc : _GEN_1113; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1115 = 8'h5b == io_state_in_0 ? 8'hb5 : _GEN_1114; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1116 = 8'h5c == io_state_in_0 ? 8'h8a : _GEN_1115; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1117 = 8'h5d == io_state_in_0 ? 8'h83 : _GEN_1116; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1118 = 8'h5e == io_state_in_0 ? 8'h98 : _GEN_1117; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1119 = 8'h5f == io_state_in_0 ? 8'h91 : _GEN_1118; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1120 = 8'h60 == io_state_in_0 ? 8'h4d : _GEN_1119; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1121 = 8'h61 == io_state_in_0 ? 8'h44 : _GEN_1120; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1122 = 8'h62 == io_state_in_0 ? 8'h5f : _GEN_1121; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1123 = 8'h63 == io_state_in_0 ? 8'h56 : _GEN_1122; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1124 = 8'h64 == io_state_in_0 ? 8'h69 : _GEN_1123; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1125 = 8'h65 == io_state_in_0 ? 8'h60 : _GEN_1124; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1126 = 8'h66 == io_state_in_0 ? 8'h7b : _GEN_1125; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1127 = 8'h67 == io_state_in_0 ? 8'h72 : _GEN_1126; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1128 = 8'h68 == io_state_in_0 ? 8'h5 : _GEN_1127; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1129 = 8'h69 == io_state_in_0 ? 8'hc : _GEN_1128; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1130 = 8'h6a == io_state_in_0 ? 8'h17 : _GEN_1129; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1131 = 8'h6b == io_state_in_0 ? 8'h1e : _GEN_1130; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1132 = 8'h6c == io_state_in_0 ? 8'h21 : _GEN_1131; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1133 = 8'h6d == io_state_in_0 ? 8'h28 : _GEN_1132; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1134 = 8'h6e == io_state_in_0 ? 8'h33 : _GEN_1133; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1135 = 8'h6f == io_state_in_0 ? 8'h3a : _GEN_1134; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1136 = 8'h70 == io_state_in_0 ? 8'hdd : _GEN_1135; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1137 = 8'h71 == io_state_in_0 ? 8'hd4 : _GEN_1136; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1138 = 8'h72 == io_state_in_0 ? 8'hcf : _GEN_1137; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1139 = 8'h73 == io_state_in_0 ? 8'hc6 : _GEN_1138; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1140 = 8'h74 == io_state_in_0 ? 8'hf9 : _GEN_1139; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1141 = 8'h75 == io_state_in_0 ? 8'hf0 : _GEN_1140; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1142 = 8'h76 == io_state_in_0 ? 8'heb : _GEN_1141; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1143 = 8'h77 == io_state_in_0 ? 8'he2 : _GEN_1142; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1144 = 8'h78 == io_state_in_0 ? 8'h95 : _GEN_1143; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1145 = 8'h79 == io_state_in_0 ? 8'h9c : _GEN_1144; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1146 = 8'h7a == io_state_in_0 ? 8'h87 : _GEN_1145; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1147 = 8'h7b == io_state_in_0 ? 8'h8e : _GEN_1146; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1148 = 8'h7c == io_state_in_0 ? 8'hb1 : _GEN_1147; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1149 = 8'h7d == io_state_in_0 ? 8'hb8 : _GEN_1148; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1150 = 8'h7e == io_state_in_0 ? 8'ha3 : _GEN_1149; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1151 = 8'h7f == io_state_in_0 ? 8'haa : _GEN_1150; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1152 = 8'h80 == io_state_in_0 ? 8'hec : _GEN_1151; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1153 = 8'h81 == io_state_in_0 ? 8'he5 : _GEN_1152; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1154 = 8'h82 == io_state_in_0 ? 8'hfe : _GEN_1153; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1155 = 8'h83 == io_state_in_0 ? 8'hf7 : _GEN_1154; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1156 = 8'h84 == io_state_in_0 ? 8'hc8 : _GEN_1155; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1157 = 8'h85 == io_state_in_0 ? 8'hc1 : _GEN_1156; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1158 = 8'h86 == io_state_in_0 ? 8'hda : _GEN_1157; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1159 = 8'h87 == io_state_in_0 ? 8'hd3 : _GEN_1158; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1160 = 8'h88 == io_state_in_0 ? 8'ha4 : _GEN_1159; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1161 = 8'h89 == io_state_in_0 ? 8'had : _GEN_1160; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1162 = 8'h8a == io_state_in_0 ? 8'hb6 : _GEN_1161; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1163 = 8'h8b == io_state_in_0 ? 8'hbf : _GEN_1162; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1164 = 8'h8c == io_state_in_0 ? 8'h80 : _GEN_1163; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1165 = 8'h8d == io_state_in_0 ? 8'h89 : _GEN_1164; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1166 = 8'h8e == io_state_in_0 ? 8'h92 : _GEN_1165; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1167 = 8'h8f == io_state_in_0 ? 8'h9b : _GEN_1166; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1168 = 8'h90 == io_state_in_0 ? 8'h7c : _GEN_1167; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1169 = 8'h91 == io_state_in_0 ? 8'h75 : _GEN_1168; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1170 = 8'h92 == io_state_in_0 ? 8'h6e : _GEN_1169; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1171 = 8'h93 == io_state_in_0 ? 8'h67 : _GEN_1170; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1172 = 8'h94 == io_state_in_0 ? 8'h58 : _GEN_1171; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1173 = 8'h95 == io_state_in_0 ? 8'h51 : _GEN_1172; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1174 = 8'h96 == io_state_in_0 ? 8'h4a : _GEN_1173; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1175 = 8'h97 == io_state_in_0 ? 8'h43 : _GEN_1174; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1176 = 8'h98 == io_state_in_0 ? 8'h34 : _GEN_1175; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1177 = 8'h99 == io_state_in_0 ? 8'h3d : _GEN_1176; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1178 = 8'h9a == io_state_in_0 ? 8'h26 : _GEN_1177; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1179 = 8'h9b == io_state_in_0 ? 8'h2f : _GEN_1178; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1180 = 8'h9c == io_state_in_0 ? 8'h10 : _GEN_1179; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1181 = 8'h9d == io_state_in_0 ? 8'h19 : _GEN_1180; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1182 = 8'h9e == io_state_in_0 ? 8'h2 : _GEN_1181; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1183 = 8'h9f == io_state_in_0 ? 8'hb : _GEN_1182; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1184 = 8'ha0 == io_state_in_0 ? 8'hd7 : _GEN_1183; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1185 = 8'ha1 == io_state_in_0 ? 8'hde : _GEN_1184; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1186 = 8'ha2 == io_state_in_0 ? 8'hc5 : _GEN_1185; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1187 = 8'ha3 == io_state_in_0 ? 8'hcc : _GEN_1186; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1188 = 8'ha4 == io_state_in_0 ? 8'hf3 : _GEN_1187; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1189 = 8'ha5 == io_state_in_0 ? 8'hfa : _GEN_1188; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1190 = 8'ha6 == io_state_in_0 ? 8'he1 : _GEN_1189; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1191 = 8'ha7 == io_state_in_0 ? 8'he8 : _GEN_1190; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1192 = 8'ha8 == io_state_in_0 ? 8'h9f : _GEN_1191; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1193 = 8'ha9 == io_state_in_0 ? 8'h96 : _GEN_1192; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1194 = 8'haa == io_state_in_0 ? 8'h8d : _GEN_1193; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1195 = 8'hab == io_state_in_0 ? 8'h84 : _GEN_1194; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1196 = 8'hac == io_state_in_0 ? 8'hbb : _GEN_1195; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1197 = 8'had == io_state_in_0 ? 8'hb2 : _GEN_1196; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1198 = 8'hae == io_state_in_0 ? 8'ha9 : _GEN_1197; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1199 = 8'haf == io_state_in_0 ? 8'ha0 : _GEN_1198; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1200 = 8'hb0 == io_state_in_0 ? 8'h47 : _GEN_1199; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1201 = 8'hb1 == io_state_in_0 ? 8'h4e : _GEN_1200; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1202 = 8'hb2 == io_state_in_0 ? 8'h55 : _GEN_1201; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1203 = 8'hb3 == io_state_in_0 ? 8'h5c : _GEN_1202; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1204 = 8'hb4 == io_state_in_0 ? 8'h63 : _GEN_1203; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1205 = 8'hb5 == io_state_in_0 ? 8'h6a : _GEN_1204; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1206 = 8'hb6 == io_state_in_0 ? 8'h71 : _GEN_1205; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1207 = 8'hb7 == io_state_in_0 ? 8'h78 : _GEN_1206; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1208 = 8'hb8 == io_state_in_0 ? 8'hf : _GEN_1207; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1209 = 8'hb9 == io_state_in_0 ? 8'h6 : _GEN_1208; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1210 = 8'hba == io_state_in_0 ? 8'h1d : _GEN_1209; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1211 = 8'hbb == io_state_in_0 ? 8'h14 : _GEN_1210; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1212 = 8'hbc == io_state_in_0 ? 8'h2b : _GEN_1211; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1213 = 8'hbd == io_state_in_0 ? 8'h22 : _GEN_1212; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1214 = 8'hbe == io_state_in_0 ? 8'h39 : _GEN_1213; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1215 = 8'hbf == io_state_in_0 ? 8'h30 : _GEN_1214; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1216 = 8'hc0 == io_state_in_0 ? 8'h9a : _GEN_1215; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1217 = 8'hc1 == io_state_in_0 ? 8'h93 : _GEN_1216; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1218 = 8'hc2 == io_state_in_0 ? 8'h88 : _GEN_1217; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1219 = 8'hc3 == io_state_in_0 ? 8'h81 : _GEN_1218; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1220 = 8'hc4 == io_state_in_0 ? 8'hbe : _GEN_1219; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1221 = 8'hc5 == io_state_in_0 ? 8'hb7 : _GEN_1220; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1222 = 8'hc6 == io_state_in_0 ? 8'hac : _GEN_1221; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1223 = 8'hc7 == io_state_in_0 ? 8'ha5 : _GEN_1222; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1224 = 8'hc8 == io_state_in_0 ? 8'hd2 : _GEN_1223; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1225 = 8'hc9 == io_state_in_0 ? 8'hdb : _GEN_1224; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1226 = 8'hca == io_state_in_0 ? 8'hc0 : _GEN_1225; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1227 = 8'hcb == io_state_in_0 ? 8'hc9 : _GEN_1226; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1228 = 8'hcc == io_state_in_0 ? 8'hf6 : _GEN_1227; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1229 = 8'hcd == io_state_in_0 ? 8'hff : _GEN_1228; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1230 = 8'hce == io_state_in_0 ? 8'he4 : _GEN_1229; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1231 = 8'hcf == io_state_in_0 ? 8'hed : _GEN_1230; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1232 = 8'hd0 == io_state_in_0 ? 8'ha : _GEN_1231; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1233 = 8'hd1 == io_state_in_0 ? 8'h3 : _GEN_1232; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1234 = 8'hd2 == io_state_in_0 ? 8'h18 : _GEN_1233; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1235 = 8'hd3 == io_state_in_0 ? 8'h11 : _GEN_1234; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1236 = 8'hd4 == io_state_in_0 ? 8'h2e : _GEN_1235; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1237 = 8'hd5 == io_state_in_0 ? 8'h27 : _GEN_1236; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1238 = 8'hd6 == io_state_in_0 ? 8'h3c : _GEN_1237; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1239 = 8'hd7 == io_state_in_0 ? 8'h35 : _GEN_1238; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1240 = 8'hd8 == io_state_in_0 ? 8'h42 : _GEN_1239; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1241 = 8'hd9 == io_state_in_0 ? 8'h4b : _GEN_1240; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1242 = 8'hda == io_state_in_0 ? 8'h50 : _GEN_1241; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1243 = 8'hdb == io_state_in_0 ? 8'h59 : _GEN_1242; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1244 = 8'hdc == io_state_in_0 ? 8'h66 : _GEN_1243; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1245 = 8'hdd == io_state_in_0 ? 8'h6f : _GEN_1244; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1246 = 8'hde == io_state_in_0 ? 8'h74 : _GEN_1245; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1247 = 8'hdf == io_state_in_0 ? 8'h7d : _GEN_1246; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1248 = 8'he0 == io_state_in_0 ? 8'ha1 : _GEN_1247; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1249 = 8'he1 == io_state_in_0 ? 8'ha8 : _GEN_1248; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1250 = 8'he2 == io_state_in_0 ? 8'hb3 : _GEN_1249; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1251 = 8'he3 == io_state_in_0 ? 8'hba : _GEN_1250; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1252 = 8'he4 == io_state_in_0 ? 8'h85 : _GEN_1251; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1253 = 8'he5 == io_state_in_0 ? 8'h8c : _GEN_1252; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1254 = 8'he6 == io_state_in_0 ? 8'h97 : _GEN_1253; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1255 = 8'he7 == io_state_in_0 ? 8'h9e : _GEN_1254; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1256 = 8'he8 == io_state_in_0 ? 8'he9 : _GEN_1255; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1257 = 8'he9 == io_state_in_0 ? 8'he0 : _GEN_1256; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1258 = 8'hea == io_state_in_0 ? 8'hfb : _GEN_1257; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1259 = 8'heb == io_state_in_0 ? 8'hf2 : _GEN_1258; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1260 = 8'hec == io_state_in_0 ? 8'hcd : _GEN_1259; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1261 = 8'hed == io_state_in_0 ? 8'hc4 : _GEN_1260; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1262 = 8'hee == io_state_in_0 ? 8'hdf : _GEN_1261; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1263 = 8'hef == io_state_in_0 ? 8'hd6 : _GEN_1262; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1264 = 8'hf0 == io_state_in_0 ? 8'h31 : _GEN_1263; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1265 = 8'hf1 == io_state_in_0 ? 8'h38 : _GEN_1264; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1266 = 8'hf2 == io_state_in_0 ? 8'h23 : _GEN_1265; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1267 = 8'hf3 == io_state_in_0 ? 8'h2a : _GEN_1266; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1268 = 8'hf4 == io_state_in_0 ? 8'h15 : _GEN_1267; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1269 = 8'hf5 == io_state_in_0 ? 8'h1c : _GEN_1268; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1270 = 8'hf6 == io_state_in_0 ? 8'h7 : _GEN_1269; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1271 = 8'hf7 == io_state_in_0 ? 8'he : _GEN_1270; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1272 = 8'hf8 == io_state_in_0 ? 8'h79 : _GEN_1271; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1273 = 8'hf9 == io_state_in_0 ? 8'h70 : _GEN_1272; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1274 = 8'hfa == io_state_in_0 ? 8'h6b : _GEN_1273; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1275 = 8'hfb == io_state_in_0 ? 8'h62 : _GEN_1274; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1276 = 8'hfc == io_state_in_0 ? 8'h5d : _GEN_1275; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1277 = 8'hfd == io_state_in_0 ? 8'h54 : _GEN_1276; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1278 = 8'hfe == io_state_in_0 ? 8'h4f : _GEN_1277; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1279 = 8'hff == io_state_in_0 ? 8'h46 : _GEN_1278; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1281 = 8'h1 == io_state_in_1 ? 8'he : 8'h0; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1282 = 8'h2 == io_state_in_1 ? 8'h1c : _GEN_1281; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1283 = 8'h3 == io_state_in_1 ? 8'h12 : _GEN_1282; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1284 = 8'h4 == io_state_in_1 ? 8'h38 : _GEN_1283; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1285 = 8'h5 == io_state_in_1 ? 8'h36 : _GEN_1284; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1286 = 8'h6 == io_state_in_1 ? 8'h24 : _GEN_1285; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1287 = 8'h7 == io_state_in_1 ? 8'h2a : _GEN_1286; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1288 = 8'h8 == io_state_in_1 ? 8'h70 : _GEN_1287; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1289 = 8'h9 == io_state_in_1 ? 8'h7e : _GEN_1288; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1290 = 8'ha == io_state_in_1 ? 8'h6c : _GEN_1289; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1291 = 8'hb == io_state_in_1 ? 8'h62 : _GEN_1290; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1292 = 8'hc == io_state_in_1 ? 8'h48 : _GEN_1291; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1293 = 8'hd == io_state_in_1 ? 8'h46 : _GEN_1292; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1294 = 8'he == io_state_in_1 ? 8'h54 : _GEN_1293; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1295 = 8'hf == io_state_in_1 ? 8'h5a : _GEN_1294; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1296 = 8'h10 == io_state_in_1 ? 8'he0 : _GEN_1295; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1297 = 8'h11 == io_state_in_1 ? 8'hee : _GEN_1296; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1298 = 8'h12 == io_state_in_1 ? 8'hfc : _GEN_1297; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1299 = 8'h13 == io_state_in_1 ? 8'hf2 : _GEN_1298; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1300 = 8'h14 == io_state_in_1 ? 8'hd8 : _GEN_1299; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1301 = 8'h15 == io_state_in_1 ? 8'hd6 : _GEN_1300; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1302 = 8'h16 == io_state_in_1 ? 8'hc4 : _GEN_1301; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1303 = 8'h17 == io_state_in_1 ? 8'hca : _GEN_1302; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1304 = 8'h18 == io_state_in_1 ? 8'h90 : _GEN_1303; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1305 = 8'h19 == io_state_in_1 ? 8'h9e : _GEN_1304; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1306 = 8'h1a == io_state_in_1 ? 8'h8c : _GEN_1305; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1307 = 8'h1b == io_state_in_1 ? 8'h82 : _GEN_1306; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1308 = 8'h1c == io_state_in_1 ? 8'ha8 : _GEN_1307; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1309 = 8'h1d == io_state_in_1 ? 8'ha6 : _GEN_1308; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1310 = 8'h1e == io_state_in_1 ? 8'hb4 : _GEN_1309; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1311 = 8'h1f == io_state_in_1 ? 8'hba : _GEN_1310; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1312 = 8'h20 == io_state_in_1 ? 8'hdb : _GEN_1311; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1313 = 8'h21 == io_state_in_1 ? 8'hd5 : _GEN_1312; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1314 = 8'h22 == io_state_in_1 ? 8'hc7 : _GEN_1313; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1315 = 8'h23 == io_state_in_1 ? 8'hc9 : _GEN_1314; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1316 = 8'h24 == io_state_in_1 ? 8'he3 : _GEN_1315; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1317 = 8'h25 == io_state_in_1 ? 8'hed : _GEN_1316; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1318 = 8'h26 == io_state_in_1 ? 8'hff : _GEN_1317; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1319 = 8'h27 == io_state_in_1 ? 8'hf1 : _GEN_1318; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1320 = 8'h28 == io_state_in_1 ? 8'hab : _GEN_1319; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1321 = 8'h29 == io_state_in_1 ? 8'ha5 : _GEN_1320; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1322 = 8'h2a == io_state_in_1 ? 8'hb7 : _GEN_1321; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1323 = 8'h2b == io_state_in_1 ? 8'hb9 : _GEN_1322; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1324 = 8'h2c == io_state_in_1 ? 8'h93 : _GEN_1323; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1325 = 8'h2d == io_state_in_1 ? 8'h9d : _GEN_1324; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1326 = 8'h2e == io_state_in_1 ? 8'h8f : _GEN_1325; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1327 = 8'h2f == io_state_in_1 ? 8'h81 : _GEN_1326; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1328 = 8'h30 == io_state_in_1 ? 8'h3b : _GEN_1327; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1329 = 8'h31 == io_state_in_1 ? 8'h35 : _GEN_1328; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1330 = 8'h32 == io_state_in_1 ? 8'h27 : _GEN_1329; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1331 = 8'h33 == io_state_in_1 ? 8'h29 : _GEN_1330; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1332 = 8'h34 == io_state_in_1 ? 8'h3 : _GEN_1331; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1333 = 8'h35 == io_state_in_1 ? 8'hd : _GEN_1332; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1334 = 8'h36 == io_state_in_1 ? 8'h1f : _GEN_1333; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1335 = 8'h37 == io_state_in_1 ? 8'h11 : _GEN_1334; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1336 = 8'h38 == io_state_in_1 ? 8'h4b : _GEN_1335; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1337 = 8'h39 == io_state_in_1 ? 8'h45 : _GEN_1336; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1338 = 8'h3a == io_state_in_1 ? 8'h57 : _GEN_1337; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1339 = 8'h3b == io_state_in_1 ? 8'h59 : _GEN_1338; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1340 = 8'h3c == io_state_in_1 ? 8'h73 : _GEN_1339; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1341 = 8'h3d == io_state_in_1 ? 8'h7d : _GEN_1340; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1342 = 8'h3e == io_state_in_1 ? 8'h6f : _GEN_1341; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1343 = 8'h3f == io_state_in_1 ? 8'h61 : _GEN_1342; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1344 = 8'h40 == io_state_in_1 ? 8'had : _GEN_1343; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1345 = 8'h41 == io_state_in_1 ? 8'ha3 : _GEN_1344; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1346 = 8'h42 == io_state_in_1 ? 8'hb1 : _GEN_1345; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1347 = 8'h43 == io_state_in_1 ? 8'hbf : _GEN_1346; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1348 = 8'h44 == io_state_in_1 ? 8'h95 : _GEN_1347; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1349 = 8'h45 == io_state_in_1 ? 8'h9b : _GEN_1348; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1350 = 8'h46 == io_state_in_1 ? 8'h89 : _GEN_1349; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1351 = 8'h47 == io_state_in_1 ? 8'h87 : _GEN_1350; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1352 = 8'h48 == io_state_in_1 ? 8'hdd : _GEN_1351; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1353 = 8'h49 == io_state_in_1 ? 8'hd3 : _GEN_1352; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1354 = 8'h4a == io_state_in_1 ? 8'hc1 : _GEN_1353; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1355 = 8'h4b == io_state_in_1 ? 8'hcf : _GEN_1354; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1356 = 8'h4c == io_state_in_1 ? 8'he5 : _GEN_1355; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1357 = 8'h4d == io_state_in_1 ? 8'heb : _GEN_1356; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1358 = 8'h4e == io_state_in_1 ? 8'hf9 : _GEN_1357; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1359 = 8'h4f == io_state_in_1 ? 8'hf7 : _GEN_1358; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1360 = 8'h50 == io_state_in_1 ? 8'h4d : _GEN_1359; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1361 = 8'h51 == io_state_in_1 ? 8'h43 : _GEN_1360; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1362 = 8'h52 == io_state_in_1 ? 8'h51 : _GEN_1361; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1363 = 8'h53 == io_state_in_1 ? 8'h5f : _GEN_1362; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1364 = 8'h54 == io_state_in_1 ? 8'h75 : _GEN_1363; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1365 = 8'h55 == io_state_in_1 ? 8'h7b : _GEN_1364; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1366 = 8'h56 == io_state_in_1 ? 8'h69 : _GEN_1365; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1367 = 8'h57 == io_state_in_1 ? 8'h67 : _GEN_1366; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1368 = 8'h58 == io_state_in_1 ? 8'h3d : _GEN_1367; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1369 = 8'h59 == io_state_in_1 ? 8'h33 : _GEN_1368; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1370 = 8'h5a == io_state_in_1 ? 8'h21 : _GEN_1369; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1371 = 8'h5b == io_state_in_1 ? 8'h2f : _GEN_1370; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1372 = 8'h5c == io_state_in_1 ? 8'h5 : _GEN_1371; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1373 = 8'h5d == io_state_in_1 ? 8'hb : _GEN_1372; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1374 = 8'h5e == io_state_in_1 ? 8'h19 : _GEN_1373; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1375 = 8'h5f == io_state_in_1 ? 8'h17 : _GEN_1374; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1376 = 8'h60 == io_state_in_1 ? 8'h76 : _GEN_1375; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1377 = 8'h61 == io_state_in_1 ? 8'h78 : _GEN_1376; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1378 = 8'h62 == io_state_in_1 ? 8'h6a : _GEN_1377; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1379 = 8'h63 == io_state_in_1 ? 8'h64 : _GEN_1378; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1380 = 8'h64 == io_state_in_1 ? 8'h4e : _GEN_1379; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1381 = 8'h65 == io_state_in_1 ? 8'h40 : _GEN_1380; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1382 = 8'h66 == io_state_in_1 ? 8'h52 : _GEN_1381; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1383 = 8'h67 == io_state_in_1 ? 8'h5c : _GEN_1382; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1384 = 8'h68 == io_state_in_1 ? 8'h6 : _GEN_1383; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1385 = 8'h69 == io_state_in_1 ? 8'h8 : _GEN_1384; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1386 = 8'h6a == io_state_in_1 ? 8'h1a : _GEN_1385; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1387 = 8'h6b == io_state_in_1 ? 8'h14 : _GEN_1386; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1388 = 8'h6c == io_state_in_1 ? 8'h3e : _GEN_1387; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1389 = 8'h6d == io_state_in_1 ? 8'h30 : _GEN_1388; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1390 = 8'h6e == io_state_in_1 ? 8'h22 : _GEN_1389; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1391 = 8'h6f == io_state_in_1 ? 8'h2c : _GEN_1390; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1392 = 8'h70 == io_state_in_1 ? 8'h96 : _GEN_1391; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1393 = 8'h71 == io_state_in_1 ? 8'h98 : _GEN_1392; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1394 = 8'h72 == io_state_in_1 ? 8'h8a : _GEN_1393; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1395 = 8'h73 == io_state_in_1 ? 8'h84 : _GEN_1394; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1396 = 8'h74 == io_state_in_1 ? 8'hae : _GEN_1395; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1397 = 8'h75 == io_state_in_1 ? 8'ha0 : _GEN_1396; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1398 = 8'h76 == io_state_in_1 ? 8'hb2 : _GEN_1397; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1399 = 8'h77 == io_state_in_1 ? 8'hbc : _GEN_1398; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1400 = 8'h78 == io_state_in_1 ? 8'he6 : _GEN_1399; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1401 = 8'h79 == io_state_in_1 ? 8'he8 : _GEN_1400; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1402 = 8'h7a == io_state_in_1 ? 8'hfa : _GEN_1401; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1403 = 8'h7b == io_state_in_1 ? 8'hf4 : _GEN_1402; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1404 = 8'h7c == io_state_in_1 ? 8'hde : _GEN_1403; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1405 = 8'h7d == io_state_in_1 ? 8'hd0 : _GEN_1404; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1406 = 8'h7e == io_state_in_1 ? 8'hc2 : _GEN_1405; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1407 = 8'h7f == io_state_in_1 ? 8'hcc : _GEN_1406; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1408 = 8'h80 == io_state_in_1 ? 8'h41 : _GEN_1407; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1409 = 8'h81 == io_state_in_1 ? 8'h4f : _GEN_1408; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1410 = 8'h82 == io_state_in_1 ? 8'h5d : _GEN_1409; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1411 = 8'h83 == io_state_in_1 ? 8'h53 : _GEN_1410; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1412 = 8'h84 == io_state_in_1 ? 8'h79 : _GEN_1411; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1413 = 8'h85 == io_state_in_1 ? 8'h77 : _GEN_1412; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1414 = 8'h86 == io_state_in_1 ? 8'h65 : _GEN_1413; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1415 = 8'h87 == io_state_in_1 ? 8'h6b : _GEN_1414; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1416 = 8'h88 == io_state_in_1 ? 8'h31 : _GEN_1415; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1417 = 8'h89 == io_state_in_1 ? 8'h3f : _GEN_1416; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1418 = 8'h8a == io_state_in_1 ? 8'h2d : _GEN_1417; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1419 = 8'h8b == io_state_in_1 ? 8'h23 : _GEN_1418; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1420 = 8'h8c == io_state_in_1 ? 8'h9 : _GEN_1419; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1421 = 8'h8d == io_state_in_1 ? 8'h7 : _GEN_1420; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1422 = 8'h8e == io_state_in_1 ? 8'h15 : _GEN_1421; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1423 = 8'h8f == io_state_in_1 ? 8'h1b : _GEN_1422; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1424 = 8'h90 == io_state_in_1 ? 8'ha1 : _GEN_1423; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1425 = 8'h91 == io_state_in_1 ? 8'haf : _GEN_1424; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1426 = 8'h92 == io_state_in_1 ? 8'hbd : _GEN_1425; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1427 = 8'h93 == io_state_in_1 ? 8'hb3 : _GEN_1426; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1428 = 8'h94 == io_state_in_1 ? 8'h99 : _GEN_1427; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1429 = 8'h95 == io_state_in_1 ? 8'h97 : _GEN_1428; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1430 = 8'h96 == io_state_in_1 ? 8'h85 : _GEN_1429; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1431 = 8'h97 == io_state_in_1 ? 8'h8b : _GEN_1430; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1432 = 8'h98 == io_state_in_1 ? 8'hd1 : _GEN_1431; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1433 = 8'h99 == io_state_in_1 ? 8'hdf : _GEN_1432; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1434 = 8'h9a == io_state_in_1 ? 8'hcd : _GEN_1433; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1435 = 8'h9b == io_state_in_1 ? 8'hc3 : _GEN_1434; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1436 = 8'h9c == io_state_in_1 ? 8'he9 : _GEN_1435; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1437 = 8'h9d == io_state_in_1 ? 8'he7 : _GEN_1436; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1438 = 8'h9e == io_state_in_1 ? 8'hf5 : _GEN_1437; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1439 = 8'h9f == io_state_in_1 ? 8'hfb : _GEN_1438; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1440 = 8'ha0 == io_state_in_1 ? 8'h9a : _GEN_1439; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1441 = 8'ha1 == io_state_in_1 ? 8'h94 : _GEN_1440; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1442 = 8'ha2 == io_state_in_1 ? 8'h86 : _GEN_1441; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1443 = 8'ha3 == io_state_in_1 ? 8'h88 : _GEN_1442; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1444 = 8'ha4 == io_state_in_1 ? 8'ha2 : _GEN_1443; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1445 = 8'ha5 == io_state_in_1 ? 8'hac : _GEN_1444; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1446 = 8'ha6 == io_state_in_1 ? 8'hbe : _GEN_1445; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1447 = 8'ha7 == io_state_in_1 ? 8'hb0 : _GEN_1446; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1448 = 8'ha8 == io_state_in_1 ? 8'hea : _GEN_1447; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1449 = 8'ha9 == io_state_in_1 ? 8'he4 : _GEN_1448; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1450 = 8'haa == io_state_in_1 ? 8'hf6 : _GEN_1449; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1451 = 8'hab == io_state_in_1 ? 8'hf8 : _GEN_1450; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1452 = 8'hac == io_state_in_1 ? 8'hd2 : _GEN_1451; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1453 = 8'had == io_state_in_1 ? 8'hdc : _GEN_1452; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1454 = 8'hae == io_state_in_1 ? 8'hce : _GEN_1453; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1455 = 8'haf == io_state_in_1 ? 8'hc0 : _GEN_1454; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1456 = 8'hb0 == io_state_in_1 ? 8'h7a : _GEN_1455; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1457 = 8'hb1 == io_state_in_1 ? 8'h74 : _GEN_1456; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1458 = 8'hb2 == io_state_in_1 ? 8'h66 : _GEN_1457; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1459 = 8'hb3 == io_state_in_1 ? 8'h68 : _GEN_1458; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1460 = 8'hb4 == io_state_in_1 ? 8'h42 : _GEN_1459; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1461 = 8'hb5 == io_state_in_1 ? 8'h4c : _GEN_1460; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1462 = 8'hb6 == io_state_in_1 ? 8'h5e : _GEN_1461; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1463 = 8'hb7 == io_state_in_1 ? 8'h50 : _GEN_1462; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1464 = 8'hb8 == io_state_in_1 ? 8'ha : _GEN_1463; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1465 = 8'hb9 == io_state_in_1 ? 8'h4 : _GEN_1464; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1466 = 8'hba == io_state_in_1 ? 8'h16 : _GEN_1465; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1467 = 8'hbb == io_state_in_1 ? 8'h18 : _GEN_1466; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1468 = 8'hbc == io_state_in_1 ? 8'h32 : _GEN_1467; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1469 = 8'hbd == io_state_in_1 ? 8'h3c : _GEN_1468; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1470 = 8'hbe == io_state_in_1 ? 8'h2e : _GEN_1469; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1471 = 8'hbf == io_state_in_1 ? 8'h20 : _GEN_1470; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1472 = 8'hc0 == io_state_in_1 ? 8'hec : _GEN_1471; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1473 = 8'hc1 == io_state_in_1 ? 8'he2 : _GEN_1472; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1474 = 8'hc2 == io_state_in_1 ? 8'hf0 : _GEN_1473; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1475 = 8'hc3 == io_state_in_1 ? 8'hfe : _GEN_1474; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1476 = 8'hc4 == io_state_in_1 ? 8'hd4 : _GEN_1475; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1477 = 8'hc5 == io_state_in_1 ? 8'hda : _GEN_1476; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1478 = 8'hc6 == io_state_in_1 ? 8'hc8 : _GEN_1477; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1479 = 8'hc7 == io_state_in_1 ? 8'hc6 : _GEN_1478; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1480 = 8'hc8 == io_state_in_1 ? 8'h9c : _GEN_1479; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1481 = 8'hc9 == io_state_in_1 ? 8'h92 : _GEN_1480; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1482 = 8'hca == io_state_in_1 ? 8'h80 : _GEN_1481; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1483 = 8'hcb == io_state_in_1 ? 8'h8e : _GEN_1482; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1484 = 8'hcc == io_state_in_1 ? 8'ha4 : _GEN_1483; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1485 = 8'hcd == io_state_in_1 ? 8'haa : _GEN_1484; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1486 = 8'hce == io_state_in_1 ? 8'hb8 : _GEN_1485; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1487 = 8'hcf == io_state_in_1 ? 8'hb6 : _GEN_1486; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1488 = 8'hd0 == io_state_in_1 ? 8'hc : _GEN_1487; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1489 = 8'hd1 == io_state_in_1 ? 8'h2 : _GEN_1488; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1490 = 8'hd2 == io_state_in_1 ? 8'h10 : _GEN_1489; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1491 = 8'hd3 == io_state_in_1 ? 8'h1e : _GEN_1490; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1492 = 8'hd4 == io_state_in_1 ? 8'h34 : _GEN_1491; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1493 = 8'hd5 == io_state_in_1 ? 8'h3a : _GEN_1492; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1494 = 8'hd6 == io_state_in_1 ? 8'h28 : _GEN_1493; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1495 = 8'hd7 == io_state_in_1 ? 8'h26 : _GEN_1494; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1496 = 8'hd8 == io_state_in_1 ? 8'h7c : _GEN_1495; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1497 = 8'hd9 == io_state_in_1 ? 8'h72 : _GEN_1496; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1498 = 8'hda == io_state_in_1 ? 8'h60 : _GEN_1497; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1499 = 8'hdb == io_state_in_1 ? 8'h6e : _GEN_1498; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1500 = 8'hdc == io_state_in_1 ? 8'h44 : _GEN_1499; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1501 = 8'hdd == io_state_in_1 ? 8'h4a : _GEN_1500; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1502 = 8'hde == io_state_in_1 ? 8'h58 : _GEN_1501; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1503 = 8'hdf == io_state_in_1 ? 8'h56 : _GEN_1502; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1504 = 8'he0 == io_state_in_1 ? 8'h37 : _GEN_1503; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1505 = 8'he1 == io_state_in_1 ? 8'h39 : _GEN_1504; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1506 = 8'he2 == io_state_in_1 ? 8'h2b : _GEN_1505; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1507 = 8'he3 == io_state_in_1 ? 8'h25 : _GEN_1506; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1508 = 8'he4 == io_state_in_1 ? 8'hf : _GEN_1507; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1509 = 8'he5 == io_state_in_1 ? 8'h1 : _GEN_1508; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1510 = 8'he6 == io_state_in_1 ? 8'h13 : _GEN_1509; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1511 = 8'he7 == io_state_in_1 ? 8'h1d : _GEN_1510; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1512 = 8'he8 == io_state_in_1 ? 8'h47 : _GEN_1511; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1513 = 8'he9 == io_state_in_1 ? 8'h49 : _GEN_1512; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1514 = 8'hea == io_state_in_1 ? 8'h5b : _GEN_1513; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1515 = 8'heb == io_state_in_1 ? 8'h55 : _GEN_1514; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1516 = 8'hec == io_state_in_1 ? 8'h7f : _GEN_1515; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1517 = 8'hed == io_state_in_1 ? 8'h71 : _GEN_1516; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1518 = 8'hee == io_state_in_1 ? 8'h63 : _GEN_1517; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1519 = 8'hef == io_state_in_1 ? 8'h6d : _GEN_1518; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1520 = 8'hf0 == io_state_in_1 ? 8'hd7 : _GEN_1519; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1521 = 8'hf1 == io_state_in_1 ? 8'hd9 : _GEN_1520; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1522 = 8'hf2 == io_state_in_1 ? 8'hcb : _GEN_1521; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1523 = 8'hf3 == io_state_in_1 ? 8'hc5 : _GEN_1522; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1524 = 8'hf4 == io_state_in_1 ? 8'hef : _GEN_1523; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1525 = 8'hf5 == io_state_in_1 ? 8'he1 : _GEN_1524; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1526 = 8'hf6 == io_state_in_1 ? 8'hf3 : _GEN_1525; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1527 = 8'hf7 == io_state_in_1 ? 8'hfd : _GEN_1526; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1528 = 8'hf8 == io_state_in_1 ? 8'ha7 : _GEN_1527; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1529 = 8'hf9 == io_state_in_1 ? 8'ha9 : _GEN_1528; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1530 = 8'hfa == io_state_in_1 ? 8'hbb : _GEN_1529; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1531 = 8'hfb == io_state_in_1 ? 8'hb5 : _GEN_1530; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1532 = 8'hfc == io_state_in_1 ? 8'h9f : _GEN_1531; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1533 = 8'hfd == io_state_in_1 ? 8'h91 : _GEN_1532; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1534 = 8'hfe == io_state_in_1 ? 8'h83 : _GEN_1533; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _GEN_1535 = 8'hff == io_state_in_1 ? 8'h8d : _GEN_1534; // @[InvMixColumns.scala 127:{41,41}]
  wire [7:0] _tmp_state_1_T = _GEN_1279 ^ _GEN_1535; // @[InvMixColumns.scala 127:41]
  wire [7:0] _GEN_1537 = 8'h1 == io_state_in_2 ? 8'hb : 8'h0; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1538 = 8'h2 == io_state_in_2 ? 8'h16 : _GEN_1537; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1539 = 8'h3 == io_state_in_2 ? 8'h1d : _GEN_1538; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1540 = 8'h4 == io_state_in_2 ? 8'h2c : _GEN_1539; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1541 = 8'h5 == io_state_in_2 ? 8'h27 : _GEN_1540; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1542 = 8'h6 == io_state_in_2 ? 8'h3a : _GEN_1541; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1543 = 8'h7 == io_state_in_2 ? 8'h31 : _GEN_1542; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1544 = 8'h8 == io_state_in_2 ? 8'h58 : _GEN_1543; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1545 = 8'h9 == io_state_in_2 ? 8'h53 : _GEN_1544; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1546 = 8'ha == io_state_in_2 ? 8'h4e : _GEN_1545; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1547 = 8'hb == io_state_in_2 ? 8'h45 : _GEN_1546; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1548 = 8'hc == io_state_in_2 ? 8'h74 : _GEN_1547; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1549 = 8'hd == io_state_in_2 ? 8'h7f : _GEN_1548; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1550 = 8'he == io_state_in_2 ? 8'h62 : _GEN_1549; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1551 = 8'hf == io_state_in_2 ? 8'h69 : _GEN_1550; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1552 = 8'h10 == io_state_in_2 ? 8'hb0 : _GEN_1551; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1553 = 8'h11 == io_state_in_2 ? 8'hbb : _GEN_1552; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1554 = 8'h12 == io_state_in_2 ? 8'ha6 : _GEN_1553; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1555 = 8'h13 == io_state_in_2 ? 8'had : _GEN_1554; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1556 = 8'h14 == io_state_in_2 ? 8'h9c : _GEN_1555; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1557 = 8'h15 == io_state_in_2 ? 8'h97 : _GEN_1556; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1558 = 8'h16 == io_state_in_2 ? 8'h8a : _GEN_1557; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1559 = 8'h17 == io_state_in_2 ? 8'h81 : _GEN_1558; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1560 = 8'h18 == io_state_in_2 ? 8'he8 : _GEN_1559; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1561 = 8'h19 == io_state_in_2 ? 8'he3 : _GEN_1560; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1562 = 8'h1a == io_state_in_2 ? 8'hfe : _GEN_1561; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1563 = 8'h1b == io_state_in_2 ? 8'hf5 : _GEN_1562; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1564 = 8'h1c == io_state_in_2 ? 8'hc4 : _GEN_1563; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1565 = 8'h1d == io_state_in_2 ? 8'hcf : _GEN_1564; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1566 = 8'h1e == io_state_in_2 ? 8'hd2 : _GEN_1565; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1567 = 8'h1f == io_state_in_2 ? 8'hd9 : _GEN_1566; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1568 = 8'h20 == io_state_in_2 ? 8'h7b : _GEN_1567; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1569 = 8'h21 == io_state_in_2 ? 8'h70 : _GEN_1568; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1570 = 8'h22 == io_state_in_2 ? 8'h6d : _GEN_1569; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1571 = 8'h23 == io_state_in_2 ? 8'h66 : _GEN_1570; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1572 = 8'h24 == io_state_in_2 ? 8'h57 : _GEN_1571; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1573 = 8'h25 == io_state_in_2 ? 8'h5c : _GEN_1572; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1574 = 8'h26 == io_state_in_2 ? 8'h41 : _GEN_1573; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1575 = 8'h27 == io_state_in_2 ? 8'h4a : _GEN_1574; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1576 = 8'h28 == io_state_in_2 ? 8'h23 : _GEN_1575; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1577 = 8'h29 == io_state_in_2 ? 8'h28 : _GEN_1576; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1578 = 8'h2a == io_state_in_2 ? 8'h35 : _GEN_1577; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1579 = 8'h2b == io_state_in_2 ? 8'h3e : _GEN_1578; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1580 = 8'h2c == io_state_in_2 ? 8'hf : _GEN_1579; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1581 = 8'h2d == io_state_in_2 ? 8'h4 : _GEN_1580; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1582 = 8'h2e == io_state_in_2 ? 8'h19 : _GEN_1581; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1583 = 8'h2f == io_state_in_2 ? 8'h12 : _GEN_1582; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1584 = 8'h30 == io_state_in_2 ? 8'hcb : _GEN_1583; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1585 = 8'h31 == io_state_in_2 ? 8'hc0 : _GEN_1584; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1586 = 8'h32 == io_state_in_2 ? 8'hdd : _GEN_1585; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1587 = 8'h33 == io_state_in_2 ? 8'hd6 : _GEN_1586; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1588 = 8'h34 == io_state_in_2 ? 8'he7 : _GEN_1587; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1589 = 8'h35 == io_state_in_2 ? 8'hec : _GEN_1588; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1590 = 8'h36 == io_state_in_2 ? 8'hf1 : _GEN_1589; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1591 = 8'h37 == io_state_in_2 ? 8'hfa : _GEN_1590; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1592 = 8'h38 == io_state_in_2 ? 8'h93 : _GEN_1591; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1593 = 8'h39 == io_state_in_2 ? 8'h98 : _GEN_1592; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1594 = 8'h3a == io_state_in_2 ? 8'h85 : _GEN_1593; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1595 = 8'h3b == io_state_in_2 ? 8'h8e : _GEN_1594; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1596 = 8'h3c == io_state_in_2 ? 8'hbf : _GEN_1595; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1597 = 8'h3d == io_state_in_2 ? 8'hb4 : _GEN_1596; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1598 = 8'h3e == io_state_in_2 ? 8'ha9 : _GEN_1597; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1599 = 8'h3f == io_state_in_2 ? 8'ha2 : _GEN_1598; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1600 = 8'h40 == io_state_in_2 ? 8'hf6 : _GEN_1599; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1601 = 8'h41 == io_state_in_2 ? 8'hfd : _GEN_1600; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1602 = 8'h42 == io_state_in_2 ? 8'he0 : _GEN_1601; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1603 = 8'h43 == io_state_in_2 ? 8'heb : _GEN_1602; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1604 = 8'h44 == io_state_in_2 ? 8'hda : _GEN_1603; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1605 = 8'h45 == io_state_in_2 ? 8'hd1 : _GEN_1604; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1606 = 8'h46 == io_state_in_2 ? 8'hcc : _GEN_1605; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1607 = 8'h47 == io_state_in_2 ? 8'hc7 : _GEN_1606; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1608 = 8'h48 == io_state_in_2 ? 8'hae : _GEN_1607; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1609 = 8'h49 == io_state_in_2 ? 8'ha5 : _GEN_1608; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1610 = 8'h4a == io_state_in_2 ? 8'hb8 : _GEN_1609; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1611 = 8'h4b == io_state_in_2 ? 8'hb3 : _GEN_1610; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1612 = 8'h4c == io_state_in_2 ? 8'h82 : _GEN_1611; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1613 = 8'h4d == io_state_in_2 ? 8'h89 : _GEN_1612; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1614 = 8'h4e == io_state_in_2 ? 8'h94 : _GEN_1613; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1615 = 8'h4f == io_state_in_2 ? 8'h9f : _GEN_1614; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1616 = 8'h50 == io_state_in_2 ? 8'h46 : _GEN_1615; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1617 = 8'h51 == io_state_in_2 ? 8'h4d : _GEN_1616; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1618 = 8'h52 == io_state_in_2 ? 8'h50 : _GEN_1617; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1619 = 8'h53 == io_state_in_2 ? 8'h5b : _GEN_1618; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1620 = 8'h54 == io_state_in_2 ? 8'h6a : _GEN_1619; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1621 = 8'h55 == io_state_in_2 ? 8'h61 : _GEN_1620; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1622 = 8'h56 == io_state_in_2 ? 8'h7c : _GEN_1621; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1623 = 8'h57 == io_state_in_2 ? 8'h77 : _GEN_1622; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1624 = 8'h58 == io_state_in_2 ? 8'h1e : _GEN_1623; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1625 = 8'h59 == io_state_in_2 ? 8'h15 : _GEN_1624; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1626 = 8'h5a == io_state_in_2 ? 8'h8 : _GEN_1625; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1627 = 8'h5b == io_state_in_2 ? 8'h3 : _GEN_1626; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1628 = 8'h5c == io_state_in_2 ? 8'h32 : _GEN_1627; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1629 = 8'h5d == io_state_in_2 ? 8'h39 : _GEN_1628; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1630 = 8'h5e == io_state_in_2 ? 8'h24 : _GEN_1629; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1631 = 8'h5f == io_state_in_2 ? 8'h2f : _GEN_1630; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1632 = 8'h60 == io_state_in_2 ? 8'h8d : _GEN_1631; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1633 = 8'h61 == io_state_in_2 ? 8'h86 : _GEN_1632; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1634 = 8'h62 == io_state_in_2 ? 8'h9b : _GEN_1633; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1635 = 8'h63 == io_state_in_2 ? 8'h90 : _GEN_1634; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1636 = 8'h64 == io_state_in_2 ? 8'ha1 : _GEN_1635; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1637 = 8'h65 == io_state_in_2 ? 8'haa : _GEN_1636; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1638 = 8'h66 == io_state_in_2 ? 8'hb7 : _GEN_1637; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1639 = 8'h67 == io_state_in_2 ? 8'hbc : _GEN_1638; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1640 = 8'h68 == io_state_in_2 ? 8'hd5 : _GEN_1639; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1641 = 8'h69 == io_state_in_2 ? 8'hde : _GEN_1640; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1642 = 8'h6a == io_state_in_2 ? 8'hc3 : _GEN_1641; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1643 = 8'h6b == io_state_in_2 ? 8'hc8 : _GEN_1642; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1644 = 8'h6c == io_state_in_2 ? 8'hf9 : _GEN_1643; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1645 = 8'h6d == io_state_in_2 ? 8'hf2 : _GEN_1644; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1646 = 8'h6e == io_state_in_2 ? 8'hef : _GEN_1645; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1647 = 8'h6f == io_state_in_2 ? 8'he4 : _GEN_1646; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1648 = 8'h70 == io_state_in_2 ? 8'h3d : _GEN_1647; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1649 = 8'h71 == io_state_in_2 ? 8'h36 : _GEN_1648; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1650 = 8'h72 == io_state_in_2 ? 8'h2b : _GEN_1649; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1651 = 8'h73 == io_state_in_2 ? 8'h20 : _GEN_1650; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1652 = 8'h74 == io_state_in_2 ? 8'h11 : _GEN_1651; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1653 = 8'h75 == io_state_in_2 ? 8'h1a : _GEN_1652; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1654 = 8'h76 == io_state_in_2 ? 8'h7 : _GEN_1653; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1655 = 8'h77 == io_state_in_2 ? 8'hc : _GEN_1654; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1656 = 8'h78 == io_state_in_2 ? 8'h65 : _GEN_1655; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1657 = 8'h79 == io_state_in_2 ? 8'h6e : _GEN_1656; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1658 = 8'h7a == io_state_in_2 ? 8'h73 : _GEN_1657; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1659 = 8'h7b == io_state_in_2 ? 8'h78 : _GEN_1658; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1660 = 8'h7c == io_state_in_2 ? 8'h49 : _GEN_1659; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1661 = 8'h7d == io_state_in_2 ? 8'h42 : _GEN_1660; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1662 = 8'h7e == io_state_in_2 ? 8'h5f : _GEN_1661; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1663 = 8'h7f == io_state_in_2 ? 8'h54 : _GEN_1662; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1664 = 8'h80 == io_state_in_2 ? 8'hf7 : _GEN_1663; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1665 = 8'h81 == io_state_in_2 ? 8'hfc : _GEN_1664; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1666 = 8'h82 == io_state_in_2 ? 8'he1 : _GEN_1665; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1667 = 8'h83 == io_state_in_2 ? 8'hea : _GEN_1666; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1668 = 8'h84 == io_state_in_2 ? 8'hdb : _GEN_1667; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1669 = 8'h85 == io_state_in_2 ? 8'hd0 : _GEN_1668; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1670 = 8'h86 == io_state_in_2 ? 8'hcd : _GEN_1669; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1671 = 8'h87 == io_state_in_2 ? 8'hc6 : _GEN_1670; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1672 = 8'h88 == io_state_in_2 ? 8'haf : _GEN_1671; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1673 = 8'h89 == io_state_in_2 ? 8'ha4 : _GEN_1672; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1674 = 8'h8a == io_state_in_2 ? 8'hb9 : _GEN_1673; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1675 = 8'h8b == io_state_in_2 ? 8'hb2 : _GEN_1674; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1676 = 8'h8c == io_state_in_2 ? 8'h83 : _GEN_1675; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1677 = 8'h8d == io_state_in_2 ? 8'h88 : _GEN_1676; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1678 = 8'h8e == io_state_in_2 ? 8'h95 : _GEN_1677; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1679 = 8'h8f == io_state_in_2 ? 8'h9e : _GEN_1678; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1680 = 8'h90 == io_state_in_2 ? 8'h47 : _GEN_1679; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1681 = 8'h91 == io_state_in_2 ? 8'h4c : _GEN_1680; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1682 = 8'h92 == io_state_in_2 ? 8'h51 : _GEN_1681; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1683 = 8'h93 == io_state_in_2 ? 8'h5a : _GEN_1682; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1684 = 8'h94 == io_state_in_2 ? 8'h6b : _GEN_1683; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1685 = 8'h95 == io_state_in_2 ? 8'h60 : _GEN_1684; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1686 = 8'h96 == io_state_in_2 ? 8'h7d : _GEN_1685; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1687 = 8'h97 == io_state_in_2 ? 8'h76 : _GEN_1686; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1688 = 8'h98 == io_state_in_2 ? 8'h1f : _GEN_1687; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1689 = 8'h99 == io_state_in_2 ? 8'h14 : _GEN_1688; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1690 = 8'h9a == io_state_in_2 ? 8'h9 : _GEN_1689; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1691 = 8'h9b == io_state_in_2 ? 8'h2 : _GEN_1690; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1692 = 8'h9c == io_state_in_2 ? 8'h33 : _GEN_1691; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1693 = 8'h9d == io_state_in_2 ? 8'h38 : _GEN_1692; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1694 = 8'h9e == io_state_in_2 ? 8'h25 : _GEN_1693; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1695 = 8'h9f == io_state_in_2 ? 8'h2e : _GEN_1694; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1696 = 8'ha0 == io_state_in_2 ? 8'h8c : _GEN_1695; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1697 = 8'ha1 == io_state_in_2 ? 8'h87 : _GEN_1696; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1698 = 8'ha2 == io_state_in_2 ? 8'h9a : _GEN_1697; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1699 = 8'ha3 == io_state_in_2 ? 8'h91 : _GEN_1698; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1700 = 8'ha4 == io_state_in_2 ? 8'ha0 : _GEN_1699; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1701 = 8'ha5 == io_state_in_2 ? 8'hab : _GEN_1700; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1702 = 8'ha6 == io_state_in_2 ? 8'hb6 : _GEN_1701; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1703 = 8'ha7 == io_state_in_2 ? 8'hbd : _GEN_1702; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1704 = 8'ha8 == io_state_in_2 ? 8'hd4 : _GEN_1703; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1705 = 8'ha9 == io_state_in_2 ? 8'hdf : _GEN_1704; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1706 = 8'haa == io_state_in_2 ? 8'hc2 : _GEN_1705; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1707 = 8'hab == io_state_in_2 ? 8'hc9 : _GEN_1706; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1708 = 8'hac == io_state_in_2 ? 8'hf8 : _GEN_1707; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1709 = 8'had == io_state_in_2 ? 8'hf3 : _GEN_1708; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1710 = 8'hae == io_state_in_2 ? 8'hee : _GEN_1709; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1711 = 8'haf == io_state_in_2 ? 8'he5 : _GEN_1710; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1712 = 8'hb0 == io_state_in_2 ? 8'h3c : _GEN_1711; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1713 = 8'hb1 == io_state_in_2 ? 8'h37 : _GEN_1712; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1714 = 8'hb2 == io_state_in_2 ? 8'h2a : _GEN_1713; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1715 = 8'hb3 == io_state_in_2 ? 8'h21 : _GEN_1714; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1716 = 8'hb4 == io_state_in_2 ? 8'h10 : _GEN_1715; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1717 = 8'hb5 == io_state_in_2 ? 8'h1b : _GEN_1716; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1718 = 8'hb6 == io_state_in_2 ? 8'h6 : _GEN_1717; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1719 = 8'hb7 == io_state_in_2 ? 8'hd : _GEN_1718; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1720 = 8'hb8 == io_state_in_2 ? 8'h64 : _GEN_1719; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1721 = 8'hb9 == io_state_in_2 ? 8'h6f : _GEN_1720; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1722 = 8'hba == io_state_in_2 ? 8'h72 : _GEN_1721; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1723 = 8'hbb == io_state_in_2 ? 8'h79 : _GEN_1722; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1724 = 8'hbc == io_state_in_2 ? 8'h48 : _GEN_1723; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1725 = 8'hbd == io_state_in_2 ? 8'h43 : _GEN_1724; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1726 = 8'hbe == io_state_in_2 ? 8'h5e : _GEN_1725; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1727 = 8'hbf == io_state_in_2 ? 8'h55 : _GEN_1726; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1728 = 8'hc0 == io_state_in_2 ? 8'h1 : _GEN_1727; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1729 = 8'hc1 == io_state_in_2 ? 8'ha : _GEN_1728; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1730 = 8'hc2 == io_state_in_2 ? 8'h17 : _GEN_1729; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1731 = 8'hc3 == io_state_in_2 ? 8'h1c : _GEN_1730; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1732 = 8'hc4 == io_state_in_2 ? 8'h2d : _GEN_1731; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1733 = 8'hc5 == io_state_in_2 ? 8'h26 : _GEN_1732; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1734 = 8'hc6 == io_state_in_2 ? 8'h3b : _GEN_1733; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1735 = 8'hc7 == io_state_in_2 ? 8'h30 : _GEN_1734; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1736 = 8'hc8 == io_state_in_2 ? 8'h59 : _GEN_1735; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1737 = 8'hc9 == io_state_in_2 ? 8'h52 : _GEN_1736; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1738 = 8'hca == io_state_in_2 ? 8'h4f : _GEN_1737; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1739 = 8'hcb == io_state_in_2 ? 8'h44 : _GEN_1738; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1740 = 8'hcc == io_state_in_2 ? 8'h75 : _GEN_1739; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1741 = 8'hcd == io_state_in_2 ? 8'h7e : _GEN_1740; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1742 = 8'hce == io_state_in_2 ? 8'h63 : _GEN_1741; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1743 = 8'hcf == io_state_in_2 ? 8'h68 : _GEN_1742; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1744 = 8'hd0 == io_state_in_2 ? 8'hb1 : _GEN_1743; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1745 = 8'hd1 == io_state_in_2 ? 8'hba : _GEN_1744; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1746 = 8'hd2 == io_state_in_2 ? 8'ha7 : _GEN_1745; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1747 = 8'hd3 == io_state_in_2 ? 8'hac : _GEN_1746; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1748 = 8'hd4 == io_state_in_2 ? 8'h9d : _GEN_1747; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1749 = 8'hd5 == io_state_in_2 ? 8'h96 : _GEN_1748; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1750 = 8'hd6 == io_state_in_2 ? 8'h8b : _GEN_1749; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1751 = 8'hd7 == io_state_in_2 ? 8'h80 : _GEN_1750; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1752 = 8'hd8 == io_state_in_2 ? 8'he9 : _GEN_1751; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1753 = 8'hd9 == io_state_in_2 ? 8'he2 : _GEN_1752; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1754 = 8'hda == io_state_in_2 ? 8'hff : _GEN_1753; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1755 = 8'hdb == io_state_in_2 ? 8'hf4 : _GEN_1754; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1756 = 8'hdc == io_state_in_2 ? 8'hc5 : _GEN_1755; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1757 = 8'hdd == io_state_in_2 ? 8'hce : _GEN_1756; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1758 = 8'hde == io_state_in_2 ? 8'hd3 : _GEN_1757; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1759 = 8'hdf == io_state_in_2 ? 8'hd8 : _GEN_1758; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1760 = 8'he0 == io_state_in_2 ? 8'h7a : _GEN_1759; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1761 = 8'he1 == io_state_in_2 ? 8'h71 : _GEN_1760; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1762 = 8'he2 == io_state_in_2 ? 8'h6c : _GEN_1761; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1763 = 8'he3 == io_state_in_2 ? 8'h67 : _GEN_1762; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1764 = 8'he4 == io_state_in_2 ? 8'h56 : _GEN_1763; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1765 = 8'he5 == io_state_in_2 ? 8'h5d : _GEN_1764; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1766 = 8'he6 == io_state_in_2 ? 8'h40 : _GEN_1765; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1767 = 8'he7 == io_state_in_2 ? 8'h4b : _GEN_1766; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1768 = 8'he8 == io_state_in_2 ? 8'h22 : _GEN_1767; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1769 = 8'he9 == io_state_in_2 ? 8'h29 : _GEN_1768; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1770 = 8'hea == io_state_in_2 ? 8'h34 : _GEN_1769; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1771 = 8'heb == io_state_in_2 ? 8'h3f : _GEN_1770; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1772 = 8'hec == io_state_in_2 ? 8'he : _GEN_1771; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1773 = 8'hed == io_state_in_2 ? 8'h5 : _GEN_1772; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1774 = 8'hee == io_state_in_2 ? 8'h18 : _GEN_1773; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1775 = 8'hef == io_state_in_2 ? 8'h13 : _GEN_1774; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1776 = 8'hf0 == io_state_in_2 ? 8'hca : _GEN_1775; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1777 = 8'hf1 == io_state_in_2 ? 8'hc1 : _GEN_1776; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1778 = 8'hf2 == io_state_in_2 ? 8'hdc : _GEN_1777; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1779 = 8'hf3 == io_state_in_2 ? 8'hd7 : _GEN_1778; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1780 = 8'hf4 == io_state_in_2 ? 8'he6 : _GEN_1779; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1781 = 8'hf5 == io_state_in_2 ? 8'hed : _GEN_1780; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1782 = 8'hf6 == io_state_in_2 ? 8'hf0 : _GEN_1781; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1783 = 8'hf7 == io_state_in_2 ? 8'hfb : _GEN_1782; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1784 = 8'hf8 == io_state_in_2 ? 8'h92 : _GEN_1783; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1785 = 8'hf9 == io_state_in_2 ? 8'h99 : _GEN_1784; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1786 = 8'hfa == io_state_in_2 ? 8'h84 : _GEN_1785; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1787 = 8'hfb == io_state_in_2 ? 8'h8f : _GEN_1786; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1788 = 8'hfc == io_state_in_2 ? 8'hbe : _GEN_1787; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1789 = 8'hfd == io_state_in_2 ? 8'hb5 : _GEN_1788; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1790 = 8'hfe == io_state_in_2 ? 8'ha8 : _GEN_1789; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _GEN_1791 = 8'hff == io_state_in_2 ? 8'ha3 : _GEN_1790; // @[InvMixColumns.scala 127:{65,65}]
  wire [7:0] _tmp_state_1_T_1 = _tmp_state_1_T ^ _GEN_1791; // @[InvMixColumns.scala 127:65]
  wire [7:0] _GEN_1793 = 8'h1 == io_state_in_3 ? 8'hd : 8'h0; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1794 = 8'h2 == io_state_in_3 ? 8'h1a : _GEN_1793; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1795 = 8'h3 == io_state_in_3 ? 8'h17 : _GEN_1794; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1796 = 8'h4 == io_state_in_3 ? 8'h34 : _GEN_1795; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1797 = 8'h5 == io_state_in_3 ? 8'h39 : _GEN_1796; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1798 = 8'h6 == io_state_in_3 ? 8'h2e : _GEN_1797; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1799 = 8'h7 == io_state_in_3 ? 8'h23 : _GEN_1798; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1800 = 8'h8 == io_state_in_3 ? 8'h68 : _GEN_1799; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1801 = 8'h9 == io_state_in_3 ? 8'h65 : _GEN_1800; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1802 = 8'ha == io_state_in_3 ? 8'h72 : _GEN_1801; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1803 = 8'hb == io_state_in_3 ? 8'h7f : _GEN_1802; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1804 = 8'hc == io_state_in_3 ? 8'h5c : _GEN_1803; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1805 = 8'hd == io_state_in_3 ? 8'h51 : _GEN_1804; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1806 = 8'he == io_state_in_3 ? 8'h46 : _GEN_1805; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1807 = 8'hf == io_state_in_3 ? 8'h4b : _GEN_1806; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1808 = 8'h10 == io_state_in_3 ? 8'hd0 : _GEN_1807; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1809 = 8'h11 == io_state_in_3 ? 8'hdd : _GEN_1808; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1810 = 8'h12 == io_state_in_3 ? 8'hca : _GEN_1809; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1811 = 8'h13 == io_state_in_3 ? 8'hc7 : _GEN_1810; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1812 = 8'h14 == io_state_in_3 ? 8'he4 : _GEN_1811; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1813 = 8'h15 == io_state_in_3 ? 8'he9 : _GEN_1812; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1814 = 8'h16 == io_state_in_3 ? 8'hfe : _GEN_1813; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1815 = 8'h17 == io_state_in_3 ? 8'hf3 : _GEN_1814; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1816 = 8'h18 == io_state_in_3 ? 8'hb8 : _GEN_1815; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1817 = 8'h19 == io_state_in_3 ? 8'hb5 : _GEN_1816; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1818 = 8'h1a == io_state_in_3 ? 8'ha2 : _GEN_1817; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1819 = 8'h1b == io_state_in_3 ? 8'haf : _GEN_1818; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1820 = 8'h1c == io_state_in_3 ? 8'h8c : _GEN_1819; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1821 = 8'h1d == io_state_in_3 ? 8'h81 : _GEN_1820; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1822 = 8'h1e == io_state_in_3 ? 8'h96 : _GEN_1821; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1823 = 8'h1f == io_state_in_3 ? 8'h9b : _GEN_1822; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1824 = 8'h20 == io_state_in_3 ? 8'hbb : _GEN_1823; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1825 = 8'h21 == io_state_in_3 ? 8'hb6 : _GEN_1824; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1826 = 8'h22 == io_state_in_3 ? 8'ha1 : _GEN_1825; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1827 = 8'h23 == io_state_in_3 ? 8'hac : _GEN_1826; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1828 = 8'h24 == io_state_in_3 ? 8'h8f : _GEN_1827; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1829 = 8'h25 == io_state_in_3 ? 8'h82 : _GEN_1828; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1830 = 8'h26 == io_state_in_3 ? 8'h95 : _GEN_1829; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1831 = 8'h27 == io_state_in_3 ? 8'h98 : _GEN_1830; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1832 = 8'h28 == io_state_in_3 ? 8'hd3 : _GEN_1831; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1833 = 8'h29 == io_state_in_3 ? 8'hde : _GEN_1832; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1834 = 8'h2a == io_state_in_3 ? 8'hc9 : _GEN_1833; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1835 = 8'h2b == io_state_in_3 ? 8'hc4 : _GEN_1834; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1836 = 8'h2c == io_state_in_3 ? 8'he7 : _GEN_1835; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1837 = 8'h2d == io_state_in_3 ? 8'hea : _GEN_1836; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1838 = 8'h2e == io_state_in_3 ? 8'hfd : _GEN_1837; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1839 = 8'h2f == io_state_in_3 ? 8'hf0 : _GEN_1838; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1840 = 8'h30 == io_state_in_3 ? 8'h6b : _GEN_1839; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1841 = 8'h31 == io_state_in_3 ? 8'h66 : _GEN_1840; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1842 = 8'h32 == io_state_in_3 ? 8'h71 : _GEN_1841; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1843 = 8'h33 == io_state_in_3 ? 8'h7c : _GEN_1842; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1844 = 8'h34 == io_state_in_3 ? 8'h5f : _GEN_1843; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1845 = 8'h35 == io_state_in_3 ? 8'h52 : _GEN_1844; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1846 = 8'h36 == io_state_in_3 ? 8'h45 : _GEN_1845; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1847 = 8'h37 == io_state_in_3 ? 8'h48 : _GEN_1846; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1848 = 8'h38 == io_state_in_3 ? 8'h3 : _GEN_1847; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1849 = 8'h39 == io_state_in_3 ? 8'he : _GEN_1848; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1850 = 8'h3a == io_state_in_3 ? 8'h19 : _GEN_1849; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1851 = 8'h3b == io_state_in_3 ? 8'h14 : _GEN_1850; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1852 = 8'h3c == io_state_in_3 ? 8'h37 : _GEN_1851; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1853 = 8'h3d == io_state_in_3 ? 8'h3a : _GEN_1852; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1854 = 8'h3e == io_state_in_3 ? 8'h2d : _GEN_1853; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1855 = 8'h3f == io_state_in_3 ? 8'h20 : _GEN_1854; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1856 = 8'h40 == io_state_in_3 ? 8'h6d : _GEN_1855; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1857 = 8'h41 == io_state_in_3 ? 8'h60 : _GEN_1856; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1858 = 8'h42 == io_state_in_3 ? 8'h77 : _GEN_1857; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1859 = 8'h43 == io_state_in_3 ? 8'h7a : _GEN_1858; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1860 = 8'h44 == io_state_in_3 ? 8'h59 : _GEN_1859; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1861 = 8'h45 == io_state_in_3 ? 8'h54 : _GEN_1860; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1862 = 8'h46 == io_state_in_3 ? 8'h43 : _GEN_1861; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1863 = 8'h47 == io_state_in_3 ? 8'h4e : _GEN_1862; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1864 = 8'h48 == io_state_in_3 ? 8'h5 : _GEN_1863; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1865 = 8'h49 == io_state_in_3 ? 8'h8 : _GEN_1864; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1866 = 8'h4a == io_state_in_3 ? 8'h1f : _GEN_1865; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1867 = 8'h4b == io_state_in_3 ? 8'h12 : _GEN_1866; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1868 = 8'h4c == io_state_in_3 ? 8'h31 : _GEN_1867; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1869 = 8'h4d == io_state_in_3 ? 8'h3c : _GEN_1868; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1870 = 8'h4e == io_state_in_3 ? 8'h2b : _GEN_1869; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1871 = 8'h4f == io_state_in_3 ? 8'h26 : _GEN_1870; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1872 = 8'h50 == io_state_in_3 ? 8'hbd : _GEN_1871; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1873 = 8'h51 == io_state_in_3 ? 8'hb0 : _GEN_1872; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1874 = 8'h52 == io_state_in_3 ? 8'ha7 : _GEN_1873; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1875 = 8'h53 == io_state_in_3 ? 8'haa : _GEN_1874; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1876 = 8'h54 == io_state_in_3 ? 8'h89 : _GEN_1875; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1877 = 8'h55 == io_state_in_3 ? 8'h84 : _GEN_1876; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1878 = 8'h56 == io_state_in_3 ? 8'h93 : _GEN_1877; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1879 = 8'h57 == io_state_in_3 ? 8'h9e : _GEN_1878; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1880 = 8'h58 == io_state_in_3 ? 8'hd5 : _GEN_1879; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1881 = 8'h59 == io_state_in_3 ? 8'hd8 : _GEN_1880; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1882 = 8'h5a == io_state_in_3 ? 8'hcf : _GEN_1881; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1883 = 8'h5b == io_state_in_3 ? 8'hc2 : _GEN_1882; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1884 = 8'h5c == io_state_in_3 ? 8'he1 : _GEN_1883; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1885 = 8'h5d == io_state_in_3 ? 8'hec : _GEN_1884; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1886 = 8'h5e == io_state_in_3 ? 8'hfb : _GEN_1885; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1887 = 8'h5f == io_state_in_3 ? 8'hf6 : _GEN_1886; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1888 = 8'h60 == io_state_in_3 ? 8'hd6 : _GEN_1887; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1889 = 8'h61 == io_state_in_3 ? 8'hdb : _GEN_1888; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1890 = 8'h62 == io_state_in_3 ? 8'hcc : _GEN_1889; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1891 = 8'h63 == io_state_in_3 ? 8'hc1 : _GEN_1890; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1892 = 8'h64 == io_state_in_3 ? 8'he2 : _GEN_1891; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1893 = 8'h65 == io_state_in_3 ? 8'hef : _GEN_1892; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1894 = 8'h66 == io_state_in_3 ? 8'hf8 : _GEN_1893; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1895 = 8'h67 == io_state_in_3 ? 8'hf5 : _GEN_1894; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1896 = 8'h68 == io_state_in_3 ? 8'hbe : _GEN_1895; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1897 = 8'h69 == io_state_in_3 ? 8'hb3 : _GEN_1896; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1898 = 8'h6a == io_state_in_3 ? 8'ha4 : _GEN_1897; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1899 = 8'h6b == io_state_in_3 ? 8'ha9 : _GEN_1898; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1900 = 8'h6c == io_state_in_3 ? 8'h8a : _GEN_1899; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1901 = 8'h6d == io_state_in_3 ? 8'h87 : _GEN_1900; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1902 = 8'h6e == io_state_in_3 ? 8'h90 : _GEN_1901; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1903 = 8'h6f == io_state_in_3 ? 8'h9d : _GEN_1902; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1904 = 8'h70 == io_state_in_3 ? 8'h6 : _GEN_1903; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1905 = 8'h71 == io_state_in_3 ? 8'hb : _GEN_1904; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1906 = 8'h72 == io_state_in_3 ? 8'h1c : _GEN_1905; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1907 = 8'h73 == io_state_in_3 ? 8'h11 : _GEN_1906; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1908 = 8'h74 == io_state_in_3 ? 8'h32 : _GEN_1907; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1909 = 8'h75 == io_state_in_3 ? 8'h3f : _GEN_1908; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1910 = 8'h76 == io_state_in_3 ? 8'h28 : _GEN_1909; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1911 = 8'h77 == io_state_in_3 ? 8'h25 : _GEN_1910; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1912 = 8'h78 == io_state_in_3 ? 8'h6e : _GEN_1911; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1913 = 8'h79 == io_state_in_3 ? 8'h63 : _GEN_1912; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1914 = 8'h7a == io_state_in_3 ? 8'h74 : _GEN_1913; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1915 = 8'h7b == io_state_in_3 ? 8'h79 : _GEN_1914; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1916 = 8'h7c == io_state_in_3 ? 8'h5a : _GEN_1915; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1917 = 8'h7d == io_state_in_3 ? 8'h57 : _GEN_1916; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1918 = 8'h7e == io_state_in_3 ? 8'h40 : _GEN_1917; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1919 = 8'h7f == io_state_in_3 ? 8'h4d : _GEN_1918; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1920 = 8'h80 == io_state_in_3 ? 8'hda : _GEN_1919; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1921 = 8'h81 == io_state_in_3 ? 8'hd7 : _GEN_1920; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1922 = 8'h82 == io_state_in_3 ? 8'hc0 : _GEN_1921; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1923 = 8'h83 == io_state_in_3 ? 8'hcd : _GEN_1922; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1924 = 8'h84 == io_state_in_3 ? 8'hee : _GEN_1923; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1925 = 8'h85 == io_state_in_3 ? 8'he3 : _GEN_1924; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1926 = 8'h86 == io_state_in_3 ? 8'hf4 : _GEN_1925; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1927 = 8'h87 == io_state_in_3 ? 8'hf9 : _GEN_1926; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1928 = 8'h88 == io_state_in_3 ? 8'hb2 : _GEN_1927; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1929 = 8'h89 == io_state_in_3 ? 8'hbf : _GEN_1928; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1930 = 8'h8a == io_state_in_3 ? 8'ha8 : _GEN_1929; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1931 = 8'h8b == io_state_in_3 ? 8'ha5 : _GEN_1930; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1932 = 8'h8c == io_state_in_3 ? 8'h86 : _GEN_1931; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1933 = 8'h8d == io_state_in_3 ? 8'h8b : _GEN_1932; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1934 = 8'h8e == io_state_in_3 ? 8'h9c : _GEN_1933; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1935 = 8'h8f == io_state_in_3 ? 8'h91 : _GEN_1934; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1936 = 8'h90 == io_state_in_3 ? 8'ha : _GEN_1935; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1937 = 8'h91 == io_state_in_3 ? 8'h7 : _GEN_1936; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1938 = 8'h92 == io_state_in_3 ? 8'h10 : _GEN_1937; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1939 = 8'h93 == io_state_in_3 ? 8'h1d : _GEN_1938; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1940 = 8'h94 == io_state_in_3 ? 8'h3e : _GEN_1939; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1941 = 8'h95 == io_state_in_3 ? 8'h33 : _GEN_1940; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1942 = 8'h96 == io_state_in_3 ? 8'h24 : _GEN_1941; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1943 = 8'h97 == io_state_in_3 ? 8'h29 : _GEN_1942; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1944 = 8'h98 == io_state_in_3 ? 8'h62 : _GEN_1943; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1945 = 8'h99 == io_state_in_3 ? 8'h6f : _GEN_1944; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1946 = 8'h9a == io_state_in_3 ? 8'h78 : _GEN_1945; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1947 = 8'h9b == io_state_in_3 ? 8'h75 : _GEN_1946; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1948 = 8'h9c == io_state_in_3 ? 8'h56 : _GEN_1947; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1949 = 8'h9d == io_state_in_3 ? 8'h5b : _GEN_1948; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1950 = 8'h9e == io_state_in_3 ? 8'h4c : _GEN_1949; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1951 = 8'h9f == io_state_in_3 ? 8'h41 : _GEN_1950; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1952 = 8'ha0 == io_state_in_3 ? 8'h61 : _GEN_1951; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1953 = 8'ha1 == io_state_in_3 ? 8'h6c : _GEN_1952; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1954 = 8'ha2 == io_state_in_3 ? 8'h7b : _GEN_1953; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1955 = 8'ha3 == io_state_in_3 ? 8'h76 : _GEN_1954; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1956 = 8'ha4 == io_state_in_3 ? 8'h55 : _GEN_1955; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1957 = 8'ha5 == io_state_in_3 ? 8'h58 : _GEN_1956; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1958 = 8'ha6 == io_state_in_3 ? 8'h4f : _GEN_1957; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1959 = 8'ha7 == io_state_in_3 ? 8'h42 : _GEN_1958; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1960 = 8'ha8 == io_state_in_3 ? 8'h9 : _GEN_1959; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1961 = 8'ha9 == io_state_in_3 ? 8'h4 : _GEN_1960; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1962 = 8'haa == io_state_in_3 ? 8'h13 : _GEN_1961; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1963 = 8'hab == io_state_in_3 ? 8'h1e : _GEN_1962; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1964 = 8'hac == io_state_in_3 ? 8'h3d : _GEN_1963; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1965 = 8'had == io_state_in_3 ? 8'h30 : _GEN_1964; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1966 = 8'hae == io_state_in_3 ? 8'h27 : _GEN_1965; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1967 = 8'haf == io_state_in_3 ? 8'h2a : _GEN_1966; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1968 = 8'hb0 == io_state_in_3 ? 8'hb1 : _GEN_1967; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1969 = 8'hb1 == io_state_in_3 ? 8'hbc : _GEN_1968; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1970 = 8'hb2 == io_state_in_3 ? 8'hab : _GEN_1969; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1971 = 8'hb3 == io_state_in_3 ? 8'ha6 : _GEN_1970; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1972 = 8'hb4 == io_state_in_3 ? 8'h85 : _GEN_1971; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1973 = 8'hb5 == io_state_in_3 ? 8'h88 : _GEN_1972; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1974 = 8'hb6 == io_state_in_3 ? 8'h9f : _GEN_1973; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1975 = 8'hb7 == io_state_in_3 ? 8'h92 : _GEN_1974; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1976 = 8'hb8 == io_state_in_3 ? 8'hd9 : _GEN_1975; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1977 = 8'hb9 == io_state_in_3 ? 8'hd4 : _GEN_1976; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1978 = 8'hba == io_state_in_3 ? 8'hc3 : _GEN_1977; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1979 = 8'hbb == io_state_in_3 ? 8'hce : _GEN_1978; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1980 = 8'hbc == io_state_in_3 ? 8'hed : _GEN_1979; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1981 = 8'hbd == io_state_in_3 ? 8'he0 : _GEN_1980; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1982 = 8'hbe == io_state_in_3 ? 8'hf7 : _GEN_1981; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1983 = 8'hbf == io_state_in_3 ? 8'hfa : _GEN_1982; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1984 = 8'hc0 == io_state_in_3 ? 8'hb7 : _GEN_1983; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1985 = 8'hc1 == io_state_in_3 ? 8'hba : _GEN_1984; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1986 = 8'hc2 == io_state_in_3 ? 8'had : _GEN_1985; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1987 = 8'hc3 == io_state_in_3 ? 8'ha0 : _GEN_1986; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1988 = 8'hc4 == io_state_in_3 ? 8'h83 : _GEN_1987; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1989 = 8'hc5 == io_state_in_3 ? 8'h8e : _GEN_1988; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1990 = 8'hc6 == io_state_in_3 ? 8'h99 : _GEN_1989; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1991 = 8'hc7 == io_state_in_3 ? 8'h94 : _GEN_1990; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1992 = 8'hc8 == io_state_in_3 ? 8'hdf : _GEN_1991; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1993 = 8'hc9 == io_state_in_3 ? 8'hd2 : _GEN_1992; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1994 = 8'hca == io_state_in_3 ? 8'hc5 : _GEN_1993; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1995 = 8'hcb == io_state_in_3 ? 8'hc8 : _GEN_1994; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1996 = 8'hcc == io_state_in_3 ? 8'heb : _GEN_1995; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1997 = 8'hcd == io_state_in_3 ? 8'he6 : _GEN_1996; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1998 = 8'hce == io_state_in_3 ? 8'hf1 : _GEN_1997; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_1999 = 8'hcf == io_state_in_3 ? 8'hfc : _GEN_1998; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2000 = 8'hd0 == io_state_in_3 ? 8'h67 : _GEN_1999; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2001 = 8'hd1 == io_state_in_3 ? 8'h6a : _GEN_2000; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2002 = 8'hd2 == io_state_in_3 ? 8'h7d : _GEN_2001; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2003 = 8'hd3 == io_state_in_3 ? 8'h70 : _GEN_2002; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2004 = 8'hd4 == io_state_in_3 ? 8'h53 : _GEN_2003; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2005 = 8'hd5 == io_state_in_3 ? 8'h5e : _GEN_2004; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2006 = 8'hd6 == io_state_in_3 ? 8'h49 : _GEN_2005; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2007 = 8'hd7 == io_state_in_3 ? 8'h44 : _GEN_2006; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2008 = 8'hd8 == io_state_in_3 ? 8'hf : _GEN_2007; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2009 = 8'hd9 == io_state_in_3 ? 8'h2 : _GEN_2008; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2010 = 8'hda == io_state_in_3 ? 8'h15 : _GEN_2009; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2011 = 8'hdb == io_state_in_3 ? 8'h18 : _GEN_2010; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2012 = 8'hdc == io_state_in_3 ? 8'h3b : _GEN_2011; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2013 = 8'hdd == io_state_in_3 ? 8'h36 : _GEN_2012; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2014 = 8'hde == io_state_in_3 ? 8'h21 : _GEN_2013; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2015 = 8'hdf == io_state_in_3 ? 8'h2c : _GEN_2014; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2016 = 8'he0 == io_state_in_3 ? 8'hc : _GEN_2015; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2017 = 8'he1 == io_state_in_3 ? 8'h1 : _GEN_2016; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2018 = 8'he2 == io_state_in_3 ? 8'h16 : _GEN_2017; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2019 = 8'he3 == io_state_in_3 ? 8'h1b : _GEN_2018; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2020 = 8'he4 == io_state_in_3 ? 8'h38 : _GEN_2019; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2021 = 8'he5 == io_state_in_3 ? 8'h35 : _GEN_2020; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2022 = 8'he6 == io_state_in_3 ? 8'h22 : _GEN_2021; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2023 = 8'he7 == io_state_in_3 ? 8'h2f : _GEN_2022; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2024 = 8'he8 == io_state_in_3 ? 8'h64 : _GEN_2023; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2025 = 8'he9 == io_state_in_3 ? 8'h69 : _GEN_2024; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2026 = 8'hea == io_state_in_3 ? 8'h7e : _GEN_2025; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2027 = 8'heb == io_state_in_3 ? 8'h73 : _GEN_2026; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2028 = 8'hec == io_state_in_3 ? 8'h50 : _GEN_2027; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2029 = 8'hed == io_state_in_3 ? 8'h5d : _GEN_2028; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2030 = 8'hee == io_state_in_3 ? 8'h4a : _GEN_2029; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2031 = 8'hef == io_state_in_3 ? 8'h47 : _GEN_2030; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2032 = 8'hf0 == io_state_in_3 ? 8'hdc : _GEN_2031; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2033 = 8'hf1 == io_state_in_3 ? 8'hd1 : _GEN_2032; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2034 = 8'hf2 == io_state_in_3 ? 8'hc6 : _GEN_2033; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2035 = 8'hf3 == io_state_in_3 ? 8'hcb : _GEN_2034; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2036 = 8'hf4 == io_state_in_3 ? 8'he8 : _GEN_2035; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2037 = 8'hf5 == io_state_in_3 ? 8'he5 : _GEN_2036; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2038 = 8'hf6 == io_state_in_3 ? 8'hf2 : _GEN_2037; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2039 = 8'hf7 == io_state_in_3 ? 8'hff : _GEN_2038; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2040 = 8'hf8 == io_state_in_3 ? 8'hb4 : _GEN_2039; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2041 = 8'hf9 == io_state_in_3 ? 8'hb9 : _GEN_2040; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2042 = 8'hfa == io_state_in_3 ? 8'hae : _GEN_2041; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2043 = 8'hfb == io_state_in_3 ? 8'ha3 : _GEN_2042; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2044 = 8'hfc == io_state_in_3 ? 8'h80 : _GEN_2043; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2045 = 8'hfd == io_state_in_3 ? 8'h8d : _GEN_2044; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2046 = 8'hfe == io_state_in_3 ? 8'h9a : _GEN_2045; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2047 = 8'hff == io_state_in_3 ? 8'h97 : _GEN_2046; // @[InvMixColumns.scala 127:{89,89}]
  wire [7:0] _GEN_2049 = 8'h1 == io_state_in_0 ? 8'hd : 8'h0; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2050 = 8'h2 == io_state_in_0 ? 8'h1a : _GEN_2049; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2051 = 8'h3 == io_state_in_0 ? 8'h17 : _GEN_2050; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2052 = 8'h4 == io_state_in_0 ? 8'h34 : _GEN_2051; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2053 = 8'h5 == io_state_in_0 ? 8'h39 : _GEN_2052; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2054 = 8'h6 == io_state_in_0 ? 8'h2e : _GEN_2053; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2055 = 8'h7 == io_state_in_0 ? 8'h23 : _GEN_2054; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2056 = 8'h8 == io_state_in_0 ? 8'h68 : _GEN_2055; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2057 = 8'h9 == io_state_in_0 ? 8'h65 : _GEN_2056; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2058 = 8'ha == io_state_in_0 ? 8'h72 : _GEN_2057; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2059 = 8'hb == io_state_in_0 ? 8'h7f : _GEN_2058; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2060 = 8'hc == io_state_in_0 ? 8'h5c : _GEN_2059; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2061 = 8'hd == io_state_in_0 ? 8'h51 : _GEN_2060; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2062 = 8'he == io_state_in_0 ? 8'h46 : _GEN_2061; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2063 = 8'hf == io_state_in_0 ? 8'h4b : _GEN_2062; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2064 = 8'h10 == io_state_in_0 ? 8'hd0 : _GEN_2063; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2065 = 8'h11 == io_state_in_0 ? 8'hdd : _GEN_2064; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2066 = 8'h12 == io_state_in_0 ? 8'hca : _GEN_2065; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2067 = 8'h13 == io_state_in_0 ? 8'hc7 : _GEN_2066; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2068 = 8'h14 == io_state_in_0 ? 8'he4 : _GEN_2067; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2069 = 8'h15 == io_state_in_0 ? 8'he9 : _GEN_2068; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2070 = 8'h16 == io_state_in_0 ? 8'hfe : _GEN_2069; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2071 = 8'h17 == io_state_in_0 ? 8'hf3 : _GEN_2070; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2072 = 8'h18 == io_state_in_0 ? 8'hb8 : _GEN_2071; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2073 = 8'h19 == io_state_in_0 ? 8'hb5 : _GEN_2072; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2074 = 8'h1a == io_state_in_0 ? 8'ha2 : _GEN_2073; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2075 = 8'h1b == io_state_in_0 ? 8'haf : _GEN_2074; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2076 = 8'h1c == io_state_in_0 ? 8'h8c : _GEN_2075; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2077 = 8'h1d == io_state_in_0 ? 8'h81 : _GEN_2076; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2078 = 8'h1e == io_state_in_0 ? 8'h96 : _GEN_2077; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2079 = 8'h1f == io_state_in_0 ? 8'h9b : _GEN_2078; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2080 = 8'h20 == io_state_in_0 ? 8'hbb : _GEN_2079; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2081 = 8'h21 == io_state_in_0 ? 8'hb6 : _GEN_2080; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2082 = 8'h22 == io_state_in_0 ? 8'ha1 : _GEN_2081; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2083 = 8'h23 == io_state_in_0 ? 8'hac : _GEN_2082; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2084 = 8'h24 == io_state_in_0 ? 8'h8f : _GEN_2083; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2085 = 8'h25 == io_state_in_0 ? 8'h82 : _GEN_2084; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2086 = 8'h26 == io_state_in_0 ? 8'h95 : _GEN_2085; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2087 = 8'h27 == io_state_in_0 ? 8'h98 : _GEN_2086; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2088 = 8'h28 == io_state_in_0 ? 8'hd3 : _GEN_2087; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2089 = 8'h29 == io_state_in_0 ? 8'hde : _GEN_2088; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2090 = 8'h2a == io_state_in_0 ? 8'hc9 : _GEN_2089; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2091 = 8'h2b == io_state_in_0 ? 8'hc4 : _GEN_2090; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2092 = 8'h2c == io_state_in_0 ? 8'he7 : _GEN_2091; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2093 = 8'h2d == io_state_in_0 ? 8'hea : _GEN_2092; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2094 = 8'h2e == io_state_in_0 ? 8'hfd : _GEN_2093; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2095 = 8'h2f == io_state_in_0 ? 8'hf0 : _GEN_2094; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2096 = 8'h30 == io_state_in_0 ? 8'h6b : _GEN_2095; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2097 = 8'h31 == io_state_in_0 ? 8'h66 : _GEN_2096; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2098 = 8'h32 == io_state_in_0 ? 8'h71 : _GEN_2097; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2099 = 8'h33 == io_state_in_0 ? 8'h7c : _GEN_2098; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2100 = 8'h34 == io_state_in_0 ? 8'h5f : _GEN_2099; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2101 = 8'h35 == io_state_in_0 ? 8'h52 : _GEN_2100; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2102 = 8'h36 == io_state_in_0 ? 8'h45 : _GEN_2101; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2103 = 8'h37 == io_state_in_0 ? 8'h48 : _GEN_2102; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2104 = 8'h38 == io_state_in_0 ? 8'h3 : _GEN_2103; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2105 = 8'h39 == io_state_in_0 ? 8'he : _GEN_2104; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2106 = 8'h3a == io_state_in_0 ? 8'h19 : _GEN_2105; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2107 = 8'h3b == io_state_in_0 ? 8'h14 : _GEN_2106; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2108 = 8'h3c == io_state_in_0 ? 8'h37 : _GEN_2107; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2109 = 8'h3d == io_state_in_0 ? 8'h3a : _GEN_2108; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2110 = 8'h3e == io_state_in_0 ? 8'h2d : _GEN_2109; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2111 = 8'h3f == io_state_in_0 ? 8'h20 : _GEN_2110; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2112 = 8'h40 == io_state_in_0 ? 8'h6d : _GEN_2111; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2113 = 8'h41 == io_state_in_0 ? 8'h60 : _GEN_2112; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2114 = 8'h42 == io_state_in_0 ? 8'h77 : _GEN_2113; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2115 = 8'h43 == io_state_in_0 ? 8'h7a : _GEN_2114; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2116 = 8'h44 == io_state_in_0 ? 8'h59 : _GEN_2115; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2117 = 8'h45 == io_state_in_0 ? 8'h54 : _GEN_2116; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2118 = 8'h46 == io_state_in_0 ? 8'h43 : _GEN_2117; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2119 = 8'h47 == io_state_in_0 ? 8'h4e : _GEN_2118; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2120 = 8'h48 == io_state_in_0 ? 8'h5 : _GEN_2119; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2121 = 8'h49 == io_state_in_0 ? 8'h8 : _GEN_2120; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2122 = 8'h4a == io_state_in_0 ? 8'h1f : _GEN_2121; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2123 = 8'h4b == io_state_in_0 ? 8'h12 : _GEN_2122; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2124 = 8'h4c == io_state_in_0 ? 8'h31 : _GEN_2123; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2125 = 8'h4d == io_state_in_0 ? 8'h3c : _GEN_2124; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2126 = 8'h4e == io_state_in_0 ? 8'h2b : _GEN_2125; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2127 = 8'h4f == io_state_in_0 ? 8'h26 : _GEN_2126; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2128 = 8'h50 == io_state_in_0 ? 8'hbd : _GEN_2127; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2129 = 8'h51 == io_state_in_0 ? 8'hb0 : _GEN_2128; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2130 = 8'h52 == io_state_in_0 ? 8'ha7 : _GEN_2129; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2131 = 8'h53 == io_state_in_0 ? 8'haa : _GEN_2130; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2132 = 8'h54 == io_state_in_0 ? 8'h89 : _GEN_2131; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2133 = 8'h55 == io_state_in_0 ? 8'h84 : _GEN_2132; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2134 = 8'h56 == io_state_in_0 ? 8'h93 : _GEN_2133; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2135 = 8'h57 == io_state_in_0 ? 8'h9e : _GEN_2134; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2136 = 8'h58 == io_state_in_0 ? 8'hd5 : _GEN_2135; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2137 = 8'h59 == io_state_in_0 ? 8'hd8 : _GEN_2136; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2138 = 8'h5a == io_state_in_0 ? 8'hcf : _GEN_2137; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2139 = 8'h5b == io_state_in_0 ? 8'hc2 : _GEN_2138; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2140 = 8'h5c == io_state_in_0 ? 8'he1 : _GEN_2139; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2141 = 8'h5d == io_state_in_0 ? 8'hec : _GEN_2140; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2142 = 8'h5e == io_state_in_0 ? 8'hfb : _GEN_2141; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2143 = 8'h5f == io_state_in_0 ? 8'hf6 : _GEN_2142; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2144 = 8'h60 == io_state_in_0 ? 8'hd6 : _GEN_2143; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2145 = 8'h61 == io_state_in_0 ? 8'hdb : _GEN_2144; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2146 = 8'h62 == io_state_in_0 ? 8'hcc : _GEN_2145; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2147 = 8'h63 == io_state_in_0 ? 8'hc1 : _GEN_2146; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2148 = 8'h64 == io_state_in_0 ? 8'he2 : _GEN_2147; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2149 = 8'h65 == io_state_in_0 ? 8'hef : _GEN_2148; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2150 = 8'h66 == io_state_in_0 ? 8'hf8 : _GEN_2149; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2151 = 8'h67 == io_state_in_0 ? 8'hf5 : _GEN_2150; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2152 = 8'h68 == io_state_in_0 ? 8'hbe : _GEN_2151; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2153 = 8'h69 == io_state_in_0 ? 8'hb3 : _GEN_2152; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2154 = 8'h6a == io_state_in_0 ? 8'ha4 : _GEN_2153; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2155 = 8'h6b == io_state_in_0 ? 8'ha9 : _GEN_2154; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2156 = 8'h6c == io_state_in_0 ? 8'h8a : _GEN_2155; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2157 = 8'h6d == io_state_in_0 ? 8'h87 : _GEN_2156; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2158 = 8'h6e == io_state_in_0 ? 8'h90 : _GEN_2157; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2159 = 8'h6f == io_state_in_0 ? 8'h9d : _GEN_2158; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2160 = 8'h70 == io_state_in_0 ? 8'h6 : _GEN_2159; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2161 = 8'h71 == io_state_in_0 ? 8'hb : _GEN_2160; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2162 = 8'h72 == io_state_in_0 ? 8'h1c : _GEN_2161; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2163 = 8'h73 == io_state_in_0 ? 8'h11 : _GEN_2162; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2164 = 8'h74 == io_state_in_0 ? 8'h32 : _GEN_2163; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2165 = 8'h75 == io_state_in_0 ? 8'h3f : _GEN_2164; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2166 = 8'h76 == io_state_in_0 ? 8'h28 : _GEN_2165; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2167 = 8'h77 == io_state_in_0 ? 8'h25 : _GEN_2166; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2168 = 8'h78 == io_state_in_0 ? 8'h6e : _GEN_2167; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2169 = 8'h79 == io_state_in_0 ? 8'h63 : _GEN_2168; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2170 = 8'h7a == io_state_in_0 ? 8'h74 : _GEN_2169; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2171 = 8'h7b == io_state_in_0 ? 8'h79 : _GEN_2170; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2172 = 8'h7c == io_state_in_0 ? 8'h5a : _GEN_2171; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2173 = 8'h7d == io_state_in_0 ? 8'h57 : _GEN_2172; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2174 = 8'h7e == io_state_in_0 ? 8'h40 : _GEN_2173; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2175 = 8'h7f == io_state_in_0 ? 8'h4d : _GEN_2174; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2176 = 8'h80 == io_state_in_0 ? 8'hda : _GEN_2175; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2177 = 8'h81 == io_state_in_0 ? 8'hd7 : _GEN_2176; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2178 = 8'h82 == io_state_in_0 ? 8'hc0 : _GEN_2177; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2179 = 8'h83 == io_state_in_0 ? 8'hcd : _GEN_2178; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2180 = 8'h84 == io_state_in_0 ? 8'hee : _GEN_2179; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2181 = 8'h85 == io_state_in_0 ? 8'he3 : _GEN_2180; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2182 = 8'h86 == io_state_in_0 ? 8'hf4 : _GEN_2181; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2183 = 8'h87 == io_state_in_0 ? 8'hf9 : _GEN_2182; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2184 = 8'h88 == io_state_in_0 ? 8'hb2 : _GEN_2183; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2185 = 8'h89 == io_state_in_0 ? 8'hbf : _GEN_2184; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2186 = 8'h8a == io_state_in_0 ? 8'ha8 : _GEN_2185; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2187 = 8'h8b == io_state_in_0 ? 8'ha5 : _GEN_2186; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2188 = 8'h8c == io_state_in_0 ? 8'h86 : _GEN_2187; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2189 = 8'h8d == io_state_in_0 ? 8'h8b : _GEN_2188; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2190 = 8'h8e == io_state_in_0 ? 8'h9c : _GEN_2189; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2191 = 8'h8f == io_state_in_0 ? 8'h91 : _GEN_2190; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2192 = 8'h90 == io_state_in_0 ? 8'ha : _GEN_2191; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2193 = 8'h91 == io_state_in_0 ? 8'h7 : _GEN_2192; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2194 = 8'h92 == io_state_in_0 ? 8'h10 : _GEN_2193; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2195 = 8'h93 == io_state_in_0 ? 8'h1d : _GEN_2194; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2196 = 8'h94 == io_state_in_0 ? 8'h3e : _GEN_2195; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2197 = 8'h95 == io_state_in_0 ? 8'h33 : _GEN_2196; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2198 = 8'h96 == io_state_in_0 ? 8'h24 : _GEN_2197; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2199 = 8'h97 == io_state_in_0 ? 8'h29 : _GEN_2198; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2200 = 8'h98 == io_state_in_0 ? 8'h62 : _GEN_2199; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2201 = 8'h99 == io_state_in_0 ? 8'h6f : _GEN_2200; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2202 = 8'h9a == io_state_in_0 ? 8'h78 : _GEN_2201; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2203 = 8'h9b == io_state_in_0 ? 8'h75 : _GEN_2202; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2204 = 8'h9c == io_state_in_0 ? 8'h56 : _GEN_2203; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2205 = 8'h9d == io_state_in_0 ? 8'h5b : _GEN_2204; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2206 = 8'h9e == io_state_in_0 ? 8'h4c : _GEN_2205; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2207 = 8'h9f == io_state_in_0 ? 8'h41 : _GEN_2206; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2208 = 8'ha0 == io_state_in_0 ? 8'h61 : _GEN_2207; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2209 = 8'ha1 == io_state_in_0 ? 8'h6c : _GEN_2208; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2210 = 8'ha2 == io_state_in_0 ? 8'h7b : _GEN_2209; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2211 = 8'ha3 == io_state_in_0 ? 8'h76 : _GEN_2210; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2212 = 8'ha4 == io_state_in_0 ? 8'h55 : _GEN_2211; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2213 = 8'ha5 == io_state_in_0 ? 8'h58 : _GEN_2212; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2214 = 8'ha6 == io_state_in_0 ? 8'h4f : _GEN_2213; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2215 = 8'ha7 == io_state_in_0 ? 8'h42 : _GEN_2214; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2216 = 8'ha8 == io_state_in_0 ? 8'h9 : _GEN_2215; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2217 = 8'ha9 == io_state_in_0 ? 8'h4 : _GEN_2216; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2218 = 8'haa == io_state_in_0 ? 8'h13 : _GEN_2217; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2219 = 8'hab == io_state_in_0 ? 8'h1e : _GEN_2218; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2220 = 8'hac == io_state_in_0 ? 8'h3d : _GEN_2219; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2221 = 8'had == io_state_in_0 ? 8'h30 : _GEN_2220; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2222 = 8'hae == io_state_in_0 ? 8'h27 : _GEN_2221; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2223 = 8'haf == io_state_in_0 ? 8'h2a : _GEN_2222; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2224 = 8'hb0 == io_state_in_0 ? 8'hb1 : _GEN_2223; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2225 = 8'hb1 == io_state_in_0 ? 8'hbc : _GEN_2224; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2226 = 8'hb2 == io_state_in_0 ? 8'hab : _GEN_2225; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2227 = 8'hb3 == io_state_in_0 ? 8'ha6 : _GEN_2226; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2228 = 8'hb4 == io_state_in_0 ? 8'h85 : _GEN_2227; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2229 = 8'hb5 == io_state_in_0 ? 8'h88 : _GEN_2228; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2230 = 8'hb6 == io_state_in_0 ? 8'h9f : _GEN_2229; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2231 = 8'hb7 == io_state_in_0 ? 8'h92 : _GEN_2230; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2232 = 8'hb8 == io_state_in_0 ? 8'hd9 : _GEN_2231; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2233 = 8'hb9 == io_state_in_0 ? 8'hd4 : _GEN_2232; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2234 = 8'hba == io_state_in_0 ? 8'hc3 : _GEN_2233; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2235 = 8'hbb == io_state_in_0 ? 8'hce : _GEN_2234; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2236 = 8'hbc == io_state_in_0 ? 8'hed : _GEN_2235; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2237 = 8'hbd == io_state_in_0 ? 8'he0 : _GEN_2236; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2238 = 8'hbe == io_state_in_0 ? 8'hf7 : _GEN_2237; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2239 = 8'hbf == io_state_in_0 ? 8'hfa : _GEN_2238; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2240 = 8'hc0 == io_state_in_0 ? 8'hb7 : _GEN_2239; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2241 = 8'hc1 == io_state_in_0 ? 8'hba : _GEN_2240; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2242 = 8'hc2 == io_state_in_0 ? 8'had : _GEN_2241; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2243 = 8'hc3 == io_state_in_0 ? 8'ha0 : _GEN_2242; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2244 = 8'hc4 == io_state_in_0 ? 8'h83 : _GEN_2243; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2245 = 8'hc5 == io_state_in_0 ? 8'h8e : _GEN_2244; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2246 = 8'hc6 == io_state_in_0 ? 8'h99 : _GEN_2245; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2247 = 8'hc7 == io_state_in_0 ? 8'h94 : _GEN_2246; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2248 = 8'hc8 == io_state_in_0 ? 8'hdf : _GEN_2247; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2249 = 8'hc9 == io_state_in_0 ? 8'hd2 : _GEN_2248; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2250 = 8'hca == io_state_in_0 ? 8'hc5 : _GEN_2249; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2251 = 8'hcb == io_state_in_0 ? 8'hc8 : _GEN_2250; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2252 = 8'hcc == io_state_in_0 ? 8'heb : _GEN_2251; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2253 = 8'hcd == io_state_in_0 ? 8'he6 : _GEN_2252; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2254 = 8'hce == io_state_in_0 ? 8'hf1 : _GEN_2253; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2255 = 8'hcf == io_state_in_0 ? 8'hfc : _GEN_2254; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2256 = 8'hd0 == io_state_in_0 ? 8'h67 : _GEN_2255; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2257 = 8'hd1 == io_state_in_0 ? 8'h6a : _GEN_2256; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2258 = 8'hd2 == io_state_in_0 ? 8'h7d : _GEN_2257; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2259 = 8'hd3 == io_state_in_0 ? 8'h70 : _GEN_2258; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2260 = 8'hd4 == io_state_in_0 ? 8'h53 : _GEN_2259; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2261 = 8'hd5 == io_state_in_0 ? 8'h5e : _GEN_2260; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2262 = 8'hd6 == io_state_in_0 ? 8'h49 : _GEN_2261; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2263 = 8'hd7 == io_state_in_0 ? 8'h44 : _GEN_2262; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2264 = 8'hd8 == io_state_in_0 ? 8'hf : _GEN_2263; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2265 = 8'hd9 == io_state_in_0 ? 8'h2 : _GEN_2264; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2266 = 8'hda == io_state_in_0 ? 8'h15 : _GEN_2265; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2267 = 8'hdb == io_state_in_0 ? 8'h18 : _GEN_2266; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2268 = 8'hdc == io_state_in_0 ? 8'h3b : _GEN_2267; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2269 = 8'hdd == io_state_in_0 ? 8'h36 : _GEN_2268; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2270 = 8'hde == io_state_in_0 ? 8'h21 : _GEN_2269; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2271 = 8'hdf == io_state_in_0 ? 8'h2c : _GEN_2270; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2272 = 8'he0 == io_state_in_0 ? 8'hc : _GEN_2271; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2273 = 8'he1 == io_state_in_0 ? 8'h1 : _GEN_2272; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2274 = 8'he2 == io_state_in_0 ? 8'h16 : _GEN_2273; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2275 = 8'he3 == io_state_in_0 ? 8'h1b : _GEN_2274; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2276 = 8'he4 == io_state_in_0 ? 8'h38 : _GEN_2275; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2277 = 8'he5 == io_state_in_0 ? 8'h35 : _GEN_2276; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2278 = 8'he6 == io_state_in_0 ? 8'h22 : _GEN_2277; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2279 = 8'he7 == io_state_in_0 ? 8'h2f : _GEN_2278; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2280 = 8'he8 == io_state_in_0 ? 8'h64 : _GEN_2279; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2281 = 8'he9 == io_state_in_0 ? 8'h69 : _GEN_2280; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2282 = 8'hea == io_state_in_0 ? 8'h7e : _GEN_2281; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2283 = 8'heb == io_state_in_0 ? 8'h73 : _GEN_2282; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2284 = 8'hec == io_state_in_0 ? 8'h50 : _GEN_2283; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2285 = 8'hed == io_state_in_0 ? 8'h5d : _GEN_2284; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2286 = 8'hee == io_state_in_0 ? 8'h4a : _GEN_2285; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2287 = 8'hef == io_state_in_0 ? 8'h47 : _GEN_2286; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2288 = 8'hf0 == io_state_in_0 ? 8'hdc : _GEN_2287; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2289 = 8'hf1 == io_state_in_0 ? 8'hd1 : _GEN_2288; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2290 = 8'hf2 == io_state_in_0 ? 8'hc6 : _GEN_2289; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2291 = 8'hf3 == io_state_in_0 ? 8'hcb : _GEN_2290; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2292 = 8'hf4 == io_state_in_0 ? 8'he8 : _GEN_2291; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2293 = 8'hf5 == io_state_in_0 ? 8'he5 : _GEN_2292; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2294 = 8'hf6 == io_state_in_0 ? 8'hf2 : _GEN_2293; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2295 = 8'hf7 == io_state_in_0 ? 8'hff : _GEN_2294; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2296 = 8'hf8 == io_state_in_0 ? 8'hb4 : _GEN_2295; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2297 = 8'hf9 == io_state_in_0 ? 8'hb9 : _GEN_2296; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2298 = 8'hfa == io_state_in_0 ? 8'hae : _GEN_2297; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2299 = 8'hfb == io_state_in_0 ? 8'ha3 : _GEN_2298; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2300 = 8'hfc == io_state_in_0 ? 8'h80 : _GEN_2299; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2301 = 8'hfd == io_state_in_0 ? 8'h8d : _GEN_2300; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2302 = 8'hfe == io_state_in_0 ? 8'h9a : _GEN_2301; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2303 = 8'hff == io_state_in_0 ? 8'h97 : _GEN_2302; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2305 = 8'h1 == io_state_in_1 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2306 = 8'h2 == io_state_in_1 ? 8'h12 : _GEN_2305; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2307 = 8'h3 == io_state_in_1 ? 8'h1b : _GEN_2306; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2308 = 8'h4 == io_state_in_1 ? 8'h24 : _GEN_2307; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2309 = 8'h5 == io_state_in_1 ? 8'h2d : _GEN_2308; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2310 = 8'h6 == io_state_in_1 ? 8'h36 : _GEN_2309; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2311 = 8'h7 == io_state_in_1 ? 8'h3f : _GEN_2310; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2312 = 8'h8 == io_state_in_1 ? 8'h48 : _GEN_2311; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2313 = 8'h9 == io_state_in_1 ? 8'h41 : _GEN_2312; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2314 = 8'ha == io_state_in_1 ? 8'h5a : _GEN_2313; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2315 = 8'hb == io_state_in_1 ? 8'h53 : _GEN_2314; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2316 = 8'hc == io_state_in_1 ? 8'h6c : _GEN_2315; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2317 = 8'hd == io_state_in_1 ? 8'h65 : _GEN_2316; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2318 = 8'he == io_state_in_1 ? 8'h7e : _GEN_2317; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2319 = 8'hf == io_state_in_1 ? 8'h77 : _GEN_2318; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2320 = 8'h10 == io_state_in_1 ? 8'h90 : _GEN_2319; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2321 = 8'h11 == io_state_in_1 ? 8'h99 : _GEN_2320; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2322 = 8'h12 == io_state_in_1 ? 8'h82 : _GEN_2321; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2323 = 8'h13 == io_state_in_1 ? 8'h8b : _GEN_2322; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2324 = 8'h14 == io_state_in_1 ? 8'hb4 : _GEN_2323; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2325 = 8'h15 == io_state_in_1 ? 8'hbd : _GEN_2324; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2326 = 8'h16 == io_state_in_1 ? 8'ha6 : _GEN_2325; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2327 = 8'h17 == io_state_in_1 ? 8'haf : _GEN_2326; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2328 = 8'h18 == io_state_in_1 ? 8'hd8 : _GEN_2327; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2329 = 8'h19 == io_state_in_1 ? 8'hd1 : _GEN_2328; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2330 = 8'h1a == io_state_in_1 ? 8'hca : _GEN_2329; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2331 = 8'h1b == io_state_in_1 ? 8'hc3 : _GEN_2330; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2332 = 8'h1c == io_state_in_1 ? 8'hfc : _GEN_2331; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2333 = 8'h1d == io_state_in_1 ? 8'hf5 : _GEN_2332; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2334 = 8'h1e == io_state_in_1 ? 8'hee : _GEN_2333; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2335 = 8'h1f == io_state_in_1 ? 8'he7 : _GEN_2334; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2336 = 8'h20 == io_state_in_1 ? 8'h3b : _GEN_2335; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2337 = 8'h21 == io_state_in_1 ? 8'h32 : _GEN_2336; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2338 = 8'h22 == io_state_in_1 ? 8'h29 : _GEN_2337; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2339 = 8'h23 == io_state_in_1 ? 8'h20 : _GEN_2338; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2340 = 8'h24 == io_state_in_1 ? 8'h1f : _GEN_2339; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2341 = 8'h25 == io_state_in_1 ? 8'h16 : _GEN_2340; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2342 = 8'h26 == io_state_in_1 ? 8'hd : _GEN_2341; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2343 = 8'h27 == io_state_in_1 ? 8'h4 : _GEN_2342; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2344 = 8'h28 == io_state_in_1 ? 8'h73 : _GEN_2343; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2345 = 8'h29 == io_state_in_1 ? 8'h7a : _GEN_2344; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2346 = 8'h2a == io_state_in_1 ? 8'h61 : _GEN_2345; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2347 = 8'h2b == io_state_in_1 ? 8'h68 : _GEN_2346; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2348 = 8'h2c == io_state_in_1 ? 8'h57 : _GEN_2347; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2349 = 8'h2d == io_state_in_1 ? 8'h5e : _GEN_2348; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2350 = 8'h2e == io_state_in_1 ? 8'h45 : _GEN_2349; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2351 = 8'h2f == io_state_in_1 ? 8'h4c : _GEN_2350; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2352 = 8'h30 == io_state_in_1 ? 8'hab : _GEN_2351; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2353 = 8'h31 == io_state_in_1 ? 8'ha2 : _GEN_2352; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2354 = 8'h32 == io_state_in_1 ? 8'hb9 : _GEN_2353; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2355 = 8'h33 == io_state_in_1 ? 8'hb0 : _GEN_2354; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2356 = 8'h34 == io_state_in_1 ? 8'h8f : _GEN_2355; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2357 = 8'h35 == io_state_in_1 ? 8'h86 : _GEN_2356; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2358 = 8'h36 == io_state_in_1 ? 8'h9d : _GEN_2357; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2359 = 8'h37 == io_state_in_1 ? 8'h94 : _GEN_2358; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2360 = 8'h38 == io_state_in_1 ? 8'he3 : _GEN_2359; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2361 = 8'h39 == io_state_in_1 ? 8'hea : _GEN_2360; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2362 = 8'h3a == io_state_in_1 ? 8'hf1 : _GEN_2361; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2363 = 8'h3b == io_state_in_1 ? 8'hf8 : _GEN_2362; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2364 = 8'h3c == io_state_in_1 ? 8'hc7 : _GEN_2363; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2365 = 8'h3d == io_state_in_1 ? 8'hce : _GEN_2364; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2366 = 8'h3e == io_state_in_1 ? 8'hd5 : _GEN_2365; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2367 = 8'h3f == io_state_in_1 ? 8'hdc : _GEN_2366; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2368 = 8'h40 == io_state_in_1 ? 8'h76 : _GEN_2367; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2369 = 8'h41 == io_state_in_1 ? 8'h7f : _GEN_2368; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2370 = 8'h42 == io_state_in_1 ? 8'h64 : _GEN_2369; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2371 = 8'h43 == io_state_in_1 ? 8'h6d : _GEN_2370; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2372 = 8'h44 == io_state_in_1 ? 8'h52 : _GEN_2371; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2373 = 8'h45 == io_state_in_1 ? 8'h5b : _GEN_2372; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2374 = 8'h46 == io_state_in_1 ? 8'h40 : _GEN_2373; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2375 = 8'h47 == io_state_in_1 ? 8'h49 : _GEN_2374; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2376 = 8'h48 == io_state_in_1 ? 8'h3e : _GEN_2375; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2377 = 8'h49 == io_state_in_1 ? 8'h37 : _GEN_2376; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2378 = 8'h4a == io_state_in_1 ? 8'h2c : _GEN_2377; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2379 = 8'h4b == io_state_in_1 ? 8'h25 : _GEN_2378; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2380 = 8'h4c == io_state_in_1 ? 8'h1a : _GEN_2379; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2381 = 8'h4d == io_state_in_1 ? 8'h13 : _GEN_2380; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2382 = 8'h4e == io_state_in_1 ? 8'h8 : _GEN_2381; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2383 = 8'h4f == io_state_in_1 ? 8'h1 : _GEN_2382; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2384 = 8'h50 == io_state_in_1 ? 8'he6 : _GEN_2383; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2385 = 8'h51 == io_state_in_1 ? 8'hef : _GEN_2384; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2386 = 8'h52 == io_state_in_1 ? 8'hf4 : _GEN_2385; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2387 = 8'h53 == io_state_in_1 ? 8'hfd : _GEN_2386; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2388 = 8'h54 == io_state_in_1 ? 8'hc2 : _GEN_2387; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2389 = 8'h55 == io_state_in_1 ? 8'hcb : _GEN_2388; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2390 = 8'h56 == io_state_in_1 ? 8'hd0 : _GEN_2389; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2391 = 8'h57 == io_state_in_1 ? 8'hd9 : _GEN_2390; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2392 = 8'h58 == io_state_in_1 ? 8'hae : _GEN_2391; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2393 = 8'h59 == io_state_in_1 ? 8'ha7 : _GEN_2392; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2394 = 8'h5a == io_state_in_1 ? 8'hbc : _GEN_2393; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2395 = 8'h5b == io_state_in_1 ? 8'hb5 : _GEN_2394; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2396 = 8'h5c == io_state_in_1 ? 8'h8a : _GEN_2395; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2397 = 8'h5d == io_state_in_1 ? 8'h83 : _GEN_2396; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2398 = 8'h5e == io_state_in_1 ? 8'h98 : _GEN_2397; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2399 = 8'h5f == io_state_in_1 ? 8'h91 : _GEN_2398; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2400 = 8'h60 == io_state_in_1 ? 8'h4d : _GEN_2399; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2401 = 8'h61 == io_state_in_1 ? 8'h44 : _GEN_2400; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2402 = 8'h62 == io_state_in_1 ? 8'h5f : _GEN_2401; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2403 = 8'h63 == io_state_in_1 ? 8'h56 : _GEN_2402; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2404 = 8'h64 == io_state_in_1 ? 8'h69 : _GEN_2403; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2405 = 8'h65 == io_state_in_1 ? 8'h60 : _GEN_2404; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2406 = 8'h66 == io_state_in_1 ? 8'h7b : _GEN_2405; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2407 = 8'h67 == io_state_in_1 ? 8'h72 : _GEN_2406; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2408 = 8'h68 == io_state_in_1 ? 8'h5 : _GEN_2407; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2409 = 8'h69 == io_state_in_1 ? 8'hc : _GEN_2408; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2410 = 8'h6a == io_state_in_1 ? 8'h17 : _GEN_2409; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2411 = 8'h6b == io_state_in_1 ? 8'h1e : _GEN_2410; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2412 = 8'h6c == io_state_in_1 ? 8'h21 : _GEN_2411; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2413 = 8'h6d == io_state_in_1 ? 8'h28 : _GEN_2412; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2414 = 8'h6e == io_state_in_1 ? 8'h33 : _GEN_2413; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2415 = 8'h6f == io_state_in_1 ? 8'h3a : _GEN_2414; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2416 = 8'h70 == io_state_in_1 ? 8'hdd : _GEN_2415; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2417 = 8'h71 == io_state_in_1 ? 8'hd4 : _GEN_2416; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2418 = 8'h72 == io_state_in_1 ? 8'hcf : _GEN_2417; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2419 = 8'h73 == io_state_in_1 ? 8'hc6 : _GEN_2418; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2420 = 8'h74 == io_state_in_1 ? 8'hf9 : _GEN_2419; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2421 = 8'h75 == io_state_in_1 ? 8'hf0 : _GEN_2420; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2422 = 8'h76 == io_state_in_1 ? 8'heb : _GEN_2421; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2423 = 8'h77 == io_state_in_1 ? 8'he2 : _GEN_2422; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2424 = 8'h78 == io_state_in_1 ? 8'h95 : _GEN_2423; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2425 = 8'h79 == io_state_in_1 ? 8'h9c : _GEN_2424; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2426 = 8'h7a == io_state_in_1 ? 8'h87 : _GEN_2425; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2427 = 8'h7b == io_state_in_1 ? 8'h8e : _GEN_2426; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2428 = 8'h7c == io_state_in_1 ? 8'hb1 : _GEN_2427; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2429 = 8'h7d == io_state_in_1 ? 8'hb8 : _GEN_2428; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2430 = 8'h7e == io_state_in_1 ? 8'ha3 : _GEN_2429; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2431 = 8'h7f == io_state_in_1 ? 8'haa : _GEN_2430; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2432 = 8'h80 == io_state_in_1 ? 8'hec : _GEN_2431; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2433 = 8'h81 == io_state_in_1 ? 8'he5 : _GEN_2432; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2434 = 8'h82 == io_state_in_1 ? 8'hfe : _GEN_2433; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2435 = 8'h83 == io_state_in_1 ? 8'hf7 : _GEN_2434; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2436 = 8'h84 == io_state_in_1 ? 8'hc8 : _GEN_2435; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2437 = 8'h85 == io_state_in_1 ? 8'hc1 : _GEN_2436; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2438 = 8'h86 == io_state_in_1 ? 8'hda : _GEN_2437; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2439 = 8'h87 == io_state_in_1 ? 8'hd3 : _GEN_2438; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2440 = 8'h88 == io_state_in_1 ? 8'ha4 : _GEN_2439; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2441 = 8'h89 == io_state_in_1 ? 8'had : _GEN_2440; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2442 = 8'h8a == io_state_in_1 ? 8'hb6 : _GEN_2441; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2443 = 8'h8b == io_state_in_1 ? 8'hbf : _GEN_2442; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2444 = 8'h8c == io_state_in_1 ? 8'h80 : _GEN_2443; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2445 = 8'h8d == io_state_in_1 ? 8'h89 : _GEN_2444; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2446 = 8'h8e == io_state_in_1 ? 8'h92 : _GEN_2445; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2447 = 8'h8f == io_state_in_1 ? 8'h9b : _GEN_2446; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2448 = 8'h90 == io_state_in_1 ? 8'h7c : _GEN_2447; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2449 = 8'h91 == io_state_in_1 ? 8'h75 : _GEN_2448; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2450 = 8'h92 == io_state_in_1 ? 8'h6e : _GEN_2449; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2451 = 8'h93 == io_state_in_1 ? 8'h67 : _GEN_2450; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2452 = 8'h94 == io_state_in_1 ? 8'h58 : _GEN_2451; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2453 = 8'h95 == io_state_in_1 ? 8'h51 : _GEN_2452; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2454 = 8'h96 == io_state_in_1 ? 8'h4a : _GEN_2453; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2455 = 8'h97 == io_state_in_1 ? 8'h43 : _GEN_2454; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2456 = 8'h98 == io_state_in_1 ? 8'h34 : _GEN_2455; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2457 = 8'h99 == io_state_in_1 ? 8'h3d : _GEN_2456; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2458 = 8'h9a == io_state_in_1 ? 8'h26 : _GEN_2457; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2459 = 8'h9b == io_state_in_1 ? 8'h2f : _GEN_2458; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2460 = 8'h9c == io_state_in_1 ? 8'h10 : _GEN_2459; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2461 = 8'h9d == io_state_in_1 ? 8'h19 : _GEN_2460; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2462 = 8'h9e == io_state_in_1 ? 8'h2 : _GEN_2461; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2463 = 8'h9f == io_state_in_1 ? 8'hb : _GEN_2462; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2464 = 8'ha0 == io_state_in_1 ? 8'hd7 : _GEN_2463; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2465 = 8'ha1 == io_state_in_1 ? 8'hde : _GEN_2464; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2466 = 8'ha2 == io_state_in_1 ? 8'hc5 : _GEN_2465; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2467 = 8'ha3 == io_state_in_1 ? 8'hcc : _GEN_2466; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2468 = 8'ha4 == io_state_in_1 ? 8'hf3 : _GEN_2467; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2469 = 8'ha5 == io_state_in_1 ? 8'hfa : _GEN_2468; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2470 = 8'ha6 == io_state_in_1 ? 8'he1 : _GEN_2469; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2471 = 8'ha7 == io_state_in_1 ? 8'he8 : _GEN_2470; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2472 = 8'ha8 == io_state_in_1 ? 8'h9f : _GEN_2471; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2473 = 8'ha9 == io_state_in_1 ? 8'h96 : _GEN_2472; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2474 = 8'haa == io_state_in_1 ? 8'h8d : _GEN_2473; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2475 = 8'hab == io_state_in_1 ? 8'h84 : _GEN_2474; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2476 = 8'hac == io_state_in_1 ? 8'hbb : _GEN_2475; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2477 = 8'had == io_state_in_1 ? 8'hb2 : _GEN_2476; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2478 = 8'hae == io_state_in_1 ? 8'ha9 : _GEN_2477; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2479 = 8'haf == io_state_in_1 ? 8'ha0 : _GEN_2478; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2480 = 8'hb0 == io_state_in_1 ? 8'h47 : _GEN_2479; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2481 = 8'hb1 == io_state_in_1 ? 8'h4e : _GEN_2480; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2482 = 8'hb2 == io_state_in_1 ? 8'h55 : _GEN_2481; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2483 = 8'hb3 == io_state_in_1 ? 8'h5c : _GEN_2482; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2484 = 8'hb4 == io_state_in_1 ? 8'h63 : _GEN_2483; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2485 = 8'hb5 == io_state_in_1 ? 8'h6a : _GEN_2484; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2486 = 8'hb6 == io_state_in_1 ? 8'h71 : _GEN_2485; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2487 = 8'hb7 == io_state_in_1 ? 8'h78 : _GEN_2486; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2488 = 8'hb8 == io_state_in_1 ? 8'hf : _GEN_2487; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2489 = 8'hb9 == io_state_in_1 ? 8'h6 : _GEN_2488; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2490 = 8'hba == io_state_in_1 ? 8'h1d : _GEN_2489; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2491 = 8'hbb == io_state_in_1 ? 8'h14 : _GEN_2490; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2492 = 8'hbc == io_state_in_1 ? 8'h2b : _GEN_2491; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2493 = 8'hbd == io_state_in_1 ? 8'h22 : _GEN_2492; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2494 = 8'hbe == io_state_in_1 ? 8'h39 : _GEN_2493; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2495 = 8'hbf == io_state_in_1 ? 8'h30 : _GEN_2494; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2496 = 8'hc0 == io_state_in_1 ? 8'h9a : _GEN_2495; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2497 = 8'hc1 == io_state_in_1 ? 8'h93 : _GEN_2496; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2498 = 8'hc2 == io_state_in_1 ? 8'h88 : _GEN_2497; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2499 = 8'hc3 == io_state_in_1 ? 8'h81 : _GEN_2498; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2500 = 8'hc4 == io_state_in_1 ? 8'hbe : _GEN_2499; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2501 = 8'hc5 == io_state_in_1 ? 8'hb7 : _GEN_2500; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2502 = 8'hc6 == io_state_in_1 ? 8'hac : _GEN_2501; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2503 = 8'hc7 == io_state_in_1 ? 8'ha5 : _GEN_2502; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2504 = 8'hc8 == io_state_in_1 ? 8'hd2 : _GEN_2503; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2505 = 8'hc9 == io_state_in_1 ? 8'hdb : _GEN_2504; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2506 = 8'hca == io_state_in_1 ? 8'hc0 : _GEN_2505; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2507 = 8'hcb == io_state_in_1 ? 8'hc9 : _GEN_2506; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2508 = 8'hcc == io_state_in_1 ? 8'hf6 : _GEN_2507; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2509 = 8'hcd == io_state_in_1 ? 8'hff : _GEN_2508; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2510 = 8'hce == io_state_in_1 ? 8'he4 : _GEN_2509; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2511 = 8'hcf == io_state_in_1 ? 8'hed : _GEN_2510; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2512 = 8'hd0 == io_state_in_1 ? 8'ha : _GEN_2511; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2513 = 8'hd1 == io_state_in_1 ? 8'h3 : _GEN_2512; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2514 = 8'hd2 == io_state_in_1 ? 8'h18 : _GEN_2513; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2515 = 8'hd3 == io_state_in_1 ? 8'h11 : _GEN_2514; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2516 = 8'hd4 == io_state_in_1 ? 8'h2e : _GEN_2515; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2517 = 8'hd5 == io_state_in_1 ? 8'h27 : _GEN_2516; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2518 = 8'hd6 == io_state_in_1 ? 8'h3c : _GEN_2517; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2519 = 8'hd7 == io_state_in_1 ? 8'h35 : _GEN_2518; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2520 = 8'hd8 == io_state_in_1 ? 8'h42 : _GEN_2519; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2521 = 8'hd9 == io_state_in_1 ? 8'h4b : _GEN_2520; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2522 = 8'hda == io_state_in_1 ? 8'h50 : _GEN_2521; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2523 = 8'hdb == io_state_in_1 ? 8'h59 : _GEN_2522; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2524 = 8'hdc == io_state_in_1 ? 8'h66 : _GEN_2523; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2525 = 8'hdd == io_state_in_1 ? 8'h6f : _GEN_2524; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2526 = 8'hde == io_state_in_1 ? 8'h74 : _GEN_2525; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2527 = 8'hdf == io_state_in_1 ? 8'h7d : _GEN_2526; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2528 = 8'he0 == io_state_in_1 ? 8'ha1 : _GEN_2527; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2529 = 8'he1 == io_state_in_1 ? 8'ha8 : _GEN_2528; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2530 = 8'he2 == io_state_in_1 ? 8'hb3 : _GEN_2529; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2531 = 8'he3 == io_state_in_1 ? 8'hba : _GEN_2530; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2532 = 8'he4 == io_state_in_1 ? 8'h85 : _GEN_2531; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2533 = 8'he5 == io_state_in_1 ? 8'h8c : _GEN_2532; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2534 = 8'he6 == io_state_in_1 ? 8'h97 : _GEN_2533; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2535 = 8'he7 == io_state_in_1 ? 8'h9e : _GEN_2534; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2536 = 8'he8 == io_state_in_1 ? 8'he9 : _GEN_2535; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2537 = 8'he9 == io_state_in_1 ? 8'he0 : _GEN_2536; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2538 = 8'hea == io_state_in_1 ? 8'hfb : _GEN_2537; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2539 = 8'heb == io_state_in_1 ? 8'hf2 : _GEN_2538; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2540 = 8'hec == io_state_in_1 ? 8'hcd : _GEN_2539; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2541 = 8'hed == io_state_in_1 ? 8'hc4 : _GEN_2540; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2542 = 8'hee == io_state_in_1 ? 8'hdf : _GEN_2541; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2543 = 8'hef == io_state_in_1 ? 8'hd6 : _GEN_2542; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2544 = 8'hf0 == io_state_in_1 ? 8'h31 : _GEN_2543; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2545 = 8'hf1 == io_state_in_1 ? 8'h38 : _GEN_2544; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2546 = 8'hf2 == io_state_in_1 ? 8'h23 : _GEN_2545; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2547 = 8'hf3 == io_state_in_1 ? 8'h2a : _GEN_2546; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2548 = 8'hf4 == io_state_in_1 ? 8'h15 : _GEN_2547; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2549 = 8'hf5 == io_state_in_1 ? 8'h1c : _GEN_2548; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2550 = 8'hf6 == io_state_in_1 ? 8'h7 : _GEN_2549; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2551 = 8'hf7 == io_state_in_1 ? 8'he : _GEN_2550; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2552 = 8'hf8 == io_state_in_1 ? 8'h79 : _GEN_2551; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2553 = 8'hf9 == io_state_in_1 ? 8'h70 : _GEN_2552; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2554 = 8'hfa == io_state_in_1 ? 8'h6b : _GEN_2553; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2555 = 8'hfb == io_state_in_1 ? 8'h62 : _GEN_2554; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2556 = 8'hfc == io_state_in_1 ? 8'h5d : _GEN_2555; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2557 = 8'hfd == io_state_in_1 ? 8'h54 : _GEN_2556; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2558 = 8'hfe == io_state_in_1 ? 8'h4f : _GEN_2557; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_2559 = 8'hff == io_state_in_1 ? 8'h46 : _GEN_2558; // @[InvMixColumns.scala 128:{41,41}]
  wire [7:0] _tmp_state_2_T = _GEN_2303 ^ _GEN_2559; // @[InvMixColumns.scala 128:41]
  wire [7:0] _GEN_2561 = 8'h1 == io_state_in_2 ? 8'he : 8'h0; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2562 = 8'h2 == io_state_in_2 ? 8'h1c : _GEN_2561; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2563 = 8'h3 == io_state_in_2 ? 8'h12 : _GEN_2562; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2564 = 8'h4 == io_state_in_2 ? 8'h38 : _GEN_2563; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2565 = 8'h5 == io_state_in_2 ? 8'h36 : _GEN_2564; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2566 = 8'h6 == io_state_in_2 ? 8'h24 : _GEN_2565; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2567 = 8'h7 == io_state_in_2 ? 8'h2a : _GEN_2566; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2568 = 8'h8 == io_state_in_2 ? 8'h70 : _GEN_2567; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2569 = 8'h9 == io_state_in_2 ? 8'h7e : _GEN_2568; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2570 = 8'ha == io_state_in_2 ? 8'h6c : _GEN_2569; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2571 = 8'hb == io_state_in_2 ? 8'h62 : _GEN_2570; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2572 = 8'hc == io_state_in_2 ? 8'h48 : _GEN_2571; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2573 = 8'hd == io_state_in_2 ? 8'h46 : _GEN_2572; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2574 = 8'he == io_state_in_2 ? 8'h54 : _GEN_2573; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2575 = 8'hf == io_state_in_2 ? 8'h5a : _GEN_2574; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2576 = 8'h10 == io_state_in_2 ? 8'he0 : _GEN_2575; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2577 = 8'h11 == io_state_in_2 ? 8'hee : _GEN_2576; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2578 = 8'h12 == io_state_in_2 ? 8'hfc : _GEN_2577; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2579 = 8'h13 == io_state_in_2 ? 8'hf2 : _GEN_2578; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2580 = 8'h14 == io_state_in_2 ? 8'hd8 : _GEN_2579; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2581 = 8'h15 == io_state_in_2 ? 8'hd6 : _GEN_2580; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2582 = 8'h16 == io_state_in_2 ? 8'hc4 : _GEN_2581; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2583 = 8'h17 == io_state_in_2 ? 8'hca : _GEN_2582; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2584 = 8'h18 == io_state_in_2 ? 8'h90 : _GEN_2583; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2585 = 8'h19 == io_state_in_2 ? 8'h9e : _GEN_2584; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2586 = 8'h1a == io_state_in_2 ? 8'h8c : _GEN_2585; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2587 = 8'h1b == io_state_in_2 ? 8'h82 : _GEN_2586; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2588 = 8'h1c == io_state_in_2 ? 8'ha8 : _GEN_2587; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2589 = 8'h1d == io_state_in_2 ? 8'ha6 : _GEN_2588; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2590 = 8'h1e == io_state_in_2 ? 8'hb4 : _GEN_2589; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2591 = 8'h1f == io_state_in_2 ? 8'hba : _GEN_2590; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2592 = 8'h20 == io_state_in_2 ? 8'hdb : _GEN_2591; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2593 = 8'h21 == io_state_in_2 ? 8'hd5 : _GEN_2592; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2594 = 8'h22 == io_state_in_2 ? 8'hc7 : _GEN_2593; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2595 = 8'h23 == io_state_in_2 ? 8'hc9 : _GEN_2594; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2596 = 8'h24 == io_state_in_2 ? 8'he3 : _GEN_2595; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2597 = 8'h25 == io_state_in_2 ? 8'hed : _GEN_2596; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2598 = 8'h26 == io_state_in_2 ? 8'hff : _GEN_2597; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2599 = 8'h27 == io_state_in_2 ? 8'hf1 : _GEN_2598; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2600 = 8'h28 == io_state_in_2 ? 8'hab : _GEN_2599; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2601 = 8'h29 == io_state_in_2 ? 8'ha5 : _GEN_2600; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2602 = 8'h2a == io_state_in_2 ? 8'hb7 : _GEN_2601; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2603 = 8'h2b == io_state_in_2 ? 8'hb9 : _GEN_2602; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2604 = 8'h2c == io_state_in_2 ? 8'h93 : _GEN_2603; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2605 = 8'h2d == io_state_in_2 ? 8'h9d : _GEN_2604; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2606 = 8'h2e == io_state_in_2 ? 8'h8f : _GEN_2605; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2607 = 8'h2f == io_state_in_2 ? 8'h81 : _GEN_2606; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2608 = 8'h30 == io_state_in_2 ? 8'h3b : _GEN_2607; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2609 = 8'h31 == io_state_in_2 ? 8'h35 : _GEN_2608; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2610 = 8'h32 == io_state_in_2 ? 8'h27 : _GEN_2609; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2611 = 8'h33 == io_state_in_2 ? 8'h29 : _GEN_2610; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2612 = 8'h34 == io_state_in_2 ? 8'h3 : _GEN_2611; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2613 = 8'h35 == io_state_in_2 ? 8'hd : _GEN_2612; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2614 = 8'h36 == io_state_in_2 ? 8'h1f : _GEN_2613; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2615 = 8'h37 == io_state_in_2 ? 8'h11 : _GEN_2614; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2616 = 8'h38 == io_state_in_2 ? 8'h4b : _GEN_2615; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2617 = 8'h39 == io_state_in_2 ? 8'h45 : _GEN_2616; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2618 = 8'h3a == io_state_in_2 ? 8'h57 : _GEN_2617; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2619 = 8'h3b == io_state_in_2 ? 8'h59 : _GEN_2618; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2620 = 8'h3c == io_state_in_2 ? 8'h73 : _GEN_2619; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2621 = 8'h3d == io_state_in_2 ? 8'h7d : _GEN_2620; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2622 = 8'h3e == io_state_in_2 ? 8'h6f : _GEN_2621; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2623 = 8'h3f == io_state_in_2 ? 8'h61 : _GEN_2622; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2624 = 8'h40 == io_state_in_2 ? 8'had : _GEN_2623; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2625 = 8'h41 == io_state_in_2 ? 8'ha3 : _GEN_2624; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2626 = 8'h42 == io_state_in_2 ? 8'hb1 : _GEN_2625; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2627 = 8'h43 == io_state_in_2 ? 8'hbf : _GEN_2626; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2628 = 8'h44 == io_state_in_2 ? 8'h95 : _GEN_2627; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2629 = 8'h45 == io_state_in_2 ? 8'h9b : _GEN_2628; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2630 = 8'h46 == io_state_in_2 ? 8'h89 : _GEN_2629; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2631 = 8'h47 == io_state_in_2 ? 8'h87 : _GEN_2630; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2632 = 8'h48 == io_state_in_2 ? 8'hdd : _GEN_2631; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2633 = 8'h49 == io_state_in_2 ? 8'hd3 : _GEN_2632; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2634 = 8'h4a == io_state_in_2 ? 8'hc1 : _GEN_2633; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2635 = 8'h4b == io_state_in_2 ? 8'hcf : _GEN_2634; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2636 = 8'h4c == io_state_in_2 ? 8'he5 : _GEN_2635; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2637 = 8'h4d == io_state_in_2 ? 8'heb : _GEN_2636; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2638 = 8'h4e == io_state_in_2 ? 8'hf9 : _GEN_2637; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2639 = 8'h4f == io_state_in_2 ? 8'hf7 : _GEN_2638; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2640 = 8'h50 == io_state_in_2 ? 8'h4d : _GEN_2639; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2641 = 8'h51 == io_state_in_2 ? 8'h43 : _GEN_2640; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2642 = 8'h52 == io_state_in_2 ? 8'h51 : _GEN_2641; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2643 = 8'h53 == io_state_in_2 ? 8'h5f : _GEN_2642; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2644 = 8'h54 == io_state_in_2 ? 8'h75 : _GEN_2643; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2645 = 8'h55 == io_state_in_2 ? 8'h7b : _GEN_2644; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2646 = 8'h56 == io_state_in_2 ? 8'h69 : _GEN_2645; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2647 = 8'h57 == io_state_in_2 ? 8'h67 : _GEN_2646; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2648 = 8'h58 == io_state_in_2 ? 8'h3d : _GEN_2647; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2649 = 8'h59 == io_state_in_2 ? 8'h33 : _GEN_2648; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2650 = 8'h5a == io_state_in_2 ? 8'h21 : _GEN_2649; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2651 = 8'h5b == io_state_in_2 ? 8'h2f : _GEN_2650; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2652 = 8'h5c == io_state_in_2 ? 8'h5 : _GEN_2651; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2653 = 8'h5d == io_state_in_2 ? 8'hb : _GEN_2652; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2654 = 8'h5e == io_state_in_2 ? 8'h19 : _GEN_2653; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2655 = 8'h5f == io_state_in_2 ? 8'h17 : _GEN_2654; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2656 = 8'h60 == io_state_in_2 ? 8'h76 : _GEN_2655; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2657 = 8'h61 == io_state_in_2 ? 8'h78 : _GEN_2656; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2658 = 8'h62 == io_state_in_2 ? 8'h6a : _GEN_2657; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2659 = 8'h63 == io_state_in_2 ? 8'h64 : _GEN_2658; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2660 = 8'h64 == io_state_in_2 ? 8'h4e : _GEN_2659; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2661 = 8'h65 == io_state_in_2 ? 8'h40 : _GEN_2660; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2662 = 8'h66 == io_state_in_2 ? 8'h52 : _GEN_2661; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2663 = 8'h67 == io_state_in_2 ? 8'h5c : _GEN_2662; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2664 = 8'h68 == io_state_in_2 ? 8'h6 : _GEN_2663; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2665 = 8'h69 == io_state_in_2 ? 8'h8 : _GEN_2664; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2666 = 8'h6a == io_state_in_2 ? 8'h1a : _GEN_2665; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2667 = 8'h6b == io_state_in_2 ? 8'h14 : _GEN_2666; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2668 = 8'h6c == io_state_in_2 ? 8'h3e : _GEN_2667; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2669 = 8'h6d == io_state_in_2 ? 8'h30 : _GEN_2668; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2670 = 8'h6e == io_state_in_2 ? 8'h22 : _GEN_2669; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2671 = 8'h6f == io_state_in_2 ? 8'h2c : _GEN_2670; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2672 = 8'h70 == io_state_in_2 ? 8'h96 : _GEN_2671; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2673 = 8'h71 == io_state_in_2 ? 8'h98 : _GEN_2672; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2674 = 8'h72 == io_state_in_2 ? 8'h8a : _GEN_2673; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2675 = 8'h73 == io_state_in_2 ? 8'h84 : _GEN_2674; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2676 = 8'h74 == io_state_in_2 ? 8'hae : _GEN_2675; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2677 = 8'h75 == io_state_in_2 ? 8'ha0 : _GEN_2676; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2678 = 8'h76 == io_state_in_2 ? 8'hb2 : _GEN_2677; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2679 = 8'h77 == io_state_in_2 ? 8'hbc : _GEN_2678; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2680 = 8'h78 == io_state_in_2 ? 8'he6 : _GEN_2679; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2681 = 8'h79 == io_state_in_2 ? 8'he8 : _GEN_2680; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2682 = 8'h7a == io_state_in_2 ? 8'hfa : _GEN_2681; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2683 = 8'h7b == io_state_in_2 ? 8'hf4 : _GEN_2682; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2684 = 8'h7c == io_state_in_2 ? 8'hde : _GEN_2683; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2685 = 8'h7d == io_state_in_2 ? 8'hd0 : _GEN_2684; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2686 = 8'h7e == io_state_in_2 ? 8'hc2 : _GEN_2685; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2687 = 8'h7f == io_state_in_2 ? 8'hcc : _GEN_2686; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2688 = 8'h80 == io_state_in_2 ? 8'h41 : _GEN_2687; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2689 = 8'h81 == io_state_in_2 ? 8'h4f : _GEN_2688; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2690 = 8'h82 == io_state_in_2 ? 8'h5d : _GEN_2689; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2691 = 8'h83 == io_state_in_2 ? 8'h53 : _GEN_2690; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2692 = 8'h84 == io_state_in_2 ? 8'h79 : _GEN_2691; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2693 = 8'h85 == io_state_in_2 ? 8'h77 : _GEN_2692; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2694 = 8'h86 == io_state_in_2 ? 8'h65 : _GEN_2693; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2695 = 8'h87 == io_state_in_2 ? 8'h6b : _GEN_2694; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2696 = 8'h88 == io_state_in_2 ? 8'h31 : _GEN_2695; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2697 = 8'h89 == io_state_in_2 ? 8'h3f : _GEN_2696; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2698 = 8'h8a == io_state_in_2 ? 8'h2d : _GEN_2697; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2699 = 8'h8b == io_state_in_2 ? 8'h23 : _GEN_2698; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2700 = 8'h8c == io_state_in_2 ? 8'h9 : _GEN_2699; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2701 = 8'h8d == io_state_in_2 ? 8'h7 : _GEN_2700; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2702 = 8'h8e == io_state_in_2 ? 8'h15 : _GEN_2701; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2703 = 8'h8f == io_state_in_2 ? 8'h1b : _GEN_2702; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2704 = 8'h90 == io_state_in_2 ? 8'ha1 : _GEN_2703; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2705 = 8'h91 == io_state_in_2 ? 8'haf : _GEN_2704; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2706 = 8'h92 == io_state_in_2 ? 8'hbd : _GEN_2705; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2707 = 8'h93 == io_state_in_2 ? 8'hb3 : _GEN_2706; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2708 = 8'h94 == io_state_in_2 ? 8'h99 : _GEN_2707; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2709 = 8'h95 == io_state_in_2 ? 8'h97 : _GEN_2708; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2710 = 8'h96 == io_state_in_2 ? 8'h85 : _GEN_2709; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2711 = 8'h97 == io_state_in_2 ? 8'h8b : _GEN_2710; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2712 = 8'h98 == io_state_in_2 ? 8'hd1 : _GEN_2711; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2713 = 8'h99 == io_state_in_2 ? 8'hdf : _GEN_2712; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2714 = 8'h9a == io_state_in_2 ? 8'hcd : _GEN_2713; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2715 = 8'h9b == io_state_in_2 ? 8'hc3 : _GEN_2714; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2716 = 8'h9c == io_state_in_2 ? 8'he9 : _GEN_2715; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2717 = 8'h9d == io_state_in_2 ? 8'he7 : _GEN_2716; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2718 = 8'h9e == io_state_in_2 ? 8'hf5 : _GEN_2717; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2719 = 8'h9f == io_state_in_2 ? 8'hfb : _GEN_2718; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2720 = 8'ha0 == io_state_in_2 ? 8'h9a : _GEN_2719; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2721 = 8'ha1 == io_state_in_2 ? 8'h94 : _GEN_2720; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2722 = 8'ha2 == io_state_in_2 ? 8'h86 : _GEN_2721; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2723 = 8'ha3 == io_state_in_2 ? 8'h88 : _GEN_2722; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2724 = 8'ha4 == io_state_in_2 ? 8'ha2 : _GEN_2723; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2725 = 8'ha5 == io_state_in_2 ? 8'hac : _GEN_2724; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2726 = 8'ha6 == io_state_in_2 ? 8'hbe : _GEN_2725; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2727 = 8'ha7 == io_state_in_2 ? 8'hb0 : _GEN_2726; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2728 = 8'ha8 == io_state_in_2 ? 8'hea : _GEN_2727; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2729 = 8'ha9 == io_state_in_2 ? 8'he4 : _GEN_2728; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2730 = 8'haa == io_state_in_2 ? 8'hf6 : _GEN_2729; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2731 = 8'hab == io_state_in_2 ? 8'hf8 : _GEN_2730; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2732 = 8'hac == io_state_in_2 ? 8'hd2 : _GEN_2731; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2733 = 8'had == io_state_in_2 ? 8'hdc : _GEN_2732; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2734 = 8'hae == io_state_in_2 ? 8'hce : _GEN_2733; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2735 = 8'haf == io_state_in_2 ? 8'hc0 : _GEN_2734; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2736 = 8'hb0 == io_state_in_2 ? 8'h7a : _GEN_2735; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2737 = 8'hb1 == io_state_in_2 ? 8'h74 : _GEN_2736; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2738 = 8'hb2 == io_state_in_2 ? 8'h66 : _GEN_2737; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2739 = 8'hb3 == io_state_in_2 ? 8'h68 : _GEN_2738; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2740 = 8'hb4 == io_state_in_2 ? 8'h42 : _GEN_2739; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2741 = 8'hb5 == io_state_in_2 ? 8'h4c : _GEN_2740; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2742 = 8'hb6 == io_state_in_2 ? 8'h5e : _GEN_2741; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2743 = 8'hb7 == io_state_in_2 ? 8'h50 : _GEN_2742; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2744 = 8'hb8 == io_state_in_2 ? 8'ha : _GEN_2743; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2745 = 8'hb9 == io_state_in_2 ? 8'h4 : _GEN_2744; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2746 = 8'hba == io_state_in_2 ? 8'h16 : _GEN_2745; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2747 = 8'hbb == io_state_in_2 ? 8'h18 : _GEN_2746; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2748 = 8'hbc == io_state_in_2 ? 8'h32 : _GEN_2747; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2749 = 8'hbd == io_state_in_2 ? 8'h3c : _GEN_2748; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2750 = 8'hbe == io_state_in_2 ? 8'h2e : _GEN_2749; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2751 = 8'hbf == io_state_in_2 ? 8'h20 : _GEN_2750; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2752 = 8'hc0 == io_state_in_2 ? 8'hec : _GEN_2751; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2753 = 8'hc1 == io_state_in_2 ? 8'he2 : _GEN_2752; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2754 = 8'hc2 == io_state_in_2 ? 8'hf0 : _GEN_2753; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2755 = 8'hc3 == io_state_in_2 ? 8'hfe : _GEN_2754; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2756 = 8'hc4 == io_state_in_2 ? 8'hd4 : _GEN_2755; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2757 = 8'hc5 == io_state_in_2 ? 8'hda : _GEN_2756; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2758 = 8'hc6 == io_state_in_2 ? 8'hc8 : _GEN_2757; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2759 = 8'hc7 == io_state_in_2 ? 8'hc6 : _GEN_2758; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2760 = 8'hc8 == io_state_in_2 ? 8'h9c : _GEN_2759; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2761 = 8'hc9 == io_state_in_2 ? 8'h92 : _GEN_2760; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2762 = 8'hca == io_state_in_2 ? 8'h80 : _GEN_2761; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2763 = 8'hcb == io_state_in_2 ? 8'h8e : _GEN_2762; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2764 = 8'hcc == io_state_in_2 ? 8'ha4 : _GEN_2763; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2765 = 8'hcd == io_state_in_2 ? 8'haa : _GEN_2764; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2766 = 8'hce == io_state_in_2 ? 8'hb8 : _GEN_2765; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2767 = 8'hcf == io_state_in_2 ? 8'hb6 : _GEN_2766; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2768 = 8'hd0 == io_state_in_2 ? 8'hc : _GEN_2767; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2769 = 8'hd1 == io_state_in_2 ? 8'h2 : _GEN_2768; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2770 = 8'hd2 == io_state_in_2 ? 8'h10 : _GEN_2769; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2771 = 8'hd3 == io_state_in_2 ? 8'h1e : _GEN_2770; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2772 = 8'hd4 == io_state_in_2 ? 8'h34 : _GEN_2771; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2773 = 8'hd5 == io_state_in_2 ? 8'h3a : _GEN_2772; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2774 = 8'hd6 == io_state_in_2 ? 8'h28 : _GEN_2773; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2775 = 8'hd7 == io_state_in_2 ? 8'h26 : _GEN_2774; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2776 = 8'hd8 == io_state_in_2 ? 8'h7c : _GEN_2775; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2777 = 8'hd9 == io_state_in_2 ? 8'h72 : _GEN_2776; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2778 = 8'hda == io_state_in_2 ? 8'h60 : _GEN_2777; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2779 = 8'hdb == io_state_in_2 ? 8'h6e : _GEN_2778; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2780 = 8'hdc == io_state_in_2 ? 8'h44 : _GEN_2779; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2781 = 8'hdd == io_state_in_2 ? 8'h4a : _GEN_2780; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2782 = 8'hde == io_state_in_2 ? 8'h58 : _GEN_2781; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2783 = 8'hdf == io_state_in_2 ? 8'h56 : _GEN_2782; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2784 = 8'he0 == io_state_in_2 ? 8'h37 : _GEN_2783; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2785 = 8'he1 == io_state_in_2 ? 8'h39 : _GEN_2784; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2786 = 8'he2 == io_state_in_2 ? 8'h2b : _GEN_2785; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2787 = 8'he3 == io_state_in_2 ? 8'h25 : _GEN_2786; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2788 = 8'he4 == io_state_in_2 ? 8'hf : _GEN_2787; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2789 = 8'he5 == io_state_in_2 ? 8'h1 : _GEN_2788; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2790 = 8'he6 == io_state_in_2 ? 8'h13 : _GEN_2789; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2791 = 8'he7 == io_state_in_2 ? 8'h1d : _GEN_2790; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2792 = 8'he8 == io_state_in_2 ? 8'h47 : _GEN_2791; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2793 = 8'he9 == io_state_in_2 ? 8'h49 : _GEN_2792; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2794 = 8'hea == io_state_in_2 ? 8'h5b : _GEN_2793; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2795 = 8'heb == io_state_in_2 ? 8'h55 : _GEN_2794; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2796 = 8'hec == io_state_in_2 ? 8'h7f : _GEN_2795; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2797 = 8'hed == io_state_in_2 ? 8'h71 : _GEN_2796; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2798 = 8'hee == io_state_in_2 ? 8'h63 : _GEN_2797; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2799 = 8'hef == io_state_in_2 ? 8'h6d : _GEN_2798; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2800 = 8'hf0 == io_state_in_2 ? 8'hd7 : _GEN_2799; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2801 = 8'hf1 == io_state_in_2 ? 8'hd9 : _GEN_2800; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2802 = 8'hf2 == io_state_in_2 ? 8'hcb : _GEN_2801; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2803 = 8'hf3 == io_state_in_2 ? 8'hc5 : _GEN_2802; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2804 = 8'hf4 == io_state_in_2 ? 8'hef : _GEN_2803; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2805 = 8'hf5 == io_state_in_2 ? 8'he1 : _GEN_2804; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2806 = 8'hf6 == io_state_in_2 ? 8'hf3 : _GEN_2805; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2807 = 8'hf7 == io_state_in_2 ? 8'hfd : _GEN_2806; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2808 = 8'hf8 == io_state_in_2 ? 8'ha7 : _GEN_2807; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2809 = 8'hf9 == io_state_in_2 ? 8'ha9 : _GEN_2808; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2810 = 8'hfa == io_state_in_2 ? 8'hbb : _GEN_2809; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2811 = 8'hfb == io_state_in_2 ? 8'hb5 : _GEN_2810; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2812 = 8'hfc == io_state_in_2 ? 8'h9f : _GEN_2811; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2813 = 8'hfd == io_state_in_2 ? 8'h91 : _GEN_2812; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2814 = 8'hfe == io_state_in_2 ? 8'h83 : _GEN_2813; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _GEN_2815 = 8'hff == io_state_in_2 ? 8'h8d : _GEN_2814; // @[InvMixColumns.scala 128:{65,65}]
  wire [7:0] _tmp_state_2_T_1 = _tmp_state_2_T ^ _GEN_2815; // @[InvMixColumns.scala 128:65]
  wire [7:0] _GEN_2817 = 8'h1 == io_state_in_3 ? 8'hb : 8'h0; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2818 = 8'h2 == io_state_in_3 ? 8'h16 : _GEN_2817; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2819 = 8'h3 == io_state_in_3 ? 8'h1d : _GEN_2818; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2820 = 8'h4 == io_state_in_3 ? 8'h2c : _GEN_2819; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2821 = 8'h5 == io_state_in_3 ? 8'h27 : _GEN_2820; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2822 = 8'h6 == io_state_in_3 ? 8'h3a : _GEN_2821; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2823 = 8'h7 == io_state_in_3 ? 8'h31 : _GEN_2822; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2824 = 8'h8 == io_state_in_3 ? 8'h58 : _GEN_2823; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2825 = 8'h9 == io_state_in_3 ? 8'h53 : _GEN_2824; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2826 = 8'ha == io_state_in_3 ? 8'h4e : _GEN_2825; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2827 = 8'hb == io_state_in_3 ? 8'h45 : _GEN_2826; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2828 = 8'hc == io_state_in_3 ? 8'h74 : _GEN_2827; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2829 = 8'hd == io_state_in_3 ? 8'h7f : _GEN_2828; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2830 = 8'he == io_state_in_3 ? 8'h62 : _GEN_2829; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2831 = 8'hf == io_state_in_3 ? 8'h69 : _GEN_2830; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2832 = 8'h10 == io_state_in_3 ? 8'hb0 : _GEN_2831; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2833 = 8'h11 == io_state_in_3 ? 8'hbb : _GEN_2832; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2834 = 8'h12 == io_state_in_3 ? 8'ha6 : _GEN_2833; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2835 = 8'h13 == io_state_in_3 ? 8'had : _GEN_2834; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2836 = 8'h14 == io_state_in_3 ? 8'h9c : _GEN_2835; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2837 = 8'h15 == io_state_in_3 ? 8'h97 : _GEN_2836; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2838 = 8'h16 == io_state_in_3 ? 8'h8a : _GEN_2837; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2839 = 8'h17 == io_state_in_3 ? 8'h81 : _GEN_2838; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2840 = 8'h18 == io_state_in_3 ? 8'he8 : _GEN_2839; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2841 = 8'h19 == io_state_in_3 ? 8'he3 : _GEN_2840; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2842 = 8'h1a == io_state_in_3 ? 8'hfe : _GEN_2841; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2843 = 8'h1b == io_state_in_3 ? 8'hf5 : _GEN_2842; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2844 = 8'h1c == io_state_in_3 ? 8'hc4 : _GEN_2843; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2845 = 8'h1d == io_state_in_3 ? 8'hcf : _GEN_2844; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2846 = 8'h1e == io_state_in_3 ? 8'hd2 : _GEN_2845; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2847 = 8'h1f == io_state_in_3 ? 8'hd9 : _GEN_2846; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2848 = 8'h20 == io_state_in_3 ? 8'h7b : _GEN_2847; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2849 = 8'h21 == io_state_in_3 ? 8'h70 : _GEN_2848; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2850 = 8'h22 == io_state_in_3 ? 8'h6d : _GEN_2849; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2851 = 8'h23 == io_state_in_3 ? 8'h66 : _GEN_2850; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2852 = 8'h24 == io_state_in_3 ? 8'h57 : _GEN_2851; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2853 = 8'h25 == io_state_in_3 ? 8'h5c : _GEN_2852; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2854 = 8'h26 == io_state_in_3 ? 8'h41 : _GEN_2853; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2855 = 8'h27 == io_state_in_3 ? 8'h4a : _GEN_2854; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2856 = 8'h28 == io_state_in_3 ? 8'h23 : _GEN_2855; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2857 = 8'h29 == io_state_in_3 ? 8'h28 : _GEN_2856; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2858 = 8'h2a == io_state_in_3 ? 8'h35 : _GEN_2857; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2859 = 8'h2b == io_state_in_3 ? 8'h3e : _GEN_2858; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2860 = 8'h2c == io_state_in_3 ? 8'hf : _GEN_2859; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2861 = 8'h2d == io_state_in_3 ? 8'h4 : _GEN_2860; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2862 = 8'h2e == io_state_in_3 ? 8'h19 : _GEN_2861; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2863 = 8'h2f == io_state_in_3 ? 8'h12 : _GEN_2862; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2864 = 8'h30 == io_state_in_3 ? 8'hcb : _GEN_2863; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2865 = 8'h31 == io_state_in_3 ? 8'hc0 : _GEN_2864; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2866 = 8'h32 == io_state_in_3 ? 8'hdd : _GEN_2865; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2867 = 8'h33 == io_state_in_3 ? 8'hd6 : _GEN_2866; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2868 = 8'h34 == io_state_in_3 ? 8'he7 : _GEN_2867; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2869 = 8'h35 == io_state_in_3 ? 8'hec : _GEN_2868; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2870 = 8'h36 == io_state_in_3 ? 8'hf1 : _GEN_2869; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2871 = 8'h37 == io_state_in_3 ? 8'hfa : _GEN_2870; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2872 = 8'h38 == io_state_in_3 ? 8'h93 : _GEN_2871; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2873 = 8'h39 == io_state_in_3 ? 8'h98 : _GEN_2872; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2874 = 8'h3a == io_state_in_3 ? 8'h85 : _GEN_2873; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2875 = 8'h3b == io_state_in_3 ? 8'h8e : _GEN_2874; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2876 = 8'h3c == io_state_in_3 ? 8'hbf : _GEN_2875; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2877 = 8'h3d == io_state_in_3 ? 8'hb4 : _GEN_2876; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2878 = 8'h3e == io_state_in_3 ? 8'ha9 : _GEN_2877; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2879 = 8'h3f == io_state_in_3 ? 8'ha2 : _GEN_2878; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2880 = 8'h40 == io_state_in_3 ? 8'hf6 : _GEN_2879; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2881 = 8'h41 == io_state_in_3 ? 8'hfd : _GEN_2880; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2882 = 8'h42 == io_state_in_3 ? 8'he0 : _GEN_2881; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2883 = 8'h43 == io_state_in_3 ? 8'heb : _GEN_2882; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2884 = 8'h44 == io_state_in_3 ? 8'hda : _GEN_2883; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2885 = 8'h45 == io_state_in_3 ? 8'hd1 : _GEN_2884; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2886 = 8'h46 == io_state_in_3 ? 8'hcc : _GEN_2885; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2887 = 8'h47 == io_state_in_3 ? 8'hc7 : _GEN_2886; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2888 = 8'h48 == io_state_in_3 ? 8'hae : _GEN_2887; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2889 = 8'h49 == io_state_in_3 ? 8'ha5 : _GEN_2888; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2890 = 8'h4a == io_state_in_3 ? 8'hb8 : _GEN_2889; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2891 = 8'h4b == io_state_in_3 ? 8'hb3 : _GEN_2890; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2892 = 8'h4c == io_state_in_3 ? 8'h82 : _GEN_2891; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2893 = 8'h4d == io_state_in_3 ? 8'h89 : _GEN_2892; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2894 = 8'h4e == io_state_in_3 ? 8'h94 : _GEN_2893; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2895 = 8'h4f == io_state_in_3 ? 8'h9f : _GEN_2894; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2896 = 8'h50 == io_state_in_3 ? 8'h46 : _GEN_2895; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2897 = 8'h51 == io_state_in_3 ? 8'h4d : _GEN_2896; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2898 = 8'h52 == io_state_in_3 ? 8'h50 : _GEN_2897; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2899 = 8'h53 == io_state_in_3 ? 8'h5b : _GEN_2898; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2900 = 8'h54 == io_state_in_3 ? 8'h6a : _GEN_2899; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2901 = 8'h55 == io_state_in_3 ? 8'h61 : _GEN_2900; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2902 = 8'h56 == io_state_in_3 ? 8'h7c : _GEN_2901; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2903 = 8'h57 == io_state_in_3 ? 8'h77 : _GEN_2902; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2904 = 8'h58 == io_state_in_3 ? 8'h1e : _GEN_2903; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2905 = 8'h59 == io_state_in_3 ? 8'h15 : _GEN_2904; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2906 = 8'h5a == io_state_in_3 ? 8'h8 : _GEN_2905; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2907 = 8'h5b == io_state_in_3 ? 8'h3 : _GEN_2906; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2908 = 8'h5c == io_state_in_3 ? 8'h32 : _GEN_2907; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2909 = 8'h5d == io_state_in_3 ? 8'h39 : _GEN_2908; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2910 = 8'h5e == io_state_in_3 ? 8'h24 : _GEN_2909; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2911 = 8'h5f == io_state_in_3 ? 8'h2f : _GEN_2910; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2912 = 8'h60 == io_state_in_3 ? 8'h8d : _GEN_2911; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2913 = 8'h61 == io_state_in_3 ? 8'h86 : _GEN_2912; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2914 = 8'h62 == io_state_in_3 ? 8'h9b : _GEN_2913; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2915 = 8'h63 == io_state_in_3 ? 8'h90 : _GEN_2914; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2916 = 8'h64 == io_state_in_3 ? 8'ha1 : _GEN_2915; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2917 = 8'h65 == io_state_in_3 ? 8'haa : _GEN_2916; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2918 = 8'h66 == io_state_in_3 ? 8'hb7 : _GEN_2917; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2919 = 8'h67 == io_state_in_3 ? 8'hbc : _GEN_2918; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2920 = 8'h68 == io_state_in_3 ? 8'hd5 : _GEN_2919; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2921 = 8'h69 == io_state_in_3 ? 8'hde : _GEN_2920; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2922 = 8'h6a == io_state_in_3 ? 8'hc3 : _GEN_2921; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2923 = 8'h6b == io_state_in_3 ? 8'hc8 : _GEN_2922; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2924 = 8'h6c == io_state_in_3 ? 8'hf9 : _GEN_2923; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2925 = 8'h6d == io_state_in_3 ? 8'hf2 : _GEN_2924; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2926 = 8'h6e == io_state_in_3 ? 8'hef : _GEN_2925; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2927 = 8'h6f == io_state_in_3 ? 8'he4 : _GEN_2926; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2928 = 8'h70 == io_state_in_3 ? 8'h3d : _GEN_2927; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2929 = 8'h71 == io_state_in_3 ? 8'h36 : _GEN_2928; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2930 = 8'h72 == io_state_in_3 ? 8'h2b : _GEN_2929; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2931 = 8'h73 == io_state_in_3 ? 8'h20 : _GEN_2930; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2932 = 8'h74 == io_state_in_3 ? 8'h11 : _GEN_2931; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2933 = 8'h75 == io_state_in_3 ? 8'h1a : _GEN_2932; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2934 = 8'h76 == io_state_in_3 ? 8'h7 : _GEN_2933; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2935 = 8'h77 == io_state_in_3 ? 8'hc : _GEN_2934; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2936 = 8'h78 == io_state_in_3 ? 8'h65 : _GEN_2935; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2937 = 8'h79 == io_state_in_3 ? 8'h6e : _GEN_2936; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2938 = 8'h7a == io_state_in_3 ? 8'h73 : _GEN_2937; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2939 = 8'h7b == io_state_in_3 ? 8'h78 : _GEN_2938; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2940 = 8'h7c == io_state_in_3 ? 8'h49 : _GEN_2939; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2941 = 8'h7d == io_state_in_3 ? 8'h42 : _GEN_2940; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2942 = 8'h7e == io_state_in_3 ? 8'h5f : _GEN_2941; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2943 = 8'h7f == io_state_in_3 ? 8'h54 : _GEN_2942; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2944 = 8'h80 == io_state_in_3 ? 8'hf7 : _GEN_2943; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2945 = 8'h81 == io_state_in_3 ? 8'hfc : _GEN_2944; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2946 = 8'h82 == io_state_in_3 ? 8'he1 : _GEN_2945; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2947 = 8'h83 == io_state_in_3 ? 8'hea : _GEN_2946; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2948 = 8'h84 == io_state_in_3 ? 8'hdb : _GEN_2947; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2949 = 8'h85 == io_state_in_3 ? 8'hd0 : _GEN_2948; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2950 = 8'h86 == io_state_in_3 ? 8'hcd : _GEN_2949; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2951 = 8'h87 == io_state_in_3 ? 8'hc6 : _GEN_2950; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2952 = 8'h88 == io_state_in_3 ? 8'haf : _GEN_2951; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2953 = 8'h89 == io_state_in_3 ? 8'ha4 : _GEN_2952; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2954 = 8'h8a == io_state_in_3 ? 8'hb9 : _GEN_2953; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2955 = 8'h8b == io_state_in_3 ? 8'hb2 : _GEN_2954; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2956 = 8'h8c == io_state_in_3 ? 8'h83 : _GEN_2955; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2957 = 8'h8d == io_state_in_3 ? 8'h88 : _GEN_2956; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2958 = 8'h8e == io_state_in_3 ? 8'h95 : _GEN_2957; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2959 = 8'h8f == io_state_in_3 ? 8'h9e : _GEN_2958; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2960 = 8'h90 == io_state_in_3 ? 8'h47 : _GEN_2959; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2961 = 8'h91 == io_state_in_3 ? 8'h4c : _GEN_2960; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2962 = 8'h92 == io_state_in_3 ? 8'h51 : _GEN_2961; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2963 = 8'h93 == io_state_in_3 ? 8'h5a : _GEN_2962; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2964 = 8'h94 == io_state_in_3 ? 8'h6b : _GEN_2963; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2965 = 8'h95 == io_state_in_3 ? 8'h60 : _GEN_2964; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2966 = 8'h96 == io_state_in_3 ? 8'h7d : _GEN_2965; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2967 = 8'h97 == io_state_in_3 ? 8'h76 : _GEN_2966; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2968 = 8'h98 == io_state_in_3 ? 8'h1f : _GEN_2967; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2969 = 8'h99 == io_state_in_3 ? 8'h14 : _GEN_2968; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2970 = 8'h9a == io_state_in_3 ? 8'h9 : _GEN_2969; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2971 = 8'h9b == io_state_in_3 ? 8'h2 : _GEN_2970; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2972 = 8'h9c == io_state_in_3 ? 8'h33 : _GEN_2971; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2973 = 8'h9d == io_state_in_3 ? 8'h38 : _GEN_2972; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2974 = 8'h9e == io_state_in_3 ? 8'h25 : _GEN_2973; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2975 = 8'h9f == io_state_in_3 ? 8'h2e : _GEN_2974; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2976 = 8'ha0 == io_state_in_3 ? 8'h8c : _GEN_2975; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2977 = 8'ha1 == io_state_in_3 ? 8'h87 : _GEN_2976; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2978 = 8'ha2 == io_state_in_3 ? 8'h9a : _GEN_2977; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2979 = 8'ha3 == io_state_in_3 ? 8'h91 : _GEN_2978; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2980 = 8'ha4 == io_state_in_3 ? 8'ha0 : _GEN_2979; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2981 = 8'ha5 == io_state_in_3 ? 8'hab : _GEN_2980; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2982 = 8'ha6 == io_state_in_3 ? 8'hb6 : _GEN_2981; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2983 = 8'ha7 == io_state_in_3 ? 8'hbd : _GEN_2982; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2984 = 8'ha8 == io_state_in_3 ? 8'hd4 : _GEN_2983; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2985 = 8'ha9 == io_state_in_3 ? 8'hdf : _GEN_2984; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2986 = 8'haa == io_state_in_3 ? 8'hc2 : _GEN_2985; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2987 = 8'hab == io_state_in_3 ? 8'hc9 : _GEN_2986; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2988 = 8'hac == io_state_in_3 ? 8'hf8 : _GEN_2987; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2989 = 8'had == io_state_in_3 ? 8'hf3 : _GEN_2988; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2990 = 8'hae == io_state_in_3 ? 8'hee : _GEN_2989; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2991 = 8'haf == io_state_in_3 ? 8'he5 : _GEN_2990; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2992 = 8'hb0 == io_state_in_3 ? 8'h3c : _GEN_2991; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2993 = 8'hb1 == io_state_in_3 ? 8'h37 : _GEN_2992; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2994 = 8'hb2 == io_state_in_3 ? 8'h2a : _GEN_2993; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2995 = 8'hb3 == io_state_in_3 ? 8'h21 : _GEN_2994; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2996 = 8'hb4 == io_state_in_3 ? 8'h10 : _GEN_2995; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2997 = 8'hb5 == io_state_in_3 ? 8'h1b : _GEN_2996; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2998 = 8'hb6 == io_state_in_3 ? 8'h6 : _GEN_2997; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_2999 = 8'hb7 == io_state_in_3 ? 8'hd : _GEN_2998; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3000 = 8'hb8 == io_state_in_3 ? 8'h64 : _GEN_2999; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3001 = 8'hb9 == io_state_in_3 ? 8'h6f : _GEN_3000; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3002 = 8'hba == io_state_in_3 ? 8'h72 : _GEN_3001; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3003 = 8'hbb == io_state_in_3 ? 8'h79 : _GEN_3002; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3004 = 8'hbc == io_state_in_3 ? 8'h48 : _GEN_3003; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3005 = 8'hbd == io_state_in_3 ? 8'h43 : _GEN_3004; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3006 = 8'hbe == io_state_in_3 ? 8'h5e : _GEN_3005; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3007 = 8'hbf == io_state_in_3 ? 8'h55 : _GEN_3006; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3008 = 8'hc0 == io_state_in_3 ? 8'h1 : _GEN_3007; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3009 = 8'hc1 == io_state_in_3 ? 8'ha : _GEN_3008; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3010 = 8'hc2 == io_state_in_3 ? 8'h17 : _GEN_3009; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3011 = 8'hc3 == io_state_in_3 ? 8'h1c : _GEN_3010; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3012 = 8'hc4 == io_state_in_3 ? 8'h2d : _GEN_3011; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3013 = 8'hc5 == io_state_in_3 ? 8'h26 : _GEN_3012; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3014 = 8'hc6 == io_state_in_3 ? 8'h3b : _GEN_3013; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3015 = 8'hc7 == io_state_in_3 ? 8'h30 : _GEN_3014; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3016 = 8'hc8 == io_state_in_3 ? 8'h59 : _GEN_3015; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3017 = 8'hc9 == io_state_in_3 ? 8'h52 : _GEN_3016; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3018 = 8'hca == io_state_in_3 ? 8'h4f : _GEN_3017; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3019 = 8'hcb == io_state_in_3 ? 8'h44 : _GEN_3018; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3020 = 8'hcc == io_state_in_3 ? 8'h75 : _GEN_3019; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3021 = 8'hcd == io_state_in_3 ? 8'h7e : _GEN_3020; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3022 = 8'hce == io_state_in_3 ? 8'h63 : _GEN_3021; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3023 = 8'hcf == io_state_in_3 ? 8'h68 : _GEN_3022; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3024 = 8'hd0 == io_state_in_3 ? 8'hb1 : _GEN_3023; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3025 = 8'hd1 == io_state_in_3 ? 8'hba : _GEN_3024; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3026 = 8'hd2 == io_state_in_3 ? 8'ha7 : _GEN_3025; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3027 = 8'hd3 == io_state_in_3 ? 8'hac : _GEN_3026; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3028 = 8'hd4 == io_state_in_3 ? 8'h9d : _GEN_3027; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3029 = 8'hd5 == io_state_in_3 ? 8'h96 : _GEN_3028; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3030 = 8'hd6 == io_state_in_3 ? 8'h8b : _GEN_3029; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3031 = 8'hd7 == io_state_in_3 ? 8'h80 : _GEN_3030; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3032 = 8'hd8 == io_state_in_3 ? 8'he9 : _GEN_3031; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3033 = 8'hd9 == io_state_in_3 ? 8'he2 : _GEN_3032; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3034 = 8'hda == io_state_in_3 ? 8'hff : _GEN_3033; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3035 = 8'hdb == io_state_in_3 ? 8'hf4 : _GEN_3034; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3036 = 8'hdc == io_state_in_3 ? 8'hc5 : _GEN_3035; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3037 = 8'hdd == io_state_in_3 ? 8'hce : _GEN_3036; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3038 = 8'hde == io_state_in_3 ? 8'hd3 : _GEN_3037; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3039 = 8'hdf == io_state_in_3 ? 8'hd8 : _GEN_3038; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3040 = 8'he0 == io_state_in_3 ? 8'h7a : _GEN_3039; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3041 = 8'he1 == io_state_in_3 ? 8'h71 : _GEN_3040; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3042 = 8'he2 == io_state_in_3 ? 8'h6c : _GEN_3041; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3043 = 8'he3 == io_state_in_3 ? 8'h67 : _GEN_3042; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3044 = 8'he4 == io_state_in_3 ? 8'h56 : _GEN_3043; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3045 = 8'he5 == io_state_in_3 ? 8'h5d : _GEN_3044; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3046 = 8'he6 == io_state_in_3 ? 8'h40 : _GEN_3045; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3047 = 8'he7 == io_state_in_3 ? 8'h4b : _GEN_3046; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3048 = 8'he8 == io_state_in_3 ? 8'h22 : _GEN_3047; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3049 = 8'he9 == io_state_in_3 ? 8'h29 : _GEN_3048; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3050 = 8'hea == io_state_in_3 ? 8'h34 : _GEN_3049; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3051 = 8'heb == io_state_in_3 ? 8'h3f : _GEN_3050; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3052 = 8'hec == io_state_in_3 ? 8'he : _GEN_3051; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3053 = 8'hed == io_state_in_3 ? 8'h5 : _GEN_3052; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3054 = 8'hee == io_state_in_3 ? 8'h18 : _GEN_3053; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3055 = 8'hef == io_state_in_3 ? 8'h13 : _GEN_3054; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3056 = 8'hf0 == io_state_in_3 ? 8'hca : _GEN_3055; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3057 = 8'hf1 == io_state_in_3 ? 8'hc1 : _GEN_3056; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3058 = 8'hf2 == io_state_in_3 ? 8'hdc : _GEN_3057; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3059 = 8'hf3 == io_state_in_3 ? 8'hd7 : _GEN_3058; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3060 = 8'hf4 == io_state_in_3 ? 8'he6 : _GEN_3059; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3061 = 8'hf5 == io_state_in_3 ? 8'hed : _GEN_3060; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3062 = 8'hf6 == io_state_in_3 ? 8'hf0 : _GEN_3061; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3063 = 8'hf7 == io_state_in_3 ? 8'hfb : _GEN_3062; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3064 = 8'hf8 == io_state_in_3 ? 8'h92 : _GEN_3063; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3065 = 8'hf9 == io_state_in_3 ? 8'h99 : _GEN_3064; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3066 = 8'hfa == io_state_in_3 ? 8'h84 : _GEN_3065; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3067 = 8'hfb == io_state_in_3 ? 8'h8f : _GEN_3066; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3068 = 8'hfc == io_state_in_3 ? 8'hbe : _GEN_3067; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3069 = 8'hfd == io_state_in_3 ? 8'hb5 : _GEN_3068; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3070 = 8'hfe == io_state_in_3 ? 8'ha8 : _GEN_3069; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3071 = 8'hff == io_state_in_3 ? 8'ha3 : _GEN_3070; // @[InvMixColumns.scala 128:{89,89}]
  wire [7:0] _GEN_3073 = 8'h1 == io_state_in_0 ? 8'hb : 8'h0; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3074 = 8'h2 == io_state_in_0 ? 8'h16 : _GEN_3073; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3075 = 8'h3 == io_state_in_0 ? 8'h1d : _GEN_3074; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3076 = 8'h4 == io_state_in_0 ? 8'h2c : _GEN_3075; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3077 = 8'h5 == io_state_in_0 ? 8'h27 : _GEN_3076; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3078 = 8'h6 == io_state_in_0 ? 8'h3a : _GEN_3077; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3079 = 8'h7 == io_state_in_0 ? 8'h31 : _GEN_3078; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3080 = 8'h8 == io_state_in_0 ? 8'h58 : _GEN_3079; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3081 = 8'h9 == io_state_in_0 ? 8'h53 : _GEN_3080; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3082 = 8'ha == io_state_in_0 ? 8'h4e : _GEN_3081; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3083 = 8'hb == io_state_in_0 ? 8'h45 : _GEN_3082; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3084 = 8'hc == io_state_in_0 ? 8'h74 : _GEN_3083; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3085 = 8'hd == io_state_in_0 ? 8'h7f : _GEN_3084; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3086 = 8'he == io_state_in_0 ? 8'h62 : _GEN_3085; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3087 = 8'hf == io_state_in_0 ? 8'h69 : _GEN_3086; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3088 = 8'h10 == io_state_in_0 ? 8'hb0 : _GEN_3087; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3089 = 8'h11 == io_state_in_0 ? 8'hbb : _GEN_3088; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3090 = 8'h12 == io_state_in_0 ? 8'ha6 : _GEN_3089; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3091 = 8'h13 == io_state_in_0 ? 8'had : _GEN_3090; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3092 = 8'h14 == io_state_in_0 ? 8'h9c : _GEN_3091; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3093 = 8'h15 == io_state_in_0 ? 8'h97 : _GEN_3092; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3094 = 8'h16 == io_state_in_0 ? 8'h8a : _GEN_3093; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3095 = 8'h17 == io_state_in_0 ? 8'h81 : _GEN_3094; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3096 = 8'h18 == io_state_in_0 ? 8'he8 : _GEN_3095; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3097 = 8'h19 == io_state_in_0 ? 8'he3 : _GEN_3096; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3098 = 8'h1a == io_state_in_0 ? 8'hfe : _GEN_3097; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3099 = 8'h1b == io_state_in_0 ? 8'hf5 : _GEN_3098; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3100 = 8'h1c == io_state_in_0 ? 8'hc4 : _GEN_3099; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3101 = 8'h1d == io_state_in_0 ? 8'hcf : _GEN_3100; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3102 = 8'h1e == io_state_in_0 ? 8'hd2 : _GEN_3101; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3103 = 8'h1f == io_state_in_0 ? 8'hd9 : _GEN_3102; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3104 = 8'h20 == io_state_in_0 ? 8'h7b : _GEN_3103; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3105 = 8'h21 == io_state_in_0 ? 8'h70 : _GEN_3104; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3106 = 8'h22 == io_state_in_0 ? 8'h6d : _GEN_3105; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3107 = 8'h23 == io_state_in_0 ? 8'h66 : _GEN_3106; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3108 = 8'h24 == io_state_in_0 ? 8'h57 : _GEN_3107; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3109 = 8'h25 == io_state_in_0 ? 8'h5c : _GEN_3108; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3110 = 8'h26 == io_state_in_0 ? 8'h41 : _GEN_3109; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3111 = 8'h27 == io_state_in_0 ? 8'h4a : _GEN_3110; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3112 = 8'h28 == io_state_in_0 ? 8'h23 : _GEN_3111; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3113 = 8'h29 == io_state_in_0 ? 8'h28 : _GEN_3112; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3114 = 8'h2a == io_state_in_0 ? 8'h35 : _GEN_3113; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3115 = 8'h2b == io_state_in_0 ? 8'h3e : _GEN_3114; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3116 = 8'h2c == io_state_in_0 ? 8'hf : _GEN_3115; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3117 = 8'h2d == io_state_in_0 ? 8'h4 : _GEN_3116; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3118 = 8'h2e == io_state_in_0 ? 8'h19 : _GEN_3117; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3119 = 8'h2f == io_state_in_0 ? 8'h12 : _GEN_3118; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3120 = 8'h30 == io_state_in_0 ? 8'hcb : _GEN_3119; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3121 = 8'h31 == io_state_in_0 ? 8'hc0 : _GEN_3120; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3122 = 8'h32 == io_state_in_0 ? 8'hdd : _GEN_3121; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3123 = 8'h33 == io_state_in_0 ? 8'hd6 : _GEN_3122; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3124 = 8'h34 == io_state_in_0 ? 8'he7 : _GEN_3123; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3125 = 8'h35 == io_state_in_0 ? 8'hec : _GEN_3124; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3126 = 8'h36 == io_state_in_0 ? 8'hf1 : _GEN_3125; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3127 = 8'h37 == io_state_in_0 ? 8'hfa : _GEN_3126; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3128 = 8'h38 == io_state_in_0 ? 8'h93 : _GEN_3127; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3129 = 8'h39 == io_state_in_0 ? 8'h98 : _GEN_3128; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3130 = 8'h3a == io_state_in_0 ? 8'h85 : _GEN_3129; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3131 = 8'h3b == io_state_in_0 ? 8'h8e : _GEN_3130; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3132 = 8'h3c == io_state_in_0 ? 8'hbf : _GEN_3131; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3133 = 8'h3d == io_state_in_0 ? 8'hb4 : _GEN_3132; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3134 = 8'h3e == io_state_in_0 ? 8'ha9 : _GEN_3133; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3135 = 8'h3f == io_state_in_0 ? 8'ha2 : _GEN_3134; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3136 = 8'h40 == io_state_in_0 ? 8'hf6 : _GEN_3135; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3137 = 8'h41 == io_state_in_0 ? 8'hfd : _GEN_3136; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3138 = 8'h42 == io_state_in_0 ? 8'he0 : _GEN_3137; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3139 = 8'h43 == io_state_in_0 ? 8'heb : _GEN_3138; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3140 = 8'h44 == io_state_in_0 ? 8'hda : _GEN_3139; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3141 = 8'h45 == io_state_in_0 ? 8'hd1 : _GEN_3140; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3142 = 8'h46 == io_state_in_0 ? 8'hcc : _GEN_3141; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3143 = 8'h47 == io_state_in_0 ? 8'hc7 : _GEN_3142; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3144 = 8'h48 == io_state_in_0 ? 8'hae : _GEN_3143; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3145 = 8'h49 == io_state_in_0 ? 8'ha5 : _GEN_3144; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3146 = 8'h4a == io_state_in_0 ? 8'hb8 : _GEN_3145; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3147 = 8'h4b == io_state_in_0 ? 8'hb3 : _GEN_3146; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3148 = 8'h4c == io_state_in_0 ? 8'h82 : _GEN_3147; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3149 = 8'h4d == io_state_in_0 ? 8'h89 : _GEN_3148; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3150 = 8'h4e == io_state_in_0 ? 8'h94 : _GEN_3149; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3151 = 8'h4f == io_state_in_0 ? 8'h9f : _GEN_3150; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3152 = 8'h50 == io_state_in_0 ? 8'h46 : _GEN_3151; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3153 = 8'h51 == io_state_in_0 ? 8'h4d : _GEN_3152; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3154 = 8'h52 == io_state_in_0 ? 8'h50 : _GEN_3153; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3155 = 8'h53 == io_state_in_0 ? 8'h5b : _GEN_3154; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3156 = 8'h54 == io_state_in_0 ? 8'h6a : _GEN_3155; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3157 = 8'h55 == io_state_in_0 ? 8'h61 : _GEN_3156; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3158 = 8'h56 == io_state_in_0 ? 8'h7c : _GEN_3157; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3159 = 8'h57 == io_state_in_0 ? 8'h77 : _GEN_3158; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3160 = 8'h58 == io_state_in_0 ? 8'h1e : _GEN_3159; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3161 = 8'h59 == io_state_in_0 ? 8'h15 : _GEN_3160; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3162 = 8'h5a == io_state_in_0 ? 8'h8 : _GEN_3161; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3163 = 8'h5b == io_state_in_0 ? 8'h3 : _GEN_3162; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3164 = 8'h5c == io_state_in_0 ? 8'h32 : _GEN_3163; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3165 = 8'h5d == io_state_in_0 ? 8'h39 : _GEN_3164; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3166 = 8'h5e == io_state_in_0 ? 8'h24 : _GEN_3165; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3167 = 8'h5f == io_state_in_0 ? 8'h2f : _GEN_3166; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3168 = 8'h60 == io_state_in_0 ? 8'h8d : _GEN_3167; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3169 = 8'h61 == io_state_in_0 ? 8'h86 : _GEN_3168; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3170 = 8'h62 == io_state_in_0 ? 8'h9b : _GEN_3169; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3171 = 8'h63 == io_state_in_0 ? 8'h90 : _GEN_3170; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3172 = 8'h64 == io_state_in_0 ? 8'ha1 : _GEN_3171; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3173 = 8'h65 == io_state_in_0 ? 8'haa : _GEN_3172; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3174 = 8'h66 == io_state_in_0 ? 8'hb7 : _GEN_3173; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3175 = 8'h67 == io_state_in_0 ? 8'hbc : _GEN_3174; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3176 = 8'h68 == io_state_in_0 ? 8'hd5 : _GEN_3175; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3177 = 8'h69 == io_state_in_0 ? 8'hde : _GEN_3176; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3178 = 8'h6a == io_state_in_0 ? 8'hc3 : _GEN_3177; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3179 = 8'h6b == io_state_in_0 ? 8'hc8 : _GEN_3178; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3180 = 8'h6c == io_state_in_0 ? 8'hf9 : _GEN_3179; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3181 = 8'h6d == io_state_in_0 ? 8'hf2 : _GEN_3180; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3182 = 8'h6e == io_state_in_0 ? 8'hef : _GEN_3181; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3183 = 8'h6f == io_state_in_0 ? 8'he4 : _GEN_3182; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3184 = 8'h70 == io_state_in_0 ? 8'h3d : _GEN_3183; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3185 = 8'h71 == io_state_in_0 ? 8'h36 : _GEN_3184; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3186 = 8'h72 == io_state_in_0 ? 8'h2b : _GEN_3185; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3187 = 8'h73 == io_state_in_0 ? 8'h20 : _GEN_3186; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3188 = 8'h74 == io_state_in_0 ? 8'h11 : _GEN_3187; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3189 = 8'h75 == io_state_in_0 ? 8'h1a : _GEN_3188; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3190 = 8'h76 == io_state_in_0 ? 8'h7 : _GEN_3189; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3191 = 8'h77 == io_state_in_0 ? 8'hc : _GEN_3190; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3192 = 8'h78 == io_state_in_0 ? 8'h65 : _GEN_3191; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3193 = 8'h79 == io_state_in_0 ? 8'h6e : _GEN_3192; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3194 = 8'h7a == io_state_in_0 ? 8'h73 : _GEN_3193; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3195 = 8'h7b == io_state_in_0 ? 8'h78 : _GEN_3194; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3196 = 8'h7c == io_state_in_0 ? 8'h49 : _GEN_3195; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3197 = 8'h7d == io_state_in_0 ? 8'h42 : _GEN_3196; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3198 = 8'h7e == io_state_in_0 ? 8'h5f : _GEN_3197; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3199 = 8'h7f == io_state_in_0 ? 8'h54 : _GEN_3198; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3200 = 8'h80 == io_state_in_0 ? 8'hf7 : _GEN_3199; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3201 = 8'h81 == io_state_in_0 ? 8'hfc : _GEN_3200; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3202 = 8'h82 == io_state_in_0 ? 8'he1 : _GEN_3201; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3203 = 8'h83 == io_state_in_0 ? 8'hea : _GEN_3202; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3204 = 8'h84 == io_state_in_0 ? 8'hdb : _GEN_3203; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3205 = 8'h85 == io_state_in_0 ? 8'hd0 : _GEN_3204; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3206 = 8'h86 == io_state_in_0 ? 8'hcd : _GEN_3205; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3207 = 8'h87 == io_state_in_0 ? 8'hc6 : _GEN_3206; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3208 = 8'h88 == io_state_in_0 ? 8'haf : _GEN_3207; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3209 = 8'h89 == io_state_in_0 ? 8'ha4 : _GEN_3208; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3210 = 8'h8a == io_state_in_0 ? 8'hb9 : _GEN_3209; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3211 = 8'h8b == io_state_in_0 ? 8'hb2 : _GEN_3210; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3212 = 8'h8c == io_state_in_0 ? 8'h83 : _GEN_3211; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3213 = 8'h8d == io_state_in_0 ? 8'h88 : _GEN_3212; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3214 = 8'h8e == io_state_in_0 ? 8'h95 : _GEN_3213; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3215 = 8'h8f == io_state_in_0 ? 8'h9e : _GEN_3214; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3216 = 8'h90 == io_state_in_0 ? 8'h47 : _GEN_3215; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3217 = 8'h91 == io_state_in_0 ? 8'h4c : _GEN_3216; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3218 = 8'h92 == io_state_in_0 ? 8'h51 : _GEN_3217; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3219 = 8'h93 == io_state_in_0 ? 8'h5a : _GEN_3218; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3220 = 8'h94 == io_state_in_0 ? 8'h6b : _GEN_3219; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3221 = 8'h95 == io_state_in_0 ? 8'h60 : _GEN_3220; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3222 = 8'h96 == io_state_in_0 ? 8'h7d : _GEN_3221; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3223 = 8'h97 == io_state_in_0 ? 8'h76 : _GEN_3222; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3224 = 8'h98 == io_state_in_0 ? 8'h1f : _GEN_3223; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3225 = 8'h99 == io_state_in_0 ? 8'h14 : _GEN_3224; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3226 = 8'h9a == io_state_in_0 ? 8'h9 : _GEN_3225; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3227 = 8'h9b == io_state_in_0 ? 8'h2 : _GEN_3226; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3228 = 8'h9c == io_state_in_0 ? 8'h33 : _GEN_3227; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3229 = 8'h9d == io_state_in_0 ? 8'h38 : _GEN_3228; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3230 = 8'h9e == io_state_in_0 ? 8'h25 : _GEN_3229; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3231 = 8'h9f == io_state_in_0 ? 8'h2e : _GEN_3230; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3232 = 8'ha0 == io_state_in_0 ? 8'h8c : _GEN_3231; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3233 = 8'ha1 == io_state_in_0 ? 8'h87 : _GEN_3232; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3234 = 8'ha2 == io_state_in_0 ? 8'h9a : _GEN_3233; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3235 = 8'ha3 == io_state_in_0 ? 8'h91 : _GEN_3234; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3236 = 8'ha4 == io_state_in_0 ? 8'ha0 : _GEN_3235; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3237 = 8'ha5 == io_state_in_0 ? 8'hab : _GEN_3236; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3238 = 8'ha6 == io_state_in_0 ? 8'hb6 : _GEN_3237; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3239 = 8'ha7 == io_state_in_0 ? 8'hbd : _GEN_3238; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3240 = 8'ha8 == io_state_in_0 ? 8'hd4 : _GEN_3239; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3241 = 8'ha9 == io_state_in_0 ? 8'hdf : _GEN_3240; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3242 = 8'haa == io_state_in_0 ? 8'hc2 : _GEN_3241; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3243 = 8'hab == io_state_in_0 ? 8'hc9 : _GEN_3242; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3244 = 8'hac == io_state_in_0 ? 8'hf8 : _GEN_3243; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3245 = 8'had == io_state_in_0 ? 8'hf3 : _GEN_3244; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3246 = 8'hae == io_state_in_0 ? 8'hee : _GEN_3245; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3247 = 8'haf == io_state_in_0 ? 8'he5 : _GEN_3246; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3248 = 8'hb0 == io_state_in_0 ? 8'h3c : _GEN_3247; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3249 = 8'hb1 == io_state_in_0 ? 8'h37 : _GEN_3248; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3250 = 8'hb2 == io_state_in_0 ? 8'h2a : _GEN_3249; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3251 = 8'hb3 == io_state_in_0 ? 8'h21 : _GEN_3250; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3252 = 8'hb4 == io_state_in_0 ? 8'h10 : _GEN_3251; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3253 = 8'hb5 == io_state_in_0 ? 8'h1b : _GEN_3252; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3254 = 8'hb6 == io_state_in_0 ? 8'h6 : _GEN_3253; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3255 = 8'hb7 == io_state_in_0 ? 8'hd : _GEN_3254; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3256 = 8'hb8 == io_state_in_0 ? 8'h64 : _GEN_3255; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3257 = 8'hb9 == io_state_in_0 ? 8'h6f : _GEN_3256; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3258 = 8'hba == io_state_in_0 ? 8'h72 : _GEN_3257; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3259 = 8'hbb == io_state_in_0 ? 8'h79 : _GEN_3258; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3260 = 8'hbc == io_state_in_0 ? 8'h48 : _GEN_3259; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3261 = 8'hbd == io_state_in_0 ? 8'h43 : _GEN_3260; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3262 = 8'hbe == io_state_in_0 ? 8'h5e : _GEN_3261; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3263 = 8'hbf == io_state_in_0 ? 8'h55 : _GEN_3262; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3264 = 8'hc0 == io_state_in_0 ? 8'h1 : _GEN_3263; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3265 = 8'hc1 == io_state_in_0 ? 8'ha : _GEN_3264; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3266 = 8'hc2 == io_state_in_0 ? 8'h17 : _GEN_3265; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3267 = 8'hc3 == io_state_in_0 ? 8'h1c : _GEN_3266; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3268 = 8'hc4 == io_state_in_0 ? 8'h2d : _GEN_3267; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3269 = 8'hc5 == io_state_in_0 ? 8'h26 : _GEN_3268; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3270 = 8'hc6 == io_state_in_0 ? 8'h3b : _GEN_3269; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3271 = 8'hc7 == io_state_in_0 ? 8'h30 : _GEN_3270; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3272 = 8'hc8 == io_state_in_0 ? 8'h59 : _GEN_3271; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3273 = 8'hc9 == io_state_in_0 ? 8'h52 : _GEN_3272; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3274 = 8'hca == io_state_in_0 ? 8'h4f : _GEN_3273; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3275 = 8'hcb == io_state_in_0 ? 8'h44 : _GEN_3274; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3276 = 8'hcc == io_state_in_0 ? 8'h75 : _GEN_3275; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3277 = 8'hcd == io_state_in_0 ? 8'h7e : _GEN_3276; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3278 = 8'hce == io_state_in_0 ? 8'h63 : _GEN_3277; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3279 = 8'hcf == io_state_in_0 ? 8'h68 : _GEN_3278; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3280 = 8'hd0 == io_state_in_0 ? 8'hb1 : _GEN_3279; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3281 = 8'hd1 == io_state_in_0 ? 8'hba : _GEN_3280; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3282 = 8'hd2 == io_state_in_0 ? 8'ha7 : _GEN_3281; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3283 = 8'hd3 == io_state_in_0 ? 8'hac : _GEN_3282; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3284 = 8'hd4 == io_state_in_0 ? 8'h9d : _GEN_3283; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3285 = 8'hd5 == io_state_in_0 ? 8'h96 : _GEN_3284; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3286 = 8'hd6 == io_state_in_0 ? 8'h8b : _GEN_3285; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3287 = 8'hd7 == io_state_in_0 ? 8'h80 : _GEN_3286; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3288 = 8'hd8 == io_state_in_0 ? 8'he9 : _GEN_3287; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3289 = 8'hd9 == io_state_in_0 ? 8'he2 : _GEN_3288; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3290 = 8'hda == io_state_in_0 ? 8'hff : _GEN_3289; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3291 = 8'hdb == io_state_in_0 ? 8'hf4 : _GEN_3290; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3292 = 8'hdc == io_state_in_0 ? 8'hc5 : _GEN_3291; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3293 = 8'hdd == io_state_in_0 ? 8'hce : _GEN_3292; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3294 = 8'hde == io_state_in_0 ? 8'hd3 : _GEN_3293; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3295 = 8'hdf == io_state_in_0 ? 8'hd8 : _GEN_3294; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3296 = 8'he0 == io_state_in_0 ? 8'h7a : _GEN_3295; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3297 = 8'he1 == io_state_in_0 ? 8'h71 : _GEN_3296; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3298 = 8'he2 == io_state_in_0 ? 8'h6c : _GEN_3297; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3299 = 8'he3 == io_state_in_0 ? 8'h67 : _GEN_3298; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3300 = 8'he4 == io_state_in_0 ? 8'h56 : _GEN_3299; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3301 = 8'he5 == io_state_in_0 ? 8'h5d : _GEN_3300; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3302 = 8'he6 == io_state_in_0 ? 8'h40 : _GEN_3301; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3303 = 8'he7 == io_state_in_0 ? 8'h4b : _GEN_3302; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3304 = 8'he8 == io_state_in_0 ? 8'h22 : _GEN_3303; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3305 = 8'he9 == io_state_in_0 ? 8'h29 : _GEN_3304; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3306 = 8'hea == io_state_in_0 ? 8'h34 : _GEN_3305; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3307 = 8'heb == io_state_in_0 ? 8'h3f : _GEN_3306; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3308 = 8'hec == io_state_in_0 ? 8'he : _GEN_3307; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3309 = 8'hed == io_state_in_0 ? 8'h5 : _GEN_3308; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3310 = 8'hee == io_state_in_0 ? 8'h18 : _GEN_3309; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3311 = 8'hef == io_state_in_0 ? 8'h13 : _GEN_3310; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3312 = 8'hf0 == io_state_in_0 ? 8'hca : _GEN_3311; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3313 = 8'hf1 == io_state_in_0 ? 8'hc1 : _GEN_3312; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3314 = 8'hf2 == io_state_in_0 ? 8'hdc : _GEN_3313; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3315 = 8'hf3 == io_state_in_0 ? 8'hd7 : _GEN_3314; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3316 = 8'hf4 == io_state_in_0 ? 8'he6 : _GEN_3315; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3317 = 8'hf5 == io_state_in_0 ? 8'hed : _GEN_3316; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3318 = 8'hf6 == io_state_in_0 ? 8'hf0 : _GEN_3317; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3319 = 8'hf7 == io_state_in_0 ? 8'hfb : _GEN_3318; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3320 = 8'hf8 == io_state_in_0 ? 8'h92 : _GEN_3319; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3321 = 8'hf9 == io_state_in_0 ? 8'h99 : _GEN_3320; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3322 = 8'hfa == io_state_in_0 ? 8'h84 : _GEN_3321; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3323 = 8'hfb == io_state_in_0 ? 8'h8f : _GEN_3322; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3324 = 8'hfc == io_state_in_0 ? 8'hbe : _GEN_3323; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3325 = 8'hfd == io_state_in_0 ? 8'hb5 : _GEN_3324; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3326 = 8'hfe == io_state_in_0 ? 8'ha8 : _GEN_3325; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3327 = 8'hff == io_state_in_0 ? 8'ha3 : _GEN_3326; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3329 = 8'h1 == io_state_in_1 ? 8'hd : 8'h0; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3330 = 8'h2 == io_state_in_1 ? 8'h1a : _GEN_3329; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3331 = 8'h3 == io_state_in_1 ? 8'h17 : _GEN_3330; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3332 = 8'h4 == io_state_in_1 ? 8'h34 : _GEN_3331; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3333 = 8'h5 == io_state_in_1 ? 8'h39 : _GEN_3332; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3334 = 8'h6 == io_state_in_1 ? 8'h2e : _GEN_3333; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3335 = 8'h7 == io_state_in_1 ? 8'h23 : _GEN_3334; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3336 = 8'h8 == io_state_in_1 ? 8'h68 : _GEN_3335; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3337 = 8'h9 == io_state_in_1 ? 8'h65 : _GEN_3336; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3338 = 8'ha == io_state_in_1 ? 8'h72 : _GEN_3337; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3339 = 8'hb == io_state_in_1 ? 8'h7f : _GEN_3338; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3340 = 8'hc == io_state_in_1 ? 8'h5c : _GEN_3339; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3341 = 8'hd == io_state_in_1 ? 8'h51 : _GEN_3340; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3342 = 8'he == io_state_in_1 ? 8'h46 : _GEN_3341; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3343 = 8'hf == io_state_in_1 ? 8'h4b : _GEN_3342; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3344 = 8'h10 == io_state_in_1 ? 8'hd0 : _GEN_3343; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3345 = 8'h11 == io_state_in_1 ? 8'hdd : _GEN_3344; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3346 = 8'h12 == io_state_in_1 ? 8'hca : _GEN_3345; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3347 = 8'h13 == io_state_in_1 ? 8'hc7 : _GEN_3346; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3348 = 8'h14 == io_state_in_1 ? 8'he4 : _GEN_3347; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3349 = 8'h15 == io_state_in_1 ? 8'he9 : _GEN_3348; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3350 = 8'h16 == io_state_in_1 ? 8'hfe : _GEN_3349; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3351 = 8'h17 == io_state_in_1 ? 8'hf3 : _GEN_3350; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3352 = 8'h18 == io_state_in_1 ? 8'hb8 : _GEN_3351; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3353 = 8'h19 == io_state_in_1 ? 8'hb5 : _GEN_3352; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3354 = 8'h1a == io_state_in_1 ? 8'ha2 : _GEN_3353; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3355 = 8'h1b == io_state_in_1 ? 8'haf : _GEN_3354; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3356 = 8'h1c == io_state_in_1 ? 8'h8c : _GEN_3355; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3357 = 8'h1d == io_state_in_1 ? 8'h81 : _GEN_3356; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3358 = 8'h1e == io_state_in_1 ? 8'h96 : _GEN_3357; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3359 = 8'h1f == io_state_in_1 ? 8'h9b : _GEN_3358; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3360 = 8'h20 == io_state_in_1 ? 8'hbb : _GEN_3359; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3361 = 8'h21 == io_state_in_1 ? 8'hb6 : _GEN_3360; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3362 = 8'h22 == io_state_in_1 ? 8'ha1 : _GEN_3361; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3363 = 8'h23 == io_state_in_1 ? 8'hac : _GEN_3362; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3364 = 8'h24 == io_state_in_1 ? 8'h8f : _GEN_3363; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3365 = 8'h25 == io_state_in_1 ? 8'h82 : _GEN_3364; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3366 = 8'h26 == io_state_in_1 ? 8'h95 : _GEN_3365; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3367 = 8'h27 == io_state_in_1 ? 8'h98 : _GEN_3366; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3368 = 8'h28 == io_state_in_1 ? 8'hd3 : _GEN_3367; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3369 = 8'h29 == io_state_in_1 ? 8'hde : _GEN_3368; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3370 = 8'h2a == io_state_in_1 ? 8'hc9 : _GEN_3369; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3371 = 8'h2b == io_state_in_1 ? 8'hc4 : _GEN_3370; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3372 = 8'h2c == io_state_in_1 ? 8'he7 : _GEN_3371; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3373 = 8'h2d == io_state_in_1 ? 8'hea : _GEN_3372; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3374 = 8'h2e == io_state_in_1 ? 8'hfd : _GEN_3373; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3375 = 8'h2f == io_state_in_1 ? 8'hf0 : _GEN_3374; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3376 = 8'h30 == io_state_in_1 ? 8'h6b : _GEN_3375; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3377 = 8'h31 == io_state_in_1 ? 8'h66 : _GEN_3376; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3378 = 8'h32 == io_state_in_1 ? 8'h71 : _GEN_3377; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3379 = 8'h33 == io_state_in_1 ? 8'h7c : _GEN_3378; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3380 = 8'h34 == io_state_in_1 ? 8'h5f : _GEN_3379; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3381 = 8'h35 == io_state_in_1 ? 8'h52 : _GEN_3380; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3382 = 8'h36 == io_state_in_1 ? 8'h45 : _GEN_3381; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3383 = 8'h37 == io_state_in_1 ? 8'h48 : _GEN_3382; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3384 = 8'h38 == io_state_in_1 ? 8'h3 : _GEN_3383; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3385 = 8'h39 == io_state_in_1 ? 8'he : _GEN_3384; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3386 = 8'h3a == io_state_in_1 ? 8'h19 : _GEN_3385; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3387 = 8'h3b == io_state_in_1 ? 8'h14 : _GEN_3386; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3388 = 8'h3c == io_state_in_1 ? 8'h37 : _GEN_3387; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3389 = 8'h3d == io_state_in_1 ? 8'h3a : _GEN_3388; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3390 = 8'h3e == io_state_in_1 ? 8'h2d : _GEN_3389; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3391 = 8'h3f == io_state_in_1 ? 8'h20 : _GEN_3390; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3392 = 8'h40 == io_state_in_1 ? 8'h6d : _GEN_3391; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3393 = 8'h41 == io_state_in_1 ? 8'h60 : _GEN_3392; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3394 = 8'h42 == io_state_in_1 ? 8'h77 : _GEN_3393; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3395 = 8'h43 == io_state_in_1 ? 8'h7a : _GEN_3394; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3396 = 8'h44 == io_state_in_1 ? 8'h59 : _GEN_3395; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3397 = 8'h45 == io_state_in_1 ? 8'h54 : _GEN_3396; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3398 = 8'h46 == io_state_in_1 ? 8'h43 : _GEN_3397; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3399 = 8'h47 == io_state_in_1 ? 8'h4e : _GEN_3398; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3400 = 8'h48 == io_state_in_1 ? 8'h5 : _GEN_3399; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3401 = 8'h49 == io_state_in_1 ? 8'h8 : _GEN_3400; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3402 = 8'h4a == io_state_in_1 ? 8'h1f : _GEN_3401; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3403 = 8'h4b == io_state_in_1 ? 8'h12 : _GEN_3402; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3404 = 8'h4c == io_state_in_1 ? 8'h31 : _GEN_3403; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3405 = 8'h4d == io_state_in_1 ? 8'h3c : _GEN_3404; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3406 = 8'h4e == io_state_in_1 ? 8'h2b : _GEN_3405; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3407 = 8'h4f == io_state_in_1 ? 8'h26 : _GEN_3406; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3408 = 8'h50 == io_state_in_1 ? 8'hbd : _GEN_3407; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3409 = 8'h51 == io_state_in_1 ? 8'hb0 : _GEN_3408; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3410 = 8'h52 == io_state_in_1 ? 8'ha7 : _GEN_3409; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3411 = 8'h53 == io_state_in_1 ? 8'haa : _GEN_3410; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3412 = 8'h54 == io_state_in_1 ? 8'h89 : _GEN_3411; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3413 = 8'h55 == io_state_in_1 ? 8'h84 : _GEN_3412; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3414 = 8'h56 == io_state_in_1 ? 8'h93 : _GEN_3413; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3415 = 8'h57 == io_state_in_1 ? 8'h9e : _GEN_3414; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3416 = 8'h58 == io_state_in_1 ? 8'hd5 : _GEN_3415; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3417 = 8'h59 == io_state_in_1 ? 8'hd8 : _GEN_3416; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3418 = 8'h5a == io_state_in_1 ? 8'hcf : _GEN_3417; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3419 = 8'h5b == io_state_in_1 ? 8'hc2 : _GEN_3418; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3420 = 8'h5c == io_state_in_1 ? 8'he1 : _GEN_3419; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3421 = 8'h5d == io_state_in_1 ? 8'hec : _GEN_3420; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3422 = 8'h5e == io_state_in_1 ? 8'hfb : _GEN_3421; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3423 = 8'h5f == io_state_in_1 ? 8'hf6 : _GEN_3422; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3424 = 8'h60 == io_state_in_1 ? 8'hd6 : _GEN_3423; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3425 = 8'h61 == io_state_in_1 ? 8'hdb : _GEN_3424; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3426 = 8'h62 == io_state_in_1 ? 8'hcc : _GEN_3425; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3427 = 8'h63 == io_state_in_1 ? 8'hc1 : _GEN_3426; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3428 = 8'h64 == io_state_in_1 ? 8'he2 : _GEN_3427; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3429 = 8'h65 == io_state_in_1 ? 8'hef : _GEN_3428; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3430 = 8'h66 == io_state_in_1 ? 8'hf8 : _GEN_3429; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3431 = 8'h67 == io_state_in_1 ? 8'hf5 : _GEN_3430; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3432 = 8'h68 == io_state_in_1 ? 8'hbe : _GEN_3431; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3433 = 8'h69 == io_state_in_1 ? 8'hb3 : _GEN_3432; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3434 = 8'h6a == io_state_in_1 ? 8'ha4 : _GEN_3433; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3435 = 8'h6b == io_state_in_1 ? 8'ha9 : _GEN_3434; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3436 = 8'h6c == io_state_in_1 ? 8'h8a : _GEN_3435; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3437 = 8'h6d == io_state_in_1 ? 8'h87 : _GEN_3436; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3438 = 8'h6e == io_state_in_1 ? 8'h90 : _GEN_3437; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3439 = 8'h6f == io_state_in_1 ? 8'h9d : _GEN_3438; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3440 = 8'h70 == io_state_in_1 ? 8'h6 : _GEN_3439; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3441 = 8'h71 == io_state_in_1 ? 8'hb : _GEN_3440; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3442 = 8'h72 == io_state_in_1 ? 8'h1c : _GEN_3441; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3443 = 8'h73 == io_state_in_1 ? 8'h11 : _GEN_3442; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3444 = 8'h74 == io_state_in_1 ? 8'h32 : _GEN_3443; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3445 = 8'h75 == io_state_in_1 ? 8'h3f : _GEN_3444; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3446 = 8'h76 == io_state_in_1 ? 8'h28 : _GEN_3445; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3447 = 8'h77 == io_state_in_1 ? 8'h25 : _GEN_3446; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3448 = 8'h78 == io_state_in_1 ? 8'h6e : _GEN_3447; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3449 = 8'h79 == io_state_in_1 ? 8'h63 : _GEN_3448; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3450 = 8'h7a == io_state_in_1 ? 8'h74 : _GEN_3449; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3451 = 8'h7b == io_state_in_1 ? 8'h79 : _GEN_3450; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3452 = 8'h7c == io_state_in_1 ? 8'h5a : _GEN_3451; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3453 = 8'h7d == io_state_in_1 ? 8'h57 : _GEN_3452; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3454 = 8'h7e == io_state_in_1 ? 8'h40 : _GEN_3453; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3455 = 8'h7f == io_state_in_1 ? 8'h4d : _GEN_3454; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3456 = 8'h80 == io_state_in_1 ? 8'hda : _GEN_3455; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3457 = 8'h81 == io_state_in_1 ? 8'hd7 : _GEN_3456; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3458 = 8'h82 == io_state_in_1 ? 8'hc0 : _GEN_3457; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3459 = 8'h83 == io_state_in_1 ? 8'hcd : _GEN_3458; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3460 = 8'h84 == io_state_in_1 ? 8'hee : _GEN_3459; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3461 = 8'h85 == io_state_in_1 ? 8'he3 : _GEN_3460; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3462 = 8'h86 == io_state_in_1 ? 8'hf4 : _GEN_3461; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3463 = 8'h87 == io_state_in_1 ? 8'hf9 : _GEN_3462; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3464 = 8'h88 == io_state_in_1 ? 8'hb2 : _GEN_3463; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3465 = 8'h89 == io_state_in_1 ? 8'hbf : _GEN_3464; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3466 = 8'h8a == io_state_in_1 ? 8'ha8 : _GEN_3465; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3467 = 8'h8b == io_state_in_1 ? 8'ha5 : _GEN_3466; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3468 = 8'h8c == io_state_in_1 ? 8'h86 : _GEN_3467; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3469 = 8'h8d == io_state_in_1 ? 8'h8b : _GEN_3468; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3470 = 8'h8e == io_state_in_1 ? 8'h9c : _GEN_3469; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3471 = 8'h8f == io_state_in_1 ? 8'h91 : _GEN_3470; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3472 = 8'h90 == io_state_in_1 ? 8'ha : _GEN_3471; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3473 = 8'h91 == io_state_in_1 ? 8'h7 : _GEN_3472; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3474 = 8'h92 == io_state_in_1 ? 8'h10 : _GEN_3473; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3475 = 8'h93 == io_state_in_1 ? 8'h1d : _GEN_3474; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3476 = 8'h94 == io_state_in_1 ? 8'h3e : _GEN_3475; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3477 = 8'h95 == io_state_in_1 ? 8'h33 : _GEN_3476; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3478 = 8'h96 == io_state_in_1 ? 8'h24 : _GEN_3477; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3479 = 8'h97 == io_state_in_1 ? 8'h29 : _GEN_3478; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3480 = 8'h98 == io_state_in_1 ? 8'h62 : _GEN_3479; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3481 = 8'h99 == io_state_in_1 ? 8'h6f : _GEN_3480; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3482 = 8'h9a == io_state_in_1 ? 8'h78 : _GEN_3481; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3483 = 8'h9b == io_state_in_1 ? 8'h75 : _GEN_3482; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3484 = 8'h9c == io_state_in_1 ? 8'h56 : _GEN_3483; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3485 = 8'h9d == io_state_in_1 ? 8'h5b : _GEN_3484; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3486 = 8'h9e == io_state_in_1 ? 8'h4c : _GEN_3485; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3487 = 8'h9f == io_state_in_1 ? 8'h41 : _GEN_3486; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3488 = 8'ha0 == io_state_in_1 ? 8'h61 : _GEN_3487; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3489 = 8'ha1 == io_state_in_1 ? 8'h6c : _GEN_3488; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3490 = 8'ha2 == io_state_in_1 ? 8'h7b : _GEN_3489; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3491 = 8'ha3 == io_state_in_1 ? 8'h76 : _GEN_3490; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3492 = 8'ha4 == io_state_in_1 ? 8'h55 : _GEN_3491; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3493 = 8'ha5 == io_state_in_1 ? 8'h58 : _GEN_3492; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3494 = 8'ha6 == io_state_in_1 ? 8'h4f : _GEN_3493; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3495 = 8'ha7 == io_state_in_1 ? 8'h42 : _GEN_3494; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3496 = 8'ha8 == io_state_in_1 ? 8'h9 : _GEN_3495; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3497 = 8'ha9 == io_state_in_1 ? 8'h4 : _GEN_3496; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3498 = 8'haa == io_state_in_1 ? 8'h13 : _GEN_3497; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3499 = 8'hab == io_state_in_1 ? 8'h1e : _GEN_3498; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3500 = 8'hac == io_state_in_1 ? 8'h3d : _GEN_3499; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3501 = 8'had == io_state_in_1 ? 8'h30 : _GEN_3500; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3502 = 8'hae == io_state_in_1 ? 8'h27 : _GEN_3501; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3503 = 8'haf == io_state_in_1 ? 8'h2a : _GEN_3502; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3504 = 8'hb0 == io_state_in_1 ? 8'hb1 : _GEN_3503; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3505 = 8'hb1 == io_state_in_1 ? 8'hbc : _GEN_3504; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3506 = 8'hb2 == io_state_in_1 ? 8'hab : _GEN_3505; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3507 = 8'hb3 == io_state_in_1 ? 8'ha6 : _GEN_3506; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3508 = 8'hb4 == io_state_in_1 ? 8'h85 : _GEN_3507; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3509 = 8'hb5 == io_state_in_1 ? 8'h88 : _GEN_3508; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3510 = 8'hb6 == io_state_in_1 ? 8'h9f : _GEN_3509; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3511 = 8'hb7 == io_state_in_1 ? 8'h92 : _GEN_3510; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3512 = 8'hb8 == io_state_in_1 ? 8'hd9 : _GEN_3511; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3513 = 8'hb9 == io_state_in_1 ? 8'hd4 : _GEN_3512; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3514 = 8'hba == io_state_in_1 ? 8'hc3 : _GEN_3513; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3515 = 8'hbb == io_state_in_1 ? 8'hce : _GEN_3514; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3516 = 8'hbc == io_state_in_1 ? 8'hed : _GEN_3515; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3517 = 8'hbd == io_state_in_1 ? 8'he0 : _GEN_3516; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3518 = 8'hbe == io_state_in_1 ? 8'hf7 : _GEN_3517; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3519 = 8'hbf == io_state_in_1 ? 8'hfa : _GEN_3518; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3520 = 8'hc0 == io_state_in_1 ? 8'hb7 : _GEN_3519; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3521 = 8'hc1 == io_state_in_1 ? 8'hba : _GEN_3520; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3522 = 8'hc2 == io_state_in_1 ? 8'had : _GEN_3521; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3523 = 8'hc3 == io_state_in_1 ? 8'ha0 : _GEN_3522; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3524 = 8'hc4 == io_state_in_1 ? 8'h83 : _GEN_3523; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3525 = 8'hc5 == io_state_in_1 ? 8'h8e : _GEN_3524; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3526 = 8'hc6 == io_state_in_1 ? 8'h99 : _GEN_3525; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3527 = 8'hc7 == io_state_in_1 ? 8'h94 : _GEN_3526; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3528 = 8'hc8 == io_state_in_1 ? 8'hdf : _GEN_3527; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3529 = 8'hc9 == io_state_in_1 ? 8'hd2 : _GEN_3528; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3530 = 8'hca == io_state_in_1 ? 8'hc5 : _GEN_3529; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3531 = 8'hcb == io_state_in_1 ? 8'hc8 : _GEN_3530; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3532 = 8'hcc == io_state_in_1 ? 8'heb : _GEN_3531; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3533 = 8'hcd == io_state_in_1 ? 8'he6 : _GEN_3532; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3534 = 8'hce == io_state_in_1 ? 8'hf1 : _GEN_3533; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3535 = 8'hcf == io_state_in_1 ? 8'hfc : _GEN_3534; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3536 = 8'hd0 == io_state_in_1 ? 8'h67 : _GEN_3535; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3537 = 8'hd1 == io_state_in_1 ? 8'h6a : _GEN_3536; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3538 = 8'hd2 == io_state_in_1 ? 8'h7d : _GEN_3537; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3539 = 8'hd3 == io_state_in_1 ? 8'h70 : _GEN_3538; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3540 = 8'hd4 == io_state_in_1 ? 8'h53 : _GEN_3539; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3541 = 8'hd5 == io_state_in_1 ? 8'h5e : _GEN_3540; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3542 = 8'hd6 == io_state_in_1 ? 8'h49 : _GEN_3541; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3543 = 8'hd7 == io_state_in_1 ? 8'h44 : _GEN_3542; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3544 = 8'hd8 == io_state_in_1 ? 8'hf : _GEN_3543; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3545 = 8'hd9 == io_state_in_1 ? 8'h2 : _GEN_3544; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3546 = 8'hda == io_state_in_1 ? 8'h15 : _GEN_3545; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3547 = 8'hdb == io_state_in_1 ? 8'h18 : _GEN_3546; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3548 = 8'hdc == io_state_in_1 ? 8'h3b : _GEN_3547; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3549 = 8'hdd == io_state_in_1 ? 8'h36 : _GEN_3548; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3550 = 8'hde == io_state_in_1 ? 8'h21 : _GEN_3549; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3551 = 8'hdf == io_state_in_1 ? 8'h2c : _GEN_3550; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3552 = 8'he0 == io_state_in_1 ? 8'hc : _GEN_3551; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3553 = 8'he1 == io_state_in_1 ? 8'h1 : _GEN_3552; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3554 = 8'he2 == io_state_in_1 ? 8'h16 : _GEN_3553; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3555 = 8'he3 == io_state_in_1 ? 8'h1b : _GEN_3554; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3556 = 8'he4 == io_state_in_1 ? 8'h38 : _GEN_3555; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3557 = 8'he5 == io_state_in_1 ? 8'h35 : _GEN_3556; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3558 = 8'he6 == io_state_in_1 ? 8'h22 : _GEN_3557; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3559 = 8'he7 == io_state_in_1 ? 8'h2f : _GEN_3558; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3560 = 8'he8 == io_state_in_1 ? 8'h64 : _GEN_3559; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3561 = 8'he9 == io_state_in_1 ? 8'h69 : _GEN_3560; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3562 = 8'hea == io_state_in_1 ? 8'h7e : _GEN_3561; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3563 = 8'heb == io_state_in_1 ? 8'h73 : _GEN_3562; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3564 = 8'hec == io_state_in_1 ? 8'h50 : _GEN_3563; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3565 = 8'hed == io_state_in_1 ? 8'h5d : _GEN_3564; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3566 = 8'hee == io_state_in_1 ? 8'h4a : _GEN_3565; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3567 = 8'hef == io_state_in_1 ? 8'h47 : _GEN_3566; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3568 = 8'hf0 == io_state_in_1 ? 8'hdc : _GEN_3567; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3569 = 8'hf1 == io_state_in_1 ? 8'hd1 : _GEN_3568; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3570 = 8'hf2 == io_state_in_1 ? 8'hc6 : _GEN_3569; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3571 = 8'hf3 == io_state_in_1 ? 8'hcb : _GEN_3570; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3572 = 8'hf4 == io_state_in_1 ? 8'he8 : _GEN_3571; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3573 = 8'hf5 == io_state_in_1 ? 8'he5 : _GEN_3572; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3574 = 8'hf6 == io_state_in_1 ? 8'hf2 : _GEN_3573; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3575 = 8'hf7 == io_state_in_1 ? 8'hff : _GEN_3574; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3576 = 8'hf8 == io_state_in_1 ? 8'hb4 : _GEN_3575; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3577 = 8'hf9 == io_state_in_1 ? 8'hb9 : _GEN_3576; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3578 = 8'hfa == io_state_in_1 ? 8'hae : _GEN_3577; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3579 = 8'hfb == io_state_in_1 ? 8'ha3 : _GEN_3578; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3580 = 8'hfc == io_state_in_1 ? 8'h80 : _GEN_3579; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3581 = 8'hfd == io_state_in_1 ? 8'h8d : _GEN_3580; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3582 = 8'hfe == io_state_in_1 ? 8'h9a : _GEN_3581; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _GEN_3583 = 8'hff == io_state_in_1 ? 8'h97 : _GEN_3582; // @[InvMixColumns.scala 129:{41,41}]
  wire [7:0] _tmp_state_3_T = _GEN_3327 ^ _GEN_3583; // @[InvMixColumns.scala 129:41]
  wire [7:0] _GEN_3585 = 8'h1 == io_state_in_2 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3586 = 8'h2 == io_state_in_2 ? 8'h12 : _GEN_3585; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3587 = 8'h3 == io_state_in_2 ? 8'h1b : _GEN_3586; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3588 = 8'h4 == io_state_in_2 ? 8'h24 : _GEN_3587; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3589 = 8'h5 == io_state_in_2 ? 8'h2d : _GEN_3588; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3590 = 8'h6 == io_state_in_2 ? 8'h36 : _GEN_3589; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3591 = 8'h7 == io_state_in_2 ? 8'h3f : _GEN_3590; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3592 = 8'h8 == io_state_in_2 ? 8'h48 : _GEN_3591; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3593 = 8'h9 == io_state_in_2 ? 8'h41 : _GEN_3592; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3594 = 8'ha == io_state_in_2 ? 8'h5a : _GEN_3593; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3595 = 8'hb == io_state_in_2 ? 8'h53 : _GEN_3594; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3596 = 8'hc == io_state_in_2 ? 8'h6c : _GEN_3595; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3597 = 8'hd == io_state_in_2 ? 8'h65 : _GEN_3596; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3598 = 8'he == io_state_in_2 ? 8'h7e : _GEN_3597; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3599 = 8'hf == io_state_in_2 ? 8'h77 : _GEN_3598; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3600 = 8'h10 == io_state_in_2 ? 8'h90 : _GEN_3599; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3601 = 8'h11 == io_state_in_2 ? 8'h99 : _GEN_3600; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3602 = 8'h12 == io_state_in_2 ? 8'h82 : _GEN_3601; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3603 = 8'h13 == io_state_in_2 ? 8'h8b : _GEN_3602; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3604 = 8'h14 == io_state_in_2 ? 8'hb4 : _GEN_3603; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3605 = 8'h15 == io_state_in_2 ? 8'hbd : _GEN_3604; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3606 = 8'h16 == io_state_in_2 ? 8'ha6 : _GEN_3605; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3607 = 8'h17 == io_state_in_2 ? 8'haf : _GEN_3606; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3608 = 8'h18 == io_state_in_2 ? 8'hd8 : _GEN_3607; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3609 = 8'h19 == io_state_in_2 ? 8'hd1 : _GEN_3608; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3610 = 8'h1a == io_state_in_2 ? 8'hca : _GEN_3609; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3611 = 8'h1b == io_state_in_2 ? 8'hc3 : _GEN_3610; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3612 = 8'h1c == io_state_in_2 ? 8'hfc : _GEN_3611; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3613 = 8'h1d == io_state_in_2 ? 8'hf5 : _GEN_3612; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3614 = 8'h1e == io_state_in_2 ? 8'hee : _GEN_3613; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3615 = 8'h1f == io_state_in_2 ? 8'he7 : _GEN_3614; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3616 = 8'h20 == io_state_in_2 ? 8'h3b : _GEN_3615; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3617 = 8'h21 == io_state_in_2 ? 8'h32 : _GEN_3616; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3618 = 8'h22 == io_state_in_2 ? 8'h29 : _GEN_3617; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3619 = 8'h23 == io_state_in_2 ? 8'h20 : _GEN_3618; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3620 = 8'h24 == io_state_in_2 ? 8'h1f : _GEN_3619; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3621 = 8'h25 == io_state_in_2 ? 8'h16 : _GEN_3620; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3622 = 8'h26 == io_state_in_2 ? 8'hd : _GEN_3621; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3623 = 8'h27 == io_state_in_2 ? 8'h4 : _GEN_3622; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3624 = 8'h28 == io_state_in_2 ? 8'h73 : _GEN_3623; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3625 = 8'h29 == io_state_in_2 ? 8'h7a : _GEN_3624; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3626 = 8'h2a == io_state_in_2 ? 8'h61 : _GEN_3625; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3627 = 8'h2b == io_state_in_2 ? 8'h68 : _GEN_3626; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3628 = 8'h2c == io_state_in_2 ? 8'h57 : _GEN_3627; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3629 = 8'h2d == io_state_in_2 ? 8'h5e : _GEN_3628; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3630 = 8'h2e == io_state_in_2 ? 8'h45 : _GEN_3629; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3631 = 8'h2f == io_state_in_2 ? 8'h4c : _GEN_3630; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3632 = 8'h30 == io_state_in_2 ? 8'hab : _GEN_3631; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3633 = 8'h31 == io_state_in_2 ? 8'ha2 : _GEN_3632; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3634 = 8'h32 == io_state_in_2 ? 8'hb9 : _GEN_3633; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3635 = 8'h33 == io_state_in_2 ? 8'hb0 : _GEN_3634; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3636 = 8'h34 == io_state_in_2 ? 8'h8f : _GEN_3635; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3637 = 8'h35 == io_state_in_2 ? 8'h86 : _GEN_3636; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3638 = 8'h36 == io_state_in_2 ? 8'h9d : _GEN_3637; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3639 = 8'h37 == io_state_in_2 ? 8'h94 : _GEN_3638; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3640 = 8'h38 == io_state_in_2 ? 8'he3 : _GEN_3639; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3641 = 8'h39 == io_state_in_2 ? 8'hea : _GEN_3640; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3642 = 8'h3a == io_state_in_2 ? 8'hf1 : _GEN_3641; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3643 = 8'h3b == io_state_in_2 ? 8'hf8 : _GEN_3642; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3644 = 8'h3c == io_state_in_2 ? 8'hc7 : _GEN_3643; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3645 = 8'h3d == io_state_in_2 ? 8'hce : _GEN_3644; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3646 = 8'h3e == io_state_in_2 ? 8'hd5 : _GEN_3645; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3647 = 8'h3f == io_state_in_2 ? 8'hdc : _GEN_3646; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3648 = 8'h40 == io_state_in_2 ? 8'h76 : _GEN_3647; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3649 = 8'h41 == io_state_in_2 ? 8'h7f : _GEN_3648; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3650 = 8'h42 == io_state_in_2 ? 8'h64 : _GEN_3649; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3651 = 8'h43 == io_state_in_2 ? 8'h6d : _GEN_3650; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3652 = 8'h44 == io_state_in_2 ? 8'h52 : _GEN_3651; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3653 = 8'h45 == io_state_in_2 ? 8'h5b : _GEN_3652; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3654 = 8'h46 == io_state_in_2 ? 8'h40 : _GEN_3653; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3655 = 8'h47 == io_state_in_2 ? 8'h49 : _GEN_3654; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3656 = 8'h48 == io_state_in_2 ? 8'h3e : _GEN_3655; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3657 = 8'h49 == io_state_in_2 ? 8'h37 : _GEN_3656; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3658 = 8'h4a == io_state_in_2 ? 8'h2c : _GEN_3657; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3659 = 8'h4b == io_state_in_2 ? 8'h25 : _GEN_3658; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3660 = 8'h4c == io_state_in_2 ? 8'h1a : _GEN_3659; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3661 = 8'h4d == io_state_in_2 ? 8'h13 : _GEN_3660; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3662 = 8'h4e == io_state_in_2 ? 8'h8 : _GEN_3661; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3663 = 8'h4f == io_state_in_2 ? 8'h1 : _GEN_3662; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3664 = 8'h50 == io_state_in_2 ? 8'he6 : _GEN_3663; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3665 = 8'h51 == io_state_in_2 ? 8'hef : _GEN_3664; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3666 = 8'h52 == io_state_in_2 ? 8'hf4 : _GEN_3665; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3667 = 8'h53 == io_state_in_2 ? 8'hfd : _GEN_3666; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3668 = 8'h54 == io_state_in_2 ? 8'hc2 : _GEN_3667; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3669 = 8'h55 == io_state_in_2 ? 8'hcb : _GEN_3668; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3670 = 8'h56 == io_state_in_2 ? 8'hd0 : _GEN_3669; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3671 = 8'h57 == io_state_in_2 ? 8'hd9 : _GEN_3670; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3672 = 8'h58 == io_state_in_2 ? 8'hae : _GEN_3671; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3673 = 8'h59 == io_state_in_2 ? 8'ha7 : _GEN_3672; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3674 = 8'h5a == io_state_in_2 ? 8'hbc : _GEN_3673; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3675 = 8'h5b == io_state_in_2 ? 8'hb5 : _GEN_3674; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3676 = 8'h5c == io_state_in_2 ? 8'h8a : _GEN_3675; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3677 = 8'h5d == io_state_in_2 ? 8'h83 : _GEN_3676; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3678 = 8'h5e == io_state_in_2 ? 8'h98 : _GEN_3677; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3679 = 8'h5f == io_state_in_2 ? 8'h91 : _GEN_3678; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3680 = 8'h60 == io_state_in_2 ? 8'h4d : _GEN_3679; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3681 = 8'h61 == io_state_in_2 ? 8'h44 : _GEN_3680; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3682 = 8'h62 == io_state_in_2 ? 8'h5f : _GEN_3681; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3683 = 8'h63 == io_state_in_2 ? 8'h56 : _GEN_3682; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3684 = 8'h64 == io_state_in_2 ? 8'h69 : _GEN_3683; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3685 = 8'h65 == io_state_in_2 ? 8'h60 : _GEN_3684; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3686 = 8'h66 == io_state_in_2 ? 8'h7b : _GEN_3685; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3687 = 8'h67 == io_state_in_2 ? 8'h72 : _GEN_3686; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3688 = 8'h68 == io_state_in_2 ? 8'h5 : _GEN_3687; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3689 = 8'h69 == io_state_in_2 ? 8'hc : _GEN_3688; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3690 = 8'h6a == io_state_in_2 ? 8'h17 : _GEN_3689; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3691 = 8'h6b == io_state_in_2 ? 8'h1e : _GEN_3690; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3692 = 8'h6c == io_state_in_2 ? 8'h21 : _GEN_3691; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3693 = 8'h6d == io_state_in_2 ? 8'h28 : _GEN_3692; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3694 = 8'h6e == io_state_in_2 ? 8'h33 : _GEN_3693; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3695 = 8'h6f == io_state_in_2 ? 8'h3a : _GEN_3694; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3696 = 8'h70 == io_state_in_2 ? 8'hdd : _GEN_3695; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3697 = 8'h71 == io_state_in_2 ? 8'hd4 : _GEN_3696; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3698 = 8'h72 == io_state_in_2 ? 8'hcf : _GEN_3697; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3699 = 8'h73 == io_state_in_2 ? 8'hc6 : _GEN_3698; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3700 = 8'h74 == io_state_in_2 ? 8'hf9 : _GEN_3699; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3701 = 8'h75 == io_state_in_2 ? 8'hf0 : _GEN_3700; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3702 = 8'h76 == io_state_in_2 ? 8'heb : _GEN_3701; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3703 = 8'h77 == io_state_in_2 ? 8'he2 : _GEN_3702; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3704 = 8'h78 == io_state_in_2 ? 8'h95 : _GEN_3703; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3705 = 8'h79 == io_state_in_2 ? 8'h9c : _GEN_3704; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3706 = 8'h7a == io_state_in_2 ? 8'h87 : _GEN_3705; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3707 = 8'h7b == io_state_in_2 ? 8'h8e : _GEN_3706; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3708 = 8'h7c == io_state_in_2 ? 8'hb1 : _GEN_3707; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3709 = 8'h7d == io_state_in_2 ? 8'hb8 : _GEN_3708; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3710 = 8'h7e == io_state_in_2 ? 8'ha3 : _GEN_3709; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3711 = 8'h7f == io_state_in_2 ? 8'haa : _GEN_3710; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3712 = 8'h80 == io_state_in_2 ? 8'hec : _GEN_3711; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3713 = 8'h81 == io_state_in_2 ? 8'he5 : _GEN_3712; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3714 = 8'h82 == io_state_in_2 ? 8'hfe : _GEN_3713; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3715 = 8'h83 == io_state_in_2 ? 8'hf7 : _GEN_3714; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3716 = 8'h84 == io_state_in_2 ? 8'hc8 : _GEN_3715; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3717 = 8'h85 == io_state_in_2 ? 8'hc1 : _GEN_3716; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3718 = 8'h86 == io_state_in_2 ? 8'hda : _GEN_3717; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3719 = 8'h87 == io_state_in_2 ? 8'hd3 : _GEN_3718; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3720 = 8'h88 == io_state_in_2 ? 8'ha4 : _GEN_3719; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3721 = 8'h89 == io_state_in_2 ? 8'had : _GEN_3720; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3722 = 8'h8a == io_state_in_2 ? 8'hb6 : _GEN_3721; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3723 = 8'h8b == io_state_in_2 ? 8'hbf : _GEN_3722; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3724 = 8'h8c == io_state_in_2 ? 8'h80 : _GEN_3723; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3725 = 8'h8d == io_state_in_2 ? 8'h89 : _GEN_3724; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3726 = 8'h8e == io_state_in_2 ? 8'h92 : _GEN_3725; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3727 = 8'h8f == io_state_in_2 ? 8'h9b : _GEN_3726; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3728 = 8'h90 == io_state_in_2 ? 8'h7c : _GEN_3727; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3729 = 8'h91 == io_state_in_2 ? 8'h75 : _GEN_3728; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3730 = 8'h92 == io_state_in_2 ? 8'h6e : _GEN_3729; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3731 = 8'h93 == io_state_in_2 ? 8'h67 : _GEN_3730; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3732 = 8'h94 == io_state_in_2 ? 8'h58 : _GEN_3731; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3733 = 8'h95 == io_state_in_2 ? 8'h51 : _GEN_3732; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3734 = 8'h96 == io_state_in_2 ? 8'h4a : _GEN_3733; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3735 = 8'h97 == io_state_in_2 ? 8'h43 : _GEN_3734; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3736 = 8'h98 == io_state_in_2 ? 8'h34 : _GEN_3735; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3737 = 8'h99 == io_state_in_2 ? 8'h3d : _GEN_3736; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3738 = 8'h9a == io_state_in_2 ? 8'h26 : _GEN_3737; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3739 = 8'h9b == io_state_in_2 ? 8'h2f : _GEN_3738; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3740 = 8'h9c == io_state_in_2 ? 8'h10 : _GEN_3739; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3741 = 8'h9d == io_state_in_2 ? 8'h19 : _GEN_3740; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3742 = 8'h9e == io_state_in_2 ? 8'h2 : _GEN_3741; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3743 = 8'h9f == io_state_in_2 ? 8'hb : _GEN_3742; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3744 = 8'ha0 == io_state_in_2 ? 8'hd7 : _GEN_3743; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3745 = 8'ha1 == io_state_in_2 ? 8'hde : _GEN_3744; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3746 = 8'ha2 == io_state_in_2 ? 8'hc5 : _GEN_3745; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3747 = 8'ha3 == io_state_in_2 ? 8'hcc : _GEN_3746; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3748 = 8'ha4 == io_state_in_2 ? 8'hf3 : _GEN_3747; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3749 = 8'ha5 == io_state_in_2 ? 8'hfa : _GEN_3748; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3750 = 8'ha6 == io_state_in_2 ? 8'he1 : _GEN_3749; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3751 = 8'ha7 == io_state_in_2 ? 8'he8 : _GEN_3750; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3752 = 8'ha8 == io_state_in_2 ? 8'h9f : _GEN_3751; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3753 = 8'ha9 == io_state_in_2 ? 8'h96 : _GEN_3752; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3754 = 8'haa == io_state_in_2 ? 8'h8d : _GEN_3753; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3755 = 8'hab == io_state_in_2 ? 8'h84 : _GEN_3754; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3756 = 8'hac == io_state_in_2 ? 8'hbb : _GEN_3755; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3757 = 8'had == io_state_in_2 ? 8'hb2 : _GEN_3756; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3758 = 8'hae == io_state_in_2 ? 8'ha9 : _GEN_3757; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3759 = 8'haf == io_state_in_2 ? 8'ha0 : _GEN_3758; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3760 = 8'hb0 == io_state_in_2 ? 8'h47 : _GEN_3759; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3761 = 8'hb1 == io_state_in_2 ? 8'h4e : _GEN_3760; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3762 = 8'hb2 == io_state_in_2 ? 8'h55 : _GEN_3761; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3763 = 8'hb3 == io_state_in_2 ? 8'h5c : _GEN_3762; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3764 = 8'hb4 == io_state_in_2 ? 8'h63 : _GEN_3763; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3765 = 8'hb5 == io_state_in_2 ? 8'h6a : _GEN_3764; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3766 = 8'hb6 == io_state_in_2 ? 8'h71 : _GEN_3765; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3767 = 8'hb7 == io_state_in_2 ? 8'h78 : _GEN_3766; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3768 = 8'hb8 == io_state_in_2 ? 8'hf : _GEN_3767; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3769 = 8'hb9 == io_state_in_2 ? 8'h6 : _GEN_3768; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3770 = 8'hba == io_state_in_2 ? 8'h1d : _GEN_3769; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3771 = 8'hbb == io_state_in_2 ? 8'h14 : _GEN_3770; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3772 = 8'hbc == io_state_in_2 ? 8'h2b : _GEN_3771; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3773 = 8'hbd == io_state_in_2 ? 8'h22 : _GEN_3772; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3774 = 8'hbe == io_state_in_2 ? 8'h39 : _GEN_3773; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3775 = 8'hbf == io_state_in_2 ? 8'h30 : _GEN_3774; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3776 = 8'hc0 == io_state_in_2 ? 8'h9a : _GEN_3775; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3777 = 8'hc1 == io_state_in_2 ? 8'h93 : _GEN_3776; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3778 = 8'hc2 == io_state_in_2 ? 8'h88 : _GEN_3777; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3779 = 8'hc3 == io_state_in_2 ? 8'h81 : _GEN_3778; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3780 = 8'hc4 == io_state_in_2 ? 8'hbe : _GEN_3779; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3781 = 8'hc5 == io_state_in_2 ? 8'hb7 : _GEN_3780; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3782 = 8'hc6 == io_state_in_2 ? 8'hac : _GEN_3781; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3783 = 8'hc7 == io_state_in_2 ? 8'ha5 : _GEN_3782; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3784 = 8'hc8 == io_state_in_2 ? 8'hd2 : _GEN_3783; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3785 = 8'hc9 == io_state_in_2 ? 8'hdb : _GEN_3784; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3786 = 8'hca == io_state_in_2 ? 8'hc0 : _GEN_3785; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3787 = 8'hcb == io_state_in_2 ? 8'hc9 : _GEN_3786; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3788 = 8'hcc == io_state_in_2 ? 8'hf6 : _GEN_3787; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3789 = 8'hcd == io_state_in_2 ? 8'hff : _GEN_3788; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3790 = 8'hce == io_state_in_2 ? 8'he4 : _GEN_3789; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3791 = 8'hcf == io_state_in_2 ? 8'hed : _GEN_3790; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3792 = 8'hd0 == io_state_in_2 ? 8'ha : _GEN_3791; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3793 = 8'hd1 == io_state_in_2 ? 8'h3 : _GEN_3792; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3794 = 8'hd2 == io_state_in_2 ? 8'h18 : _GEN_3793; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3795 = 8'hd3 == io_state_in_2 ? 8'h11 : _GEN_3794; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3796 = 8'hd4 == io_state_in_2 ? 8'h2e : _GEN_3795; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3797 = 8'hd5 == io_state_in_2 ? 8'h27 : _GEN_3796; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3798 = 8'hd6 == io_state_in_2 ? 8'h3c : _GEN_3797; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3799 = 8'hd7 == io_state_in_2 ? 8'h35 : _GEN_3798; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3800 = 8'hd8 == io_state_in_2 ? 8'h42 : _GEN_3799; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3801 = 8'hd9 == io_state_in_2 ? 8'h4b : _GEN_3800; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3802 = 8'hda == io_state_in_2 ? 8'h50 : _GEN_3801; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3803 = 8'hdb == io_state_in_2 ? 8'h59 : _GEN_3802; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3804 = 8'hdc == io_state_in_2 ? 8'h66 : _GEN_3803; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3805 = 8'hdd == io_state_in_2 ? 8'h6f : _GEN_3804; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3806 = 8'hde == io_state_in_2 ? 8'h74 : _GEN_3805; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3807 = 8'hdf == io_state_in_2 ? 8'h7d : _GEN_3806; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3808 = 8'he0 == io_state_in_2 ? 8'ha1 : _GEN_3807; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3809 = 8'he1 == io_state_in_2 ? 8'ha8 : _GEN_3808; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3810 = 8'he2 == io_state_in_2 ? 8'hb3 : _GEN_3809; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3811 = 8'he3 == io_state_in_2 ? 8'hba : _GEN_3810; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3812 = 8'he4 == io_state_in_2 ? 8'h85 : _GEN_3811; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3813 = 8'he5 == io_state_in_2 ? 8'h8c : _GEN_3812; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3814 = 8'he6 == io_state_in_2 ? 8'h97 : _GEN_3813; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3815 = 8'he7 == io_state_in_2 ? 8'h9e : _GEN_3814; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3816 = 8'he8 == io_state_in_2 ? 8'he9 : _GEN_3815; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3817 = 8'he9 == io_state_in_2 ? 8'he0 : _GEN_3816; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3818 = 8'hea == io_state_in_2 ? 8'hfb : _GEN_3817; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3819 = 8'heb == io_state_in_2 ? 8'hf2 : _GEN_3818; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3820 = 8'hec == io_state_in_2 ? 8'hcd : _GEN_3819; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3821 = 8'hed == io_state_in_2 ? 8'hc4 : _GEN_3820; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3822 = 8'hee == io_state_in_2 ? 8'hdf : _GEN_3821; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3823 = 8'hef == io_state_in_2 ? 8'hd6 : _GEN_3822; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3824 = 8'hf0 == io_state_in_2 ? 8'h31 : _GEN_3823; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3825 = 8'hf1 == io_state_in_2 ? 8'h38 : _GEN_3824; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3826 = 8'hf2 == io_state_in_2 ? 8'h23 : _GEN_3825; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3827 = 8'hf3 == io_state_in_2 ? 8'h2a : _GEN_3826; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3828 = 8'hf4 == io_state_in_2 ? 8'h15 : _GEN_3827; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3829 = 8'hf5 == io_state_in_2 ? 8'h1c : _GEN_3828; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3830 = 8'hf6 == io_state_in_2 ? 8'h7 : _GEN_3829; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3831 = 8'hf7 == io_state_in_2 ? 8'he : _GEN_3830; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3832 = 8'hf8 == io_state_in_2 ? 8'h79 : _GEN_3831; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3833 = 8'hf9 == io_state_in_2 ? 8'h70 : _GEN_3832; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3834 = 8'hfa == io_state_in_2 ? 8'h6b : _GEN_3833; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3835 = 8'hfb == io_state_in_2 ? 8'h62 : _GEN_3834; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3836 = 8'hfc == io_state_in_2 ? 8'h5d : _GEN_3835; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3837 = 8'hfd == io_state_in_2 ? 8'h54 : _GEN_3836; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3838 = 8'hfe == io_state_in_2 ? 8'h4f : _GEN_3837; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _GEN_3839 = 8'hff == io_state_in_2 ? 8'h46 : _GEN_3838; // @[InvMixColumns.scala 129:{65,65}]
  wire [7:0] _tmp_state_3_T_1 = _tmp_state_3_T ^ _GEN_3839; // @[InvMixColumns.scala 129:65]
  wire [7:0] _GEN_3841 = 8'h1 == io_state_in_3 ? 8'he : 8'h0; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3842 = 8'h2 == io_state_in_3 ? 8'h1c : _GEN_3841; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3843 = 8'h3 == io_state_in_3 ? 8'h12 : _GEN_3842; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3844 = 8'h4 == io_state_in_3 ? 8'h38 : _GEN_3843; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3845 = 8'h5 == io_state_in_3 ? 8'h36 : _GEN_3844; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3846 = 8'h6 == io_state_in_3 ? 8'h24 : _GEN_3845; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3847 = 8'h7 == io_state_in_3 ? 8'h2a : _GEN_3846; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3848 = 8'h8 == io_state_in_3 ? 8'h70 : _GEN_3847; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3849 = 8'h9 == io_state_in_3 ? 8'h7e : _GEN_3848; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3850 = 8'ha == io_state_in_3 ? 8'h6c : _GEN_3849; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3851 = 8'hb == io_state_in_3 ? 8'h62 : _GEN_3850; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3852 = 8'hc == io_state_in_3 ? 8'h48 : _GEN_3851; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3853 = 8'hd == io_state_in_3 ? 8'h46 : _GEN_3852; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3854 = 8'he == io_state_in_3 ? 8'h54 : _GEN_3853; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3855 = 8'hf == io_state_in_3 ? 8'h5a : _GEN_3854; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3856 = 8'h10 == io_state_in_3 ? 8'he0 : _GEN_3855; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3857 = 8'h11 == io_state_in_3 ? 8'hee : _GEN_3856; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3858 = 8'h12 == io_state_in_3 ? 8'hfc : _GEN_3857; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3859 = 8'h13 == io_state_in_3 ? 8'hf2 : _GEN_3858; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3860 = 8'h14 == io_state_in_3 ? 8'hd8 : _GEN_3859; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3861 = 8'h15 == io_state_in_3 ? 8'hd6 : _GEN_3860; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3862 = 8'h16 == io_state_in_3 ? 8'hc4 : _GEN_3861; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3863 = 8'h17 == io_state_in_3 ? 8'hca : _GEN_3862; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3864 = 8'h18 == io_state_in_3 ? 8'h90 : _GEN_3863; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3865 = 8'h19 == io_state_in_3 ? 8'h9e : _GEN_3864; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3866 = 8'h1a == io_state_in_3 ? 8'h8c : _GEN_3865; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3867 = 8'h1b == io_state_in_3 ? 8'h82 : _GEN_3866; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3868 = 8'h1c == io_state_in_3 ? 8'ha8 : _GEN_3867; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3869 = 8'h1d == io_state_in_3 ? 8'ha6 : _GEN_3868; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3870 = 8'h1e == io_state_in_3 ? 8'hb4 : _GEN_3869; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3871 = 8'h1f == io_state_in_3 ? 8'hba : _GEN_3870; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3872 = 8'h20 == io_state_in_3 ? 8'hdb : _GEN_3871; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3873 = 8'h21 == io_state_in_3 ? 8'hd5 : _GEN_3872; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3874 = 8'h22 == io_state_in_3 ? 8'hc7 : _GEN_3873; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3875 = 8'h23 == io_state_in_3 ? 8'hc9 : _GEN_3874; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3876 = 8'h24 == io_state_in_3 ? 8'he3 : _GEN_3875; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3877 = 8'h25 == io_state_in_3 ? 8'hed : _GEN_3876; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3878 = 8'h26 == io_state_in_3 ? 8'hff : _GEN_3877; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3879 = 8'h27 == io_state_in_3 ? 8'hf1 : _GEN_3878; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3880 = 8'h28 == io_state_in_3 ? 8'hab : _GEN_3879; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3881 = 8'h29 == io_state_in_3 ? 8'ha5 : _GEN_3880; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3882 = 8'h2a == io_state_in_3 ? 8'hb7 : _GEN_3881; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3883 = 8'h2b == io_state_in_3 ? 8'hb9 : _GEN_3882; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3884 = 8'h2c == io_state_in_3 ? 8'h93 : _GEN_3883; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3885 = 8'h2d == io_state_in_3 ? 8'h9d : _GEN_3884; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3886 = 8'h2e == io_state_in_3 ? 8'h8f : _GEN_3885; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3887 = 8'h2f == io_state_in_3 ? 8'h81 : _GEN_3886; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3888 = 8'h30 == io_state_in_3 ? 8'h3b : _GEN_3887; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3889 = 8'h31 == io_state_in_3 ? 8'h35 : _GEN_3888; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3890 = 8'h32 == io_state_in_3 ? 8'h27 : _GEN_3889; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3891 = 8'h33 == io_state_in_3 ? 8'h29 : _GEN_3890; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3892 = 8'h34 == io_state_in_3 ? 8'h3 : _GEN_3891; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3893 = 8'h35 == io_state_in_3 ? 8'hd : _GEN_3892; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3894 = 8'h36 == io_state_in_3 ? 8'h1f : _GEN_3893; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3895 = 8'h37 == io_state_in_3 ? 8'h11 : _GEN_3894; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3896 = 8'h38 == io_state_in_3 ? 8'h4b : _GEN_3895; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3897 = 8'h39 == io_state_in_3 ? 8'h45 : _GEN_3896; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3898 = 8'h3a == io_state_in_3 ? 8'h57 : _GEN_3897; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3899 = 8'h3b == io_state_in_3 ? 8'h59 : _GEN_3898; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3900 = 8'h3c == io_state_in_3 ? 8'h73 : _GEN_3899; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3901 = 8'h3d == io_state_in_3 ? 8'h7d : _GEN_3900; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3902 = 8'h3e == io_state_in_3 ? 8'h6f : _GEN_3901; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3903 = 8'h3f == io_state_in_3 ? 8'h61 : _GEN_3902; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3904 = 8'h40 == io_state_in_3 ? 8'had : _GEN_3903; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3905 = 8'h41 == io_state_in_3 ? 8'ha3 : _GEN_3904; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3906 = 8'h42 == io_state_in_3 ? 8'hb1 : _GEN_3905; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3907 = 8'h43 == io_state_in_3 ? 8'hbf : _GEN_3906; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3908 = 8'h44 == io_state_in_3 ? 8'h95 : _GEN_3907; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3909 = 8'h45 == io_state_in_3 ? 8'h9b : _GEN_3908; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3910 = 8'h46 == io_state_in_3 ? 8'h89 : _GEN_3909; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3911 = 8'h47 == io_state_in_3 ? 8'h87 : _GEN_3910; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3912 = 8'h48 == io_state_in_3 ? 8'hdd : _GEN_3911; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3913 = 8'h49 == io_state_in_3 ? 8'hd3 : _GEN_3912; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3914 = 8'h4a == io_state_in_3 ? 8'hc1 : _GEN_3913; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3915 = 8'h4b == io_state_in_3 ? 8'hcf : _GEN_3914; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3916 = 8'h4c == io_state_in_3 ? 8'he5 : _GEN_3915; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3917 = 8'h4d == io_state_in_3 ? 8'heb : _GEN_3916; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3918 = 8'h4e == io_state_in_3 ? 8'hf9 : _GEN_3917; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3919 = 8'h4f == io_state_in_3 ? 8'hf7 : _GEN_3918; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3920 = 8'h50 == io_state_in_3 ? 8'h4d : _GEN_3919; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3921 = 8'h51 == io_state_in_3 ? 8'h43 : _GEN_3920; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3922 = 8'h52 == io_state_in_3 ? 8'h51 : _GEN_3921; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3923 = 8'h53 == io_state_in_3 ? 8'h5f : _GEN_3922; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3924 = 8'h54 == io_state_in_3 ? 8'h75 : _GEN_3923; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3925 = 8'h55 == io_state_in_3 ? 8'h7b : _GEN_3924; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3926 = 8'h56 == io_state_in_3 ? 8'h69 : _GEN_3925; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3927 = 8'h57 == io_state_in_3 ? 8'h67 : _GEN_3926; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3928 = 8'h58 == io_state_in_3 ? 8'h3d : _GEN_3927; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3929 = 8'h59 == io_state_in_3 ? 8'h33 : _GEN_3928; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3930 = 8'h5a == io_state_in_3 ? 8'h21 : _GEN_3929; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3931 = 8'h5b == io_state_in_3 ? 8'h2f : _GEN_3930; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3932 = 8'h5c == io_state_in_3 ? 8'h5 : _GEN_3931; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3933 = 8'h5d == io_state_in_3 ? 8'hb : _GEN_3932; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3934 = 8'h5e == io_state_in_3 ? 8'h19 : _GEN_3933; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3935 = 8'h5f == io_state_in_3 ? 8'h17 : _GEN_3934; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3936 = 8'h60 == io_state_in_3 ? 8'h76 : _GEN_3935; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3937 = 8'h61 == io_state_in_3 ? 8'h78 : _GEN_3936; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3938 = 8'h62 == io_state_in_3 ? 8'h6a : _GEN_3937; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3939 = 8'h63 == io_state_in_3 ? 8'h64 : _GEN_3938; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3940 = 8'h64 == io_state_in_3 ? 8'h4e : _GEN_3939; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3941 = 8'h65 == io_state_in_3 ? 8'h40 : _GEN_3940; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3942 = 8'h66 == io_state_in_3 ? 8'h52 : _GEN_3941; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3943 = 8'h67 == io_state_in_3 ? 8'h5c : _GEN_3942; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3944 = 8'h68 == io_state_in_3 ? 8'h6 : _GEN_3943; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3945 = 8'h69 == io_state_in_3 ? 8'h8 : _GEN_3944; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3946 = 8'h6a == io_state_in_3 ? 8'h1a : _GEN_3945; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3947 = 8'h6b == io_state_in_3 ? 8'h14 : _GEN_3946; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3948 = 8'h6c == io_state_in_3 ? 8'h3e : _GEN_3947; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3949 = 8'h6d == io_state_in_3 ? 8'h30 : _GEN_3948; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3950 = 8'h6e == io_state_in_3 ? 8'h22 : _GEN_3949; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3951 = 8'h6f == io_state_in_3 ? 8'h2c : _GEN_3950; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3952 = 8'h70 == io_state_in_3 ? 8'h96 : _GEN_3951; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3953 = 8'h71 == io_state_in_3 ? 8'h98 : _GEN_3952; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3954 = 8'h72 == io_state_in_3 ? 8'h8a : _GEN_3953; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3955 = 8'h73 == io_state_in_3 ? 8'h84 : _GEN_3954; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3956 = 8'h74 == io_state_in_3 ? 8'hae : _GEN_3955; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3957 = 8'h75 == io_state_in_3 ? 8'ha0 : _GEN_3956; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3958 = 8'h76 == io_state_in_3 ? 8'hb2 : _GEN_3957; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3959 = 8'h77 == io_state_in_3 ? 8'hbc : _GEN_3958; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3960 = 8'h78 == io_state_in_3 ? 8'he6 : _GEN_3959; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3961 = 8'h79 == io_state_in_3 ? 8'he8 : _GEN_3960; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3962 = 8'h7a == io_state_in_3 ? 8'hfa : _GEN_3961; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3963 = 8'h7b == io_state_in_3 ? 8'hf4 : _GEN_3962; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3964 = 8'h7c == io_state_in_3 ? 8'hde : _GEN_3963; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3965 = 8'h7d == io_state_in_3 ? 8'hd0 : _GEN_3964; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3966 = 8'h7e == io_state_in_3 ? 8'hc2 : _GEN_3965; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3967 = 8'h7f == io_state_in_3 ? 8'hcc : _GEN_3966; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3968 = 8'h80 == io_state_in_3 ? 8'h41 : _GEN_3967; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3969 = 8'h81 == io_state_in_3 ? 8'h4f : _GEN_3968; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3970 = 8'h82 == io_state_in_3 ? 8'h5d : _GEN_3969; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3971 = 8'h83 == io_state_in_3 ? 8'h53 : _GEN_3970; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3972 = 8'h84 == io_state_in_3 ? 8'h79 : _GEN_3971; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3973 = 8'h85 == io_state_in_3 ? 8'h77 : _GEN_3972; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3974 = 8'h86 == io_state_in_3 ? 8'h65 : _GEN_3973; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3975 = 8'h87 == io_state_in_3 ? 8'h6b : _GEN_3974; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3976 = 8'h88 == io_state_in_3 ? 8'h31 : _GEN_3975; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3977 = 8'h89 == io_state_in_3 ? 8'h3f : _GEN_3976; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3978 = 8'h8a == io_state_in_3 ? 8'h2d : _GEN_3977; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3979 = 8'h8b == io_state_in_3 ? 8'h23 : _GEN_3978; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3980 = 8'h8c == io_state_in_3 ? 8'h9 : _GEN_3979; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3981 = 8'h8d == io_state_in_3 ? 8'h7 : _GEN_3980; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3982 = 8'h8e == io_state_in_3 ? 8'h15 : _GEN_3981; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3983 = 8'h8f == io_state_in_3 ? 8'h1b : _GEN_3982; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3984 = 8'h90 == io_state_in_3 ? 8'ha1 : _GEN_3983; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3985 = 8'h91 == io_state_in_3 ? 8'haf : _GEN_3984; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3986 = 8'h92 == io_state_in_3 ? 8'hbd : _GEN_3985; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3987 = 8'h93 == io_state_in_3 ? 8'hb3 : _GEN_3986; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3988 = 8'h94 == io_state_in_3 ? 8'h99 : _GEN_3987; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3989 = 8'h95 == io_state_in_3 ? 8'h97 : _GEN_3988; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3990 = 8'h96 == io_state_in_3 ? 8'h85 : _GEN_3989; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3991 = 8'h97 == io_state_in_3 ? 8'h8b : _GEN_3990; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3992 = 8'h98 == io_state_in_3 ? 8'hd1 : _GEN_3991; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3993 = 8'h99 == io_state_in_3 ? 8'hdf : _GEN_3992; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3994 = 8'h9a == io_state_in_3 ? 8'hcd : _GEN_3993; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3995 = 8'h9b == io_state_in_3 ? 8'hc3 : _GEN_3994; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3996 = 8'h9c == io_state_in_3 ? 8'he9 : _GEN_3995; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3997 = 8'h9d == io_state_in_3 ? 8'he7 : _GEN_3996; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3998 = 8'h9e == io_state_in_3 ? 8'hf5 : _GEN_3997; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_3999 = 8'h9f == io_state_in_3 ? 8'hfb : _GEN_3998; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4000 = 8'ha0 == io_state_in_3 ? 8'h9a : _GEN_3999; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4001 = 8'ha1 == io_state_in_3 ? 8'h94 : _GEN_4000; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4002 = 8'ha2 == io_state_in_3 ? 8'h86 : _GEN_4001; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4003 = 8'ha3 == io_state_in_3 ? 8'h88 : _GEN_4002; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4004 = 8'ha4 == io_state_in_3 ? 8'ha2 : _GEN_4003; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4005 = 8'ha5 == io_state_in_3 ? 8'hac : _GEN_4004; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4006 = 8'ha6 == io_state_in_3 ? 8'hbe : _GEN_4005; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4007 = 8'ha7 == io_state_in_3 ? 8'hb0 : _GEN_4006; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4008 = 8'ha8 == io_state_in_3 ? 8'hea : _GEN_4007; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4009 = 8'ha9 == io_state_in_3 ? 8'he4 : _GEN_4008; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4010 = 8'haa == io_state_in_3 ? 8'hf6 : _GEN_4009; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4011 = 8'hab == io_state_in_3 ? 8'hf8 : _GEN_4010; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4012 = 8'hac == io_state_in_3 ? 8'hd2 : _GEN_4011; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4013 = 8'had == io_state_in_3 ? 8'hdc : _GEN_4012; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4014 = 8'hae == io_state_in_3 ? 8'hce : _GEN_4013; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4015 = 8'haf == io_state_in_3 ? 8'hc0 : _GEN_4014; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4016 = 8'hb0 == io_state_in_3 ? 8'h7a : _GEN_4015; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4017 = 8'hb1 == io_state_in_3 ? 8'h74 : _GEN_4016; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4018 = 8'hb2 == io_state_in_3 ? 8'h66 : _GEN_4017; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4019 = 8'hb3 == io_state_in_3 ? 8'h68 : _GEN_4018; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4020 = 8'hb4 == io_state_in_3 ? 8'h42 : _GEN_4019; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4021 = 8'hb5 == io_state_in_3 ? 8'h4c : _GEN_4020; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4022 = 8'hb6 == io_state_in_3 ? 8'h5e : _GEN_4021; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4023 = 8'hb7 == io_state_in_3 ? 8'h50 : _GEN_4022; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4024 = 8'hb8 == io_state_in_3 ? 8'ha : _GEN_4023; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4025 = 8'hb9 == io_state_in_3 ? 8'h4 : _GEN_4024; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4026 = 8'hba == io_state_in_3 ? 8'h16 : _GEN_4025; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4027 = 8'hbb == io_state_in_3 ? 8'h18 : _GEN_4026; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4028 = 8'hbc == io_state_in_3 ? 8'h32 : _GEN_4027; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4029 = 8'hbd == io_state_in_3 ? 8'h3c : _GEN_4028; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4030 = 8'hbe == io_state_in_3 ? 8'h2e : _GEN_4029; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4031 = 8'hbf == io_state_in_3 ? 8'h20 : _GEN_4030; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4032 = 8'hc0 == io_state_in_3 ? 8'hec : _GEN_4031; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4033 = 8'hc1 == io_state_in_3 ? 8'he2 : _GEN_4032; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4034 = 8'hc2 == io_state_in_3 ? 8'hf0 : _GEN_4033; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4035 = 8'hc3 == io_state_in_3 ? 8'hfe : _GEN_4034; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4036 = 8'hc4 == io_state_in_3 ? 8'hd4 : _GEN_4035; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4037 = 8'hc5 == io_state_in_3 ? 8'hda : _GEN_4036; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4038 = 8'hc6 == io_state_in_3 ? 8'hc8 : _GEN_4037; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4039 = 8'hc7 == io_state_in_3 ? 8'hc6 : _GEN_4038; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4040 = 8'hc8 == io_state_in_3 ? 8'h9c : _GEN_4039; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4041 = 8'hc9 == io_state_in_3 ? 8'h92 : _GEN_4040; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4042 = 8'hca == io_state_in_3 ? 8'h80 : _GEN_4041; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4043 = 8'hcb == io_state_in_3 ? 8'h8e : _GEN_4042; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4044 = 8'hcc == io_state_in_3 ? 8'ha4 : _GEN_4043; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4045 = 8'hcd == io_state_in_3 ? 8'haa : _GEN_4044; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4046 = 8'hce == io_state_in_3 ? 8'hb8 : _GEN_4045; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4047 = 8'hcf == io_state_in_3 ? 8'hb6 : _GEN_4046; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4048 = 8'hd0 == io_state_in_3 ? 8'hc : _GEN_4047; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4049 = 8'hd1 == io_state_in_3 ? 8'h2 : _GEN_4048; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4050 = 8'hd2 == io_state_in_3 ? 8'h10 : _GEN_4049; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4051 = 8'hd3 == io_state_in_3 ? 8'h1e : _GEN_4050; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4052 = 8'hd4 == io_state_in_3 ? 8'h34 : _GEN_4051; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4053 = 8'hd5 == io_state_in_3 ? 8'h3a : _GEN_4052; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4054 = 8'hd6 == io_state_in_3 ? 8'h28 : _GEN_4053; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4055 = 8'hd7 == io_state_in_3 ? 8'h26 : _GEN_4054; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4056 = 8'hd8 == io_state_in_3 ? 8'h7c : _GEN_4055; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4057 = 8'hd9 == io_state_in_3 ? 8'h72 : _GEN_4056; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4058 = 8'hda == io_state_in_3 ? 8'h60 : _GEN_4057; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4059 = 8'hdb == io_state_in_3 ? 8'h6e : _GEN_4058; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4060 = 8'hdc == io_state_in_3 ? 8'h44 : _GEN_4059; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4061 = 8'hdd == io_state_in_3 ? 8'h4a : _GEN_4060; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4062 = 8'hde == io_state_in_3 ? 8'h58 : _GEN_4061; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4063 = 8'hdf == io_state_in_3 ? 8'h56 : _GEN_4062; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4064 = 8'he0 == io_state_in_3 ? 8'h37 : _GEN_4063; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4065 = 8'he1 == io_state_in_3 ? 8'h39 : _GEN_4064; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4066 = 8'he2 == io_state_in_3 ? 8'h2b : _GEN_4065; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4067 = 8'he3 == io_state_in_3 ? 8'h25 : _GEN_4066; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4068 = 8'he4 == io_state_in_3 ? 8'hf : _GEN_4067; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4069 = 8'he5 == io_state_in_3 ? 8'h1 : _GEN_4068; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4070 = 8'he6 == io_state_in_3 ? 8'h13 : _GEN_4069; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4071 = 8'he7 == io_state_in_3 ? 8'h1d : _GEN_4070; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4072 = 8'he8 == io_state_in_3 ? 8'h47 : _GEN_4071; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4073 = 8'he9 == io_state_in_3 ? 8'h49 : _GEN_4072; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4074 = 8'hea == io_state_in_3 ? 8'h5b : _GEN_4073; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4075 = 8'heb == io_state_in_3 ? 8'h55 : _GEN_4074; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4076 = 8'hec == io_state_in_3 ? 8'h7f : _GEN_4075; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4077 = 8'hed == io_state_in_3 ? 8'h71 : _GEN_4076; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4078 = 8'hee == io_state_in_3 ? 8'h63 : _GEN_4077; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4079 = 8'hef == io_state_in_3 ? 8'h6d : _GEN_4078; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4080 = 8'hf0 == io_state_in_3 ? 8'hd7 : _GEN_4079; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4081 = 8'hf1 == io_state_in_3 ? 8'hd9 : _GEN_4080; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4082 = 8'hf2 == io_state_in_3 ? 8'hcb : _GEN_4081; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4083 = 8'hf3 == io_state_in_3 ? 8'hc5 : _GEN_4082; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4084 = 8'hf4 == io_state_in_3 ? 8'hef : _GEN_4083; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4085 = 8'hf5 == io_state_in_3 ? 8'he1 : _GEN_4084; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4086 = 8'hf6 == io_state_in_3 ? 8'hf3 : _GEN_4085; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4087 = 8'hf7 == io_state_in_3 ? 8'hfd : _GEN_4086; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4088 = 8'hf8 == io_state_in_3 ? 8'ha7 : _GEN_4087; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4089 = 8'hf9 == io_state_in_3 ? 8'ha9 : _GEN_4088; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4090 = 8'hfa == io_state_in_3 ? 8'hbb : _GEN_4089; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4091 = 8'hfb == io_state_in_3 ? 8'hb5 : _GEN_4090; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4092 = 8'hfc == io_state_in_3 ? 8'h9f : _GEN_4091; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4093 = 8'hfd == io_state_in_3 ? 8'h91 : _GEN_4092; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4094 = 8'hfe == io_state_in_3 ? 8'h83 : _GEN_4093; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4095 = 8'hff == io_state_in_3 ? 8'h8d : _GEN_4094; // @[InvMixColumns.scala 129:{89,89}]
  wire [7:0] _GEN_4097 = 8'h1 == io_state_in_4 ? 8'he : 8'h0; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4098 = 8'h2 == io_state_in_4 ? 8'h1c : _GEN_4097; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4099 = 8'h3 == io_state_in_4 ? 8'h12 : _GEN_4098; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4100 = 8'h4 == io_state_in_4 ? 8'h38 : _GEN_4099; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4101 = 8'h5 == io_state_in_4 ? 8'h36 : _GEN_4100; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4102 = 8'h6 == io_state_in_4 ? 8'h24 : _GEN_4101; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4103 = 8'h7 == io_state_in_4 ? 8'h2a : _GEN_4102; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4104 = 8'h8 == io_state_in_4 ? 8'h70 : _GEN_4103; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4105 = 8'h9 == io_state_in_4 ? 8'h7e : _GEN_4104; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4106 = 8'ha == io_state_in_4 ? 8'h6c : _GEN_4105; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4107 = 8'hb == io_state_in_4 ? 8'h62 : _GEN_4106; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4108 = 8'hc == io_state_in_4 ? 8'h48 : _GEN_4107; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4109 = 8'hd == io_state_in_4 ? 8'h46 : _GEN_4108; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4110 = 8'he == io_state_in_4 ? 8'h54 : _GEN_4109; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4111 = 8'hf == io_state_in_4 ? 8'h5a : _GEN_4110; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4112 = 8'h10 == io_state_in_4 ? 8'he0 : _GEN_4111; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4113 = 8'h11 == io_state_in_4 ? 8'hee : _GEN_4112; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4114 = 8'h12 == io_state_in_4 ? 8'hfc : _GEN_4113; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4115 = 8'h13 == io_state_in_4 ? 8'hf2 : _GEN_4114; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4116 = 8'h14 == io_state_in_4 ? 8'hd8 : _GEN_4115; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4117 = 8'h15 == io_state_in_4 ? 8'hd6 : _GEN_4116; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4118 = 8'h16 == io_state_in_4 ? 8'hc4 : _GEN_4117; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4119 = 8'h17 == io_state_in_4 ? 8'hca : _GEN_4118; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4120 = 8'h18 == io_state_in_4 ? 8'h90 : _GEN_4119; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4121 = 8'h19 == io_state_in_4 ? 8'h9e : _GEN_4120; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4122 = 8'h1a == io_state_in_4 ? 8'h8c : _GEN_4121; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4123 = 8'h1b == io_state_in_4 ? 8'h82 : _GEN_4122; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4124 = 8'h1c == io_state_in_4 ? 8'ha8 : _GEN_4123; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4125 = 8'h1d == io_state_in_4 ? 8'ha6 : _GEN_4124; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4126 = 8'h1e == io_state_in_4 ? 8'hb4 : _GEN_4125; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4127 = 8'h1f == io_state_in_4 ? 8'hba : _GEN_4126; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4128 = 8'h20 == io_state_in_4 ? 8'hdb : _GEN_4127; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4129 = 8'h21 == io_state_in_4 ? 8'hd5 : _GEN_4128; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4130 = 8'h22 == io_state_in_4 ? 8'hc7 : _GEN_4129; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4131 = 8'h23 == io_state_in_4 ? 8'hc9 : _GEN_4130; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4132 = 8'h24 == io_state_in_4 ? 8'he3 : _GEN_4131; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4133 = 8'h25 == io_state_in_4 ? 8'hed : _GEN_4132; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4134 = 8'h26 == io_state_in_4 ? 8'hff : _GEN_4133; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4135 = 8'h27 == io_state_in_4 ? 8'hf1 : _GEN_4134; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4136 = 8'h28 == io_state_in_4 ? 8'hab : _GEN_4135; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4137 = 8'h29 == io_state_in_4 ? 8'ha5 : _GEN_4136; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4138 = 8'h2a == io_state_in_4 ? 8'hb7 : _GEN_4137; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4139 = 8'h2b == io_state_in_4 ? 8'hb9 : _GEN_4138; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4140 = 8'h2c == io_state_in_4 ? 8'h93 : _GEN_4139; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4141 = 8'h2d == io_state_in_4 ? 8'h9d : _GEN_4140; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4142 = 8'h2e == io_state_in_4 ? 8'h8f : _GEN_4141; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4143 = 8'h2f == io_state_in_4 ? 8'h81 : _GEN_4142; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4144 = 8'h30 == io_state_in_4 ? 8'h3b : _GEN_4143; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4145 = 8'h31 == io_state_in_4 ? 8'h35 : _GEN_4144; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4146 = 8'h32 == io_state_in_4 ? 8'h27 : _GEN_4145; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4147 = 8'h33 == io_state_in_4 ? 8'h29 : _GEN_4146; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4148 = 8'h34 == io_state_in_4 ? 8'h3 : _GEN_4147; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4149 = 8'h35 == io_state_in_4 ? 8'hd : _GEN_4148; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4150 = 8'h36 == io_state_in_4 ? 8'h1f : _GEN_4149; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4151 = 8'h37 == io_state_in_4 ? 8'h11 : _GEN_4150; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4152 = 8'h38 == io_state_in_4 ? 8'h4b : _GEN_4151; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4153 = 8'h39 == io_state_in_4 ? 8'h45 : _GEN_4152; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4154 = 8'h3a == io_state_in_4 ? 8'h57 : _GEN_4153; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4155 = 8'h3b == io_state_in_4 ? 8'h59 : _GEN_4154; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4156 = 8'h3c == io_state_in_4 ? 8'h73 : _GEN_4155; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4157 = 8'h3d == io_state_in_4 ? 8'h7d : _GEN_4156; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4158 = 8'h3e == io_state_in_4 ? 8'h6f : _GEN_4157; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4159 = 8'h3f == io_state_in_4 ? 8'h61 : _GEN_4158; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4160 = 8'h40 == io_state_in_4 ? 8'had : _GEN_4159; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4161 = 8'h41 == io_state_in_4 ? 8'ha3 : _GEN_4160; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4162 = 8'h42 == io_state_in_4 ? 8'hb1 : _GEN_4161; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4163 = 8'h43 == io_state_in_4 ? 8'hbf : _GEN_4162; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4164 = 8'h44 == io_state_in_4 ? 8'h95 : _GEN_4163; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4165 = 8'h45 == io_state_in_4 ? 8'h9b : _GEN_4164; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4166 = 8'h46 == io_state_in_4 ? 8'h89 : _GEN_4165; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4167 = 8'h47 == io_state_in_4 ? 8'h87 : _GEN_4166; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4168 = 8'h48 == io_state_in_4 ? 8'hdd : _GEN_4167; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4169 = 8'h49 == io_state_in_4 ? 8'hd3 : _GEN_4168; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4170 = 8'h4a == io_state_in_4 ? 8'hc1 : _GEN_4169; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4171 = 8'h4b == io_state_in_4 ? 8'hcf : _GEN_4170; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4172 = 8'h4c == io_state_in_4 ? 8'he5 : _GEN_4171; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4173 = 8'h4d == io_state_in_4 ? 8'heb : _GEN_4172; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4174 = 8'h4e == io_state_in_4 ? 8'hf9 : _GEN_4173; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4175 = 8'h4f == io_state_in_4 ? 8'hf7 : _GEN_4174; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4176 = 8'h50 == io_state_in_4 ? 8'h4d : _GEN_4175; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4177 = 8'h51 == io_state_in_4 ? 8'h43 : _GEN_4176; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4178 = 8'h52 == io_state_in_4 ? 8'h51 : _GEN_4177; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4179 = 8'h53 == io_state_in_4 ? 8'h5f : _GEN_4178; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4180 = 8'h54 == io_state_in_4 ? 8'h75 : _GEN_4179; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4181 = 8'h55 == io_state_in_4 ? 8'h7b : _GEN_4180; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4182 = 8'h56 == io_state_in_4 ? 8'h69 : _GEN_4181; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4183 = 8'h57 == io_state_in_4 ? 8'h67 : _GEN_4182; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4184 = 8'h58 == io_state_in_4 ? 8'h3d : _GEN_4183; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4185 = 8'h59 == io_state_in_4 ? 8'h33 : _GEN_4184; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4186 = 8'h5a == io_state_in_4 ? 8'h21 : _GEN_4185; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4187 = 8'h5b == io_state_in_4 ? 8'h2f : _GEN_4186; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4188 = 8'h5c == io_state_in_4 ? 8'h5 : _GEN_4187; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4189 = 8'h5d == io_state_in_4 ? 8'hb : _GEN_4188; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4190 = 8'h5e == io_state_in_4 ? 8'h19 : _GEN_4189; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4191 = 8'h5f == io_state_in_4 ? 8'h17 : _GEN_4190; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4192 = 8'h60 == io_state_in_4 ? 8'h76 : _GEN_4191; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4193 = 8'h61 == io_state_in_4 ? 8'h78 : _GEN_4192; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4194 = 8'h62 == io_state_in_4 ? 8'h6a : _GEN_4193; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4195 = 8'h63 == io_state_in_4 ? 8'h64 : _GEN_4194; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4196 = 8'h64 == io_state_in_4 ? 8'h4e : _GEN_4195; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4197 = 8'h65 == io_state_in_4 ? 8'h40 : _GEN_4196; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4198 = 8'h66 == io_state_in_4 ? 8'h52 : _GEN_4197; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4199 = 8'h67 == io_state_in_4 ? 8'h5c : _GEN_4198; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4200 = 8'h68 == io_state_in_4 ? 8'h6 : _GEN_4199; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4201 = 8'h69 == io_state_in_4 ? 8'h8 : _GEN_4200; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4202 = 8'h6a == io_state_in_4 ? 8'h1a : _GEN_4201; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4203 = 8'h6b == io_state_in_4 ? 8'h14 : _GEN_4202; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4204 = 8'h6c == io_state_in_4 ? 8'h3e : _GEN_4203; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4205 = 8'h6d == io_state_in_4 ? 8'h30 : _GEN_4204; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4206 = 8'h6e == io_state_in_4 ? 8'h22 : _GEN_4205; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4207 = 8'h6f == io_state_in_4 ? 8'h2c : _GEN_4206; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4208 = 8'h70 == io_state_in_4 ? 8'h96 : _GEN_4207; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4209 = 8'h71 == io_state_in_4 ? 8'h98 : _GEN_4208; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4210 = 8'h72 == io_state_in_4 ? 8'h8a : _GEN_4209; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4211 = 8'h73 == io_state_in_4 ? 8'h84 : _GEN_4210; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4212 = 8'h74 == io_state_in_4 ? 8'hae : _GEN_4211; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4213 = 8'h75 == io_state_in_4 ? 8'ha0 : _GEN_4212; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4214 = 8'h76 == io_state_in_4 ? 8'hb2 : _GEN_4213; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4215 = 8'h77 == io_state_in_4 ? 8'hbc : _GEN_4214; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4216 = 8'h78 == io_state_in_4 ? 8'he6 : _GEN_4215; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4217 = 8'h79 == io_state_in_4 ? 8'he8 : _GEN_4216; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4218 = 8'h7a == io_state_in_4 ? 8'hfa : _GEN_4217; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4219 = 8'h7b == io_state_in_4 ? 8'hf4 : _GEN_4218; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4220 = 8'h7c == io_state_in_4 ? 8'hde : _GEN_4219; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4221 = 8'h7d == io_state_in_4 ? 8'hd0 : _GEN_4220; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4222 = 8'h7e == io_state_in_4 ? 8'hc2 : _GEN_4221; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4223 = 8'h7f == io_state_in_4 ? 8'hcc : _GEN_4222; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4224 = 8'h80 == io_state_in_4 ? 8'h41 : _GEN_4223; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4225 = 8'h81 == io_state_in_4 ? 8'h4f : _GEN_4224; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4226 = 8'h82 == io_state_in_4 ? 8'h5d : _GEN_4225; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4227 = 8'h83 == io_state_in_4 ? 8'h53 : _GEN_4226; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4228 = 8'h84 == io_state_in_4 ? 8'h79 : _GEN_4227; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4229 = 8'h85 == io_state_in_4 ? 8'h77 : _GEN_4228; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4230 = 8'h86 == io_state_in_4 ? 8'h65 : _GEN_4229; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4231 = 8'h87 == io_state_in_4 ? 8'h6b : _GEN_4230; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4232 = 8'h88 == io_state_in_4 ? 8'h31 : _GEN_4231; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4233 = 8'h89 == io_state_in_4 ? 8'h3f : _GEN_4232; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4234 = 8'h8a == io_state_in_4 ? 8'h2d : _GEN_4233; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4235 = 8'h8b == io_state_in_4 ? 8'h23 : _GEN_4234; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4236 = 8'h8c == io_state_in_4 ? 8'h9 : _GEN_4235; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4237 = 8'h8d == io_state_in_4 ? 8'h7 : _GEN_4236; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4238 = 8'h8e == io_state_in_4 ? 8'h15 : _GEN_4237; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4239 = 8'h8f == io_state_in_4 ? 8'h1b : _GEN_4238; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4240 = 8'h90 == io_state_in_4 ? 8'ha1 : _GEN_4239; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4241 = 8'h91 == io_state_in_4 ? 8'haf : _GEN_4240; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4242 = 8'h92 == io_state_in_4 ? 8'hbd : _GEN_4241; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4243 = 8'h93 == io_state_in_4 ? 8'hb3 : _GEN_4242; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4244 = 8'h94 == io_state_in_4 ? 8'h99 : _GEN_4243; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4245 = 8'h95 == io_state_in_4 ? 8'h97 : _GEN_4244; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4246 = 8'h96 == io_state_in_4 ? 8'h85 : _GEN_4245; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4247 = 8'h97 == io_state_in_4 ? 8'h8b : _GEN_4246; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4248 = 8'h98 == io_state_in_4 ? 8'hd1 : _GEN_4247; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4249 = 8'h99 == io_state_in_4 ? 8'hdf : _GEN_4248; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4250 = 8'h9a == io_state_in_4 ? 8'hcd : _GEN_4249; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4251 = 8'h9b == io_state_in_4 ? 8'hc3 : _GEN_4250; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4252 = 8'h9c == io_state_in_4 ? 8'he9 : _GEN_4251; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4253 = 8'h9d == io_state_in_4 ? 8'he7 : _GEN_4252; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4254 = 8'h9e == io_state_in_4 ? 8'hf5 : _GEN_4253; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4255 = 8'h9f == io_state_in_4 ? 8'hfb : _GEN_4254; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4256 = 8'ha0 == io_state_in_4 ? 8'h9a : _GEN_4255; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4257 = 8'ha1 == io_state_in_4 ? 8'h94 : _GEN_4256; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4258 = 8'ha2 == io_state_in_4 ? 8'h86 : _GEN_4257; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4259 = 8'ha3 == io_state_in_4 ? 8'h88 : _GEN_4258; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4260 = 8'ha4 == io_state_in_4 ? 8'ha2 : _GEN_4259; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4261 = 8'ha5 == io_state_in_4 ? 8'hac : _GEN_4260; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4262 = 8'ha6 == io_state_in_4 ? 8'hbe : _GEN_4261; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4263 = 8'ha7 == io_state_in_4 ? 8'hb0 : _GEN_4262; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4264 = 8'ha8 == io_state_in_4 ? 8'hea : _GEN_4263; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4265 = 8'ha9 == io_state_in_4 ? 8'he4 : _GEN_4264; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4266 = 8'haa == io_state_in_4 ? 8'hf6 : _GEN_4265; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4267 = 8'hab == io_state_in_4 ? 8'hf8 : _GEN_4266; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4268 = 8'hac == io_state_in_4 ? 8'hd2 : _GEN_4267; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4269 = 8'had == io_state_in_4 ? 8'hdc : _GEN_4268; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4270 = 8'hae == io_state_in_4 ? 8'hce : _GEN_4269; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4271 = 8'haf == io_state_in_4 ? 8'hc0 : _GEN_4270; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4272 = 8'hb0 == io_state_in_4 ? 8'h7a : _GEN_4271; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4273 = 8'hb1 == io_state_in_4 ? 8'h74 : _GEN_4272; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4274 = 8'hb2 == io_state_in_4 ? 8'h66 : _GEN_4273; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4275 = 8'hb3 == io_state_in_4 ? 8'h68 : _GEN_4274; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4276 = 8'hb4 == io_state_in_4 ? 8'h42 : _GEN_4275; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4277 = 8'hb5 == io_state_in_4 ? 8'h4c : _GEN_4276; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4278 = 8'hb6 == io_state_in_4 ? 8'h5e : _GEN_4277; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4279 = 8'hb7 == io_state_in_4 ? 8'h50 : _GEN_4278; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4280 = 8'hb8 == io_state_in_4 ? 8'ha : _GEN_4279; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4281 = 8'hb9 == io_state_in_4 ? 8'h4 : _GEN_4280; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4282 = 8'hba == io_state_in_4 ? 8'h16 : _GEN_4281; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4283 = 8'hbb == io_state_in_4 ? 8'h18 : _GEN_4282; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4284 = 8'hbc == io_state_in_4 ? 8'h32 : _GEN_4283; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4285 = 8'hbd == io_state_in_4 ? 8'h3c : _GEN_4284; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4286 = 8'hbe == io_state_in_4 ? 8'h2e : _GEN_4285; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4287 = 8'hbf == io_state_in_4 ? 8'h20 : _GEN_4286; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4288 = 8'hc0 == io_state_in_4 ? 8'hec : _GEN_4287; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4289 = 8'hc1 == io_state_in_4 ? 8'he2 : _GEN_4288; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4290 = 8'hc2 == io_state_in_4 ? 8'hf0 : _GEN_4289; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4291 = 8'hc3 == io_state_in_4 ? 8'hfe : _GEN_4290; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4292 = 8'hc4 == io_state_in_4 ? 8'hd4 : _GEN_4291; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4293 = 8'hc5 == io_state_in_4 ? 8'hda : _GEN_4292; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4294 = 8'hc6 == io_state_in_4 ? 8'hc8 : _GEN_4293; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4295 = 8'hc7 == io_state_in_4 ? 8'hc6 : _GEN_4294; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4296 = 8'hc8 == io_state_in_4 ? 8'h9c : _GEN_4295; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4297 = 8'hc9 == io_state_in_4 ? 8'h92 : _GEN_4296; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4298 = 8'hca == io_state_in_4 ? 8'h80 : _GEN_4297; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4299 = 8'hcb == io_state_in_4 ? 8'h8e : _GEN_4298; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4300 = 8'hcc == io_state_in_4 ? 8'ha4 : _GEN_4299; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4301 = 8'hcd == io_state_in_4 ? 8'haa : _GEN_4300; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4302 = 8'hce == io_state_in_4 ? 8'hb8 : _GEN_4301; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4303 = 8'hcf == io_state_in_4 ? 8'hb6 : _GEN_4302; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4304 = 8'hd0 == io_state_in_4 ? 8'hc : _GEN_4303; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4305 = 8'hd1 == io_state_in_4 ? 8'h2 : _GEN_4304; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4306 = 8'hd2 == io_state_in_4 ? 8'h10 : _GEN_4305; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4307 = 8'hd3 == io_state_in_4 ? 8'h1e : _GEN_4306; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4308 = 8'hd4 == io_state_in_4 ? 8'h34 : _GEN_4307; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4309 = 8'hd5 == io_state_in_4 ? 8'h3a : _GEN_4308; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4310 = 8'hd6 == io_state_in_4 ? 8'h28 : _GEN_4309; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4311 = 8'hd7 == io_state_in_4 ? 8'h26 : _GEN_4310; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4312 = 8'hd8 == io_state_in_4 ? 8'h7c : _GEN_4311; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4313 = 8'hd9 == io_state_in_4 ? 8'h72 : _GEN_4312; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4314 = 8'hda == io_state_in_4 ? 8'h60 : _GEN_4313; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4315 = 8'hdb == io_state_in_4 ? 8'h6e : _GEN_4314; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4316 = 8'hdc == io_state_in_4 ? 8'h44 : _GEN_4315; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4317 = 8'hdd == io_state_in_4 ? 8'h4a : _GEN_4316; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4318 = 8'hde == io_state_in_4 ? 8'h58 : _GEN_4317; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4319 = 8'hdf == io_state_in_4 ? 8'h56 : _GEN_4318; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4320 = 8'he0 == io_state_in_4 ? 8'h37 : _GEN_4319; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4321 = 8'he1 == io_state_in_4 ? 8'h39 : _GEN_4320; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4322 = 8'he2 == io_state_in_4 ? 8'h2b : _GEN_4321; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4323 = 8'he3 == io_state_in_4 ? 8'h25 : _GEN_4322; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4324 = 8'he4 == io_state_in_4 ? 8'hf : _GEN_4323; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4325 = 8'he5 == io_state_in_4 ? 8'h1 : _GEN_4324; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4326 = 8'he6 == io_state_in_4 ? 8'h13 : _GEN_4325; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4327 = 8'he7 == io_state_in_4 ? 8'h1d : _GEN_4326; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4328 = 8'he8 == io_state_in_4 ? 8'h47 : _GEN_4327; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4329 = 8'he9 == io_state_in_4 ? 8'h49 : _GEN_4328; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4330 = 8'hea == io_state_in_4 ? 8'h5b : _GEN_4329; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4331 = 8'heb == io_state_in_4 ? 8'h55 : _GEN_4330; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4332 = 8'hec == io_state_in_4 ? 8'h7f : _GEN_4331; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4333 = 8'hed == io_state_in_4 ? 8'h71 : _GEN_4332; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4334 = 8'hee == io_state_in_4 ? 8'h63 : _GEN_4333; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4335 = 8'hef == io_state_in_4 ? 8'h6d : _GEN_4334; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4336 = 8'hf0 == io_state_in_4 ? 8'hd7 : _GEN_4335; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4337 = 8'hf1 == io_state_in_4 ? 8'hd9 : _GEN_4336; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4338 = 8'hf2 == io_state_in_4 ? 8'hcb : _GEN_4337; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4339 = 8'hf3 == io_state_in_4 ? 8'hc5 : _GEN_4338; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4340 = 8'hf4 == io_state_in_4 ? 8'hef : _GEN_4339; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4341 = 8'hf5 == io_state_in_4 ? 8'he1 : _GEN_4340; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4342 = 8'hf6 == io_state_in_4 ? 8'hf3 : _GEN_4341; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4343 = 8'hf7 == io_state_in_4 ? 8'hfd : _GEN_4342; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4344 = 8'hf8 == io_state_in_4 ? 8'ha7 : _GEN_4343; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4345 = 8'hf9 == io_state_in_4 ? 8'ha9 : _GEN_4344; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4346 = 8'hfa == io_state_in_4 ? 8'hbb : _GEN_4345; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4347 = 8'hfb == io_state_in_4 ? 8'hb5 : _GEN_4346; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4348 = 8'hfc == io_state_in_4 ? 8'h9f : _GEN_4347; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4349 = 8'hfd == io_state_in_4 ? 8'h91 : _GEN_4348; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4350 = 8'hfe == io_state_in_4 ? 8'h83 : _GEN_4349; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4351 = 8'hff == io_state_in_4 ? 8'h8d : _GEN_4350; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4353 = 8'h1 == io_state_in_5 ? 8'hb : 8'h0; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4354 = 8'h2 == io_state_in_5 ? 8'h16 : _GEN_4353; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4355 = 8'h3 == io_state_in_5 ? 8'h1d : _GEN_4354; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4356 = 8'h4 == io_state_in_5 ? 8'h2c : _GEN_4355; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4357 = 8'h5 == io_state_in_5 ? 8'h27 : _GEN_4356; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4358 = 8'h6 == io_state_in_5 ? 8'h3a : _GEN_4357; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4359 = 8'h7 == io_state_in_5 ? 8'h31 : _GEN_4358; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4360 = 8'h8 == io_state_in_5 ? 8'h58 : _GEN_4359; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4361 = 8'h9 == io_state_in_5 ? 8'h53 : _GEN_4360; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4362 = 8'ha == io_state_in_5 ? 8'h4e : _GEN_4361; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4363 = 8'hb == io_state_in_5 ? 8'h45 : _GEN_4362; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4364 = 8'hc == io_state_in_5 ? 8'h74 : _GEN_4363; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4365 = 8'hd == io_state_in_5 ? 8'h7f : _GEN_4364; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4366 = 8'he == io_state_in_5 ? 8'h62 : _GEN_4365; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4367 = 8'hf == io_state_in_5 ? 8'h69 : _GEN_4366; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4368 = 8'h10 == io_state_in_5 ? 8'hb0 : _GEN_4367; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4369 = 8'h11 == io_state_in_5 ? 8'hbb : _GEN_4368; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4370 = 8'h12 == io_state_in_5 ? 8'ha6 : _GEN_4369; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4371 = 8'h13 == io_state_in_5 ? 8'had : _GEN_4370; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4372 = 8'h14 == io_state_in_5 ? 8'h9c : _GEN_4371; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4373 = 8'h15 == io_state_in_5 ? 8'h97 : _GEN_4372; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4374 = 8'h16 == io_state_in_5 ? 8'h8a : _GEN_4373; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4375 = 8'h17 == io_state_in_5 ? 8'h81 : _GEN_4374; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4376 = 8'h18 == io_state_in_5 ? 8'he8 : _GEN_4375; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4377 = 8'h19 == io_state_in_5 ? 8'he3 : _GEN_4376; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4378 = 8'h1a == io_state_in_5 ? 8'hfe : _GEN_4377; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4379 = 8'h1b == io_state_in_5 ? 8'hf5 : _GEN_4378; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4380 = 8'h1c == io_state_in_5 ? 8'hc4 : _GEN_4379; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4381 = 8'h1d == io_state_in_5 ? 8'hcf : _GEN_4380; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4382 = 8'h1e == io_state_in_5 ? 8'hd2 : _GEN_4381; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4383 = 8'h1f == io_state_in_5 ? 8'hd9 : _GEN_4382; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4384 = 8'h20 == io_state_in_5 ? 8'h7b : _GEN_4383; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4385 = 8'h21 == io_state_in_5 ? 8'h70 : _GEN_4384; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4386 = 8'h22 == io_state_in_5 ? 8'h6d : _GEN_4385; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4387 = 8'h23 == io_state_in_5 ? 8'h66 : _GEN_4386; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4388 = 8'h24 == io_state_in_5 ? 8'h57 : _GEN_4387; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4389 = 8'h25 == io_state_in_5 ? 8'h5c : _GEN_4388; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4390 = 8'h26 == io_state_in_5 ? 8'h41 : _GEN_4389; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4391 = 8'h27 == io_state_in_5 ? 8'h4a : _GEN_4390; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4392 = 8'h28 == io_state_in_5 ? 8'h23 : _GEN_4391; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4393 = 8'h29 == io_state_in_5 ? 8'h28 : _GEN_4392; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4394 = 8'h2a == io_state_in_5 ? 8'h35 : _GEN_4393; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4395 = 8'h2b == io_state_in_5 ? 8'h3e : _GEN_4394; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4396 = 8'h2c == io_state_in_5 ? 8'hf : _GEN_4395; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4397 = 8'h2d == io_state_in_5 ? 8'h4 : _GEN_4396; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4398 = 8'h2e == io_state_in_5 ? 8'h19 : _GEN_4397; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4399 = 8'h2f == io_state_in_5 ? 8'h12 : _GEN_4398; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4400 = 8'h30 == io_state_in_5 ? 8'hcb : _GEN_4399; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4401 = 8'h31 == io_state_in_5 ? 8'hc0 : _GEN_4400; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4402 = 8'h32 == io_state_in_5 ? 8'hdd : _GEN_4401; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4403 = 8'h33 == io_state_in_5 ? 8'hd6 : _GEN_4402; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4404 = 8'h34 == io_state_in_5 ? 8'he7 : _GEN_4403; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4405 = 8'h35 == io_state_in_5 ? 8'hec : _GEN_4404; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4406 = 8'h36 == io_state_in_5 ? 8'hf1 : _GEN_4405; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4407 = 8'h37 == io_state_in_5 ? 8'hfa : _GEN_4406; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4408 = 8'h38 == io_state_in_5 ? 8'h93 : _GEN_4407; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4409 = 8'h39 == io_state_in_5 ? 8'h98 : _GEN_4408; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4410 = 8'h3a == io_state_in_5 ? 8'h85 : _GEN_4409; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4411 = 8'h3b == io_state_in_5 ? 8'h8e : _GEN_4410; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4412 = 8'h3c == io_state_in_5 ? 8'hbf : _GEN_4411; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4413 = 8'h3d == io_state_in_5 ? 8'hb4 : _GEN_4412; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4414 = 8'h3e == io_state_in_5 ? 8'ha9 : _GEN_4413; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4415 = 8'h3f == io_state_in_5 ? 8'ha2 : _GEN_4414; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4416 = 8'h40 == io_state_in_5 ? 8'hf6 : _GEN_4415; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4417 = 8'h41 == io_state_in_5 ? 8'hfd : _GEN_4416; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4418 = 8'h42 == io_state_in_5 ? 8'he0 : _GEN_4417; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4419 = 8'h43 == io_state_in_5 ? 8'heb : _GEN_4418; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4420 = 8'h44 == io_state_in_5 ? 8'hda : _GEN_4419; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4421 = 8'h45 == io_state_in_5 ? 8'hd1 : _GEN_4420; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4422 = 8'h46 == io_state_in_5 ? 8'hcc : _GEN_4421; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4423 = 8'h47 == io_state_in_5 ? 8'hc7 : _GEN_4422; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4424 = 8'h48 == io_state_in_5 ? 8'hae : _GEN_4423; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4425 = 8'h49 == io_state_in_5 ? 8'ha5 : _GEN_4424; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4426 = 8'h4a == io_state_in_5 ? 8'hb8 : _GEN_4425; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4427 = 8'h4b == io_state_in_5 ? 8'hb3 : _GEN_4426; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4428 = 8'h4c == io_state_in_5 ? 8'h82 : _GEN_4427; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4429 = 8'h4d == io_state_in_5 ? 8'h89 : _GEN_4428; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4430 = 8'h4e == io_state_in_5 ? 8'h94 : _GEN_4429; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4431 = 8'h4f == io_state_in_5 ? 8'h9f : _GEN_4430; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4432 = 8'h50 == io_state_in_5 ? 8'h46 : _GEN_4431; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4433 = 8'h51 == io_state_in_5 ? 8'h4d : _GEN_4432; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4434 = 8'h52 == io_state_in_5 ? 8'h50 : _GEN_4433; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4435 = 8'h53 == io_state_in_5 ? 8'h5b : _GEN_4434; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4436 = 8'h54 == io_state_in_5 ? 8'h6a : _GEN_4435; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4437 = 8'h55 == io_state_in_5 ? 8'h61 : _GEN_4436; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4438 = 8'h56 == io_state_in_5 ? 8'h7c : _GEN_4437; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4439 = 8'h57 == io_state_in_5 ? 8'h77 : _GEN_4438; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4440 = 8'h58 == io_state_in_5 ? 8'h1e : _GEN_4439; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4441 = 8'h59 == io_state_in_5 ? 8'h15 : _GEN_4440; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4442 = 8'h5a == io_state_in_5 ? 8'h8 : _GEN_4441; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4443 = 8'h5b == io_state_in_5 ? 8'h3 : _GEN_4442; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4444 = 8'h5c == io_state_in_5 ? 8'h32 : _GEN_4443; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4445 = 8'h5d == io_state_in_5 ? 8'h39 : _GEN_4444; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4446 = 8'h5e == io_state_in_5 ? 8'h24 : _GEN_4445; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4447 = 8'h5f == io_state_in_5 ? 8'h2f : _GEN_4446; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4448 = 8'h60 == io_state_in_5 ? 8'h8d : _GEN_4447; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4449 = 8'h61 == io_state_in_5 ? 8'h86 : _GEN_4448; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4450 = 8'h62 == io_state_in_5 ? 8'h9b : _GEN_4449; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4451 = 8'h63 == io_state_in_5 ? 8'h90 : _GEN_4450; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4452 = 8'h64 == io_state_in_5 ? 8'ha1 : _GEN_4451; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4453 = 8'h65 == io_state_in_5 ? 8'haa : _GEN_4452; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4454 = 8'h66 == io_state_in_5 ? 8'hb7 : _GEN_4453; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4455 = 8'h67 == io_state_in_5 ? 8'hbc : _GEN_4454; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4456 = 8'h68 == io_state_in_5 ? 8'hd5 : _GEN_4455; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4457 = 8'h69 == io_state_in_5 ? 8'hde : _GEN_4456; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4458 = 8'h6a == io_state_in_5 ? 8'hc3 : _GEN_4457; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4459 = 8'h6b == io_state_in_5 ? 8'hc8 : _GEN_4458; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4460 = 8'h6c == io_state_in_5 ? 8'hf9 : _GEN_4459; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4461 = 8'h6d == io_state_in_5 ? 8'hf2 : _GEN_4460; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4462 = 8'h6e == io_state_in_5 ? 8'hef : _GEN_4461; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4463 = 8'h6f == io_state_in_5 ? 8'he4 : _GEN_4462; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4464 = 8'h70 == io_state_in_5 ? 8'h3d : _GEN_4463; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4465 = 8'h71 == io_state_in_5 ? 8'h36 : _GEN_4464; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4466 = 8'h72 == io_state_in_5 ? 8'h2b : _GEN_4465; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4467 = 8'h73 == io_state_in_5 ? 8'h20 : _GEN_4466; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4468 = 8'h74 == io_state_in_5 ? 8'h11 : _GEN_4467; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4469 = 8'h75 == io_state_in_5 ? 8'h1a : _GEN_4468; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4470 = 8'h76 == io_state_in_5 ? 8'h7 : _GEN_4469; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4471 = 8'h77 == io_state_in_5 ? 8'hc : _GEN_4470; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4472 = 8'h78 == io_state_in_5 ? 8'h65 : _GEN_4471; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4473 = 8'h79 == io_state_in_5 ? 8'h6e : _GEN_4472; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4474 = 8'h7a == io_state_in_5 ? 8'h73 : _GEN_4473; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4475 = 8'h7b == io_state_in_5 ? 8'h78 : _GEN_4474; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4476 = 8'h7c == io_state_in_5 ? 8'h49 : _GEN_4475; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4477 = 8'h7d == io_state_in_5 ? 8'h42 : _GEN_4476; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4478 = 8'h7e == io_state_in_5 ? 8'h5f : _GEN_4477; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4479 = 8'h7f == io_state_in_5 ? 8'h54 : _GEN_4478; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4480 = 8'h80 == io_state_in_5 ? 8'hf7 : _GEN_4479; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4481 = 8'h81 == io_state_in_5 ? 8'hfc : _GEN_4480; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4482 = 8'h82 == io_state_in_5 ? 8'he1 : _GEN_4481; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4483 = 8'h83 == io_state_in_5 ? 8'hea : _GEN_4482; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4484 = 8'h84 == io_state_in_5 ? 8'hdb : _GEN_4483; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4485 = 8'h85 == io_state_in_5 ? 8'hd0 : _GEN_4484; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4486 = 8'h86 == io_state_in_5 ? 8'hcd : _GEN_4485; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4487 = 8'h87 == io_state_in_5 ? 8'hc6 : _GEN_4486; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4488 = 8'h88 == io_state_in_5 ? 8'haf : _GEN_4487; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4489 = 8'h89 == io_state_in_5 ? 8'ha4 : _GEN_4488; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4490 = 8'h8a == io_state_in_5 ? 8'hb9 : _GEN_4489; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4491 = 8'h8b == io_state_in_5 ? 8'hb2 : _GEN_4490; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4492 = 8'h8c == io_state_in_5 ? 8'h83 : _GEN_4491; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4493 = 8'h8d == io_state_in_5 ? 8'h88 : _GEN_4492; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4494 = 8'h8e == io_state_in_5 ? 8'h95 : _GEN_4493; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4495 = 8'h8f == io_state_in_5 ? 8'h9e : _GEN_4494; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4496 = 8'h90 == io_state_in_5 ? 8'h47 : _GEN_4495; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4497 = 8'h91 == io_state_in_5 ? 8'h4c : _GEN_4496; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4498 = 8'h92 == io_state_in_5 ? 8'h51 : _GEN_4497; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4499 = 8'h93 == io_state_in_5 ? 8'h5a : _GEN_4498; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4500 = 8'h94 == io_state_in_5 ? 8'h6b : _GEN_4499; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4501 = 8'h95 == io_state_in_5 ? 8'h60 : _GEN_4500; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4502 = 8'h96 == io_state_in_5 ? 8'h7d : _GEN_4501; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4503 = 8'h97 == io_state_in_5 ? 8'h76 : _GEN_4502; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4504 = 8'h98 == io_state_in_5 ? 8'h1f : _GEN_4503; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4505 = 8'h99 == io_state_in_5 ? 8'h14 : _GEN_4504; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4506 = 8'h9a == io_state_in_5 ? 8'h9 : _GEN_4505; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4507 = 8'h9b == io_state_in_5 ? 8'h2 : _GEN_4506; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4508 = 8'h9c == io_state_in_5 ? 8'h33 : _GEN_4507; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4509 = 8'h9d == io_state_in_5 ? 8'h38 : _GEN_4508; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4510 = 8'h9e == io_state_in_5 ? 8'h25 : _GEN_4509; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4511 = 8'h9f == io_state_in_5 ? 8'h2e : _GEN_4510; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4512 = 8'ha0 == io_state_in_5 ? 8'h8c : _GEN_4511; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4513 = 8'ha1 == io_state_in_5 ? 8'h87 : _GEN_4512; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4514 = 8'ha2 == io_state_in_5 ? 8'h9a : _GEN_4513; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4515 = 8'ha3 == io_state_in_5 ? 8'h91 : _GEN_4514; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4516 = 8'ha4 == io_state_in_5 ? 8'ha0 : _GEN_4515; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4517 = 8'ha5 == io_state_in_5 ? 8'hab : _GEN_4516; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4518 = 8'ha6 == io_state_in_5 ? 8'hb6 : _GEN_4517; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4519 = 8'ha7 == io_state_in_5 ? 8'hbd : _GEN_4518; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4520 = 8'ha8 == io_state_in_5 ? 8'hd4 : _GEN_4519; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4521 = 8'ha9 == io_state_in_5 ? 8'hdf : _GEN_4520; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4522 = 8'haa == io_state_in_5 ? 8'hc2 : _GEN_4521; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4523 = 8'hab == io_state_in_5 ? 8'hc9 : _GEN_4522; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4524 = 8'hac == io_state_in_5 ? 8'hf8 : _GEN_4523; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4525 = 8'had == io_state_in_5 ? 8'hf3 : _GEN_4524; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4526 = 8'hae == io_state_in_5 ? 8'hee : _GEN_4525; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4527 = 8'haf == io_state_in_5 ? 8'he5 : _GEN_4526; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4528 = 8'hb0 == io_state_in_5 ? 8'h3c : _GEN_4527; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4529 = 8'hb1 == io_state_in_5 ? 8'h37 : _GEN_4528; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4530 = 8'hb2 == io_state_in_5 ? 8'h2a : _GEN_4529; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4531 = 8'hb3 == io_state_in_5 ? 8'h21 : _GEN_4530; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4532 = 8'hb4 == io_state_in_5 ? 8'h10 : _GEN_4531; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4533 = 8'hb5 == io_state_in_5 ? 8'h1b : _GEN_4532; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4534 = 8'hb6 == io_state_in_5 ? 8'h6 : _GEN_4533; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4535 = 8'hb7 == io_state_in_5 ? 8'hd : _GEN_4534; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4536 = 8'hb8 == io_state_in_5 ? 8'h64 : _GEN_4535; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4537 = 8'hb9 == io_state_in_5 ? 8'h6f : _GEN_4536; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4538 = 8'hba == io_state_in_5 ? 8'h72 : _GEN_4537; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4539 = 8'hbb == io_state_in_5 ? 8'h79 : _GEN_4538; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4540 = 8'hbc == io_state_in_5 ? 8'h48 : _GEN_4539; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4541 = 8'hbd == io_state_in_5 ? 8'h43 : _GEN_4540; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4542 = 8'hbe == io_state_in_5 ? 8'h5e : _GEN_4541; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4543 = 8'hbf == io_state_in_5 ? 8'h55 : _GEN_4542; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4544 = 8'hc0 == io_state_in_5 ? 8'h1 : _GEN_4543; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4545 = 8'hc1 == io_state_in_5 ? 8'ha : _GEN_4544; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4546 = 8'hc2 == io_state_in_5 ? 8'h17 : _GEN_4545; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4547 = 8'hc3 == io_state_in_5 ? 8'h1c : _GEN_4546; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4548 = 8'hc4 == io_state_in_5 ? 8'h2d : _GEN_4547; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4549 = 8'hc5 == io_state_in_5 ? 8'h26 : _GEN_4548; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4550 = 8'hc6 == io_state_in_5 ? 8'h3b : _GEN_4549; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4551 = 8'hc7 == io_state_in_5 ? 8'h30 : _GEN_4550; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4552 = 8'hc8 == io_state_in_5 ? 8'h59 : _GEN_4551; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4553 = 8'hc9 == io_state_in_5 ? 8'h52 : _GEN_4552; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4554 = 8'hca == io_state_in_5 ? 8'h4f : _GEN_4553; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4555 = 8'hcb == io_state_in_5 ? 8'h44 : _GEN_4554; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4556 = 8'hcc == io_state_in_5 ? 8'h75 : _GEN_4555; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4557 = 8'hcd == io_state_in_5 ? 8'h7e : _GEN_4556; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4558 = 8'hce == io_state_in_5 ? 8'h63 : _GEN_4557; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4559 = 8'hcf == io_state_in_5 ? 8'h68 : _GEN_4558; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4560 = 8'hd0 == io_state_in_5 ? 8'hb1 : _GEN_4559; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4561 = 8'hd1 == io_state_in_5 ? 8'hba : _GEN_4560; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4562 = 8'hd2 == io_state_in_5 ? 8'ha7 : _GEN_4561; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4563 = 8'hd3 == io_state_in_5 ? 8'hac : _GEN_4562; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4564 = 8'hd4 == io_state_in_5 ? 8'h9d : _GEN_4563; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4565 = 8'hd5 == io_state_in_5 ? 8'h96 : _GEN_4564; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4566 = 8'hd6 == io_state_in_5 ? 8'h8b : _GEN_4565; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4567 = 8'hd7 == io_state_in_5 ? 8'h80 : _GEN_4566; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4568 = 8'hd8 == io_state_in_5 ? 8'he9 : _GEN_4567; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4569 = 8'hd9 == io_state_in_5 ? 8'he2 : _GEN_4568; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4570 = 8'hda == io_state_in_5 ? 8'hff : _GEN_4569; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4571 = 8'hdb == io_state_in_5 ? 8'hf4 : _GEN_4570; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4572 = 8'hdc == io_state_in_5 ? 8'hc5 : _GEN_4571; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4573 = 8'hdd == io_state_in_5 ? 8'hce : _GEN_4572; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4574 = 8'hde == io_state_in_5 ? 8'hd3 : _GEN_4573; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4575 = 8'hdf == io_state_in_5 ? 8'hd8 : _GEN_4574; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4576 = 8'he0 == io_state_in_5 ? 8'h7a : _GEN_4575; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4577 = 8'he1 == io_state_in_5 ? 8'h71 : _GEN_4576; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4578 = 8'he2 == io_state_in_5 ? 8'h6c : _GEN_4577; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4579 = 8'he3 == io_state_in_5 ? 8'h67 : _GEN_4578; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4580 = 8'he4 == io_state_in_5 ? 8'h56 : _GEN_4579; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4581 = 8'he5 == io_state_in_5 ? 8'h5d : _GEN_4580; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4582 = 8'he6 == io_state_in_5 ? 8'h40 : _GEN_4581; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4583 = 8'he7 == io_state_in_5 ? 8'h4b : _GEN_4582; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4584 = 8'he8 == io_state_in_5 ? 8'h22 : _GEN_4583; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4585 = 8'he9 == io_state_in_5 ? 8'h29 : _GEN_4584; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4586 = 8'hea == io_state_in_5 ? 8'h34 : _GEN_4585; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4587 = 8'heb == io_state_in_5 ? 8'h3f : _GEN_4586; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4588 = 8'hec == io_state_in_5 ? 8'he : _GEN_4587; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4589 = 8'hed == io_state_in_5 ? 8'h5 : _GEN_4588; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4590 = 8'hee == io_state_in_5 ? 8'h18 : _GEN_4589; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4591 = 8'hef == io_state_in_5 ? 8'h13 : _GEN_4590; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4592 = 8'hf0 == io_state_in_5 ? 8'hca : _GEN_4591; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4593 = 8'hf1 == io_state_in_5 ? 8'hc1 : _GEN_4592; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4594 = 8'hf2 == io_state_in_5 ? 8'hdc : _GEN_4593; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4595 = 8'hf3 == io_state_in_5 ? 8'hd7 : _GEN_4594; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4596 = 8'hf4 == io_state_in_5 ? 8'he6 : _GEN_4595; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4597 = 8'hf5 == io_state_in_5 ? 8'hed : _GEN_4596; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4598 = 8'hf6 == io_state_in_5 ? 8'hf0 : _GEN_4597; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4599 = 8'hf7 == io_state_in_5 ? 8'hfb : _GEN_4598; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4600 = 8'hf8 == io_state_in_5 ? 8'h92 : _GEN_4599; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4601 = 8'hf9 == io_state_in_5 ? 8'h99 : _GEN_4600; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4602 = 8'hfa == io_state_in_5 ? 8'h84 : _GEN_4601; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4603 = 8'hfb == io_state_in_5 ? 8'h8f : _GEN_4602; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4604 = 8'hfc == io_state_in_5 ? 8'hbe : _GEN_4603; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4605 = 8'hfd == io_state_in_5 ? 8'hb5 : _GEN_4604; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4606 = 8'hfe == io_state_in_5 ? 8'ha8 : _GEN_4605; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _GEN_4607 = 8'hff == io_state_in_5 ? 8'ha3 : _GEN_4606; // @[InvMixColumns.scala 131:{41,41}]
  wire [7:0] _tmp_state_4_T = _GEN_4351 ^ _GEN_4607; // @[InvMixColumns.scala 131:41]
  wire [7:0] _GEN_4609 = 8'h1 == io_state_in_6 ? 8'hd : 8'h0; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4610 = 8'h2 == io_state_in_6 ? 8'h1a : _GEN_4609; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4611 = 8'h3 == io_state_in_6 ? 8'h17 : _GEN_4610; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4612 = 8'h4 == io_state_in_6 ? 8'h34 : _GEN_4611; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4613 = 8'h5 == io_state_in_6 ? 8'h39 : _GEN_4612; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4614 = 8'h6 == io_state_in_6 ? 8'h2e : _GEN_4613; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4615 = 8'h7 == io_state_in_6 ? 8'h23 : _GEN_4614; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4616 = 8'h8 == io_state_in_6 ? 8'h68 : _GEN_4615; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4617 = 8'h9 == io_state_in_6 ? 8'h65 : _GEN_4616; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4618 = 8'ha == io_state_in_6 ? 8'h72 : _GEN_4617; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4619 = 8'hb == io_state_in_6 ? 8'h7f : _GEN_4618; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4620 = 8'hc == io_state_in_6 ? 8'h5c : _GEN_4619; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4621 = 8'hd == io_state_in_6 ? 8'h51 : _GEN_4620; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4622 = 8'he == io_state_in_6 ? 8'h46 : _GEN_4621; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4623 = 8'hf == io_state_in_6 ? 8'h4b : _GEN_4622; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4624 = 8'h10 == io_state_in_6 ? 8'hd0 : _GEN_4623; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4625 = 8'h11 == io_state_in_6 ? 8'hdd : _GEN_4624; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4626 = 8'h12 == io_state_in_6 ? 8'hca : _GEN_4625; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4627 = 8'h13 == io_state_in_6 ? 8'hc7 : _GEN_4626; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4628 = 8'h14 == io_state_in_6 ? 8'he4 : _GEN_4627; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4629 = 8'h15 == io_state_in_6 ? 8'he9 : _GEN_4628; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4630 = 8'h16 == io_state_in_6 ? 8'hfe : _GEN_4629; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4631 = 8'h17 == io_state_in_6 ? 8'hf3 : _GEN_4630; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4632 = 8'h18 == io_state_in_6 ? 8'hb8 : _GEN_4631; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4633 = 8'h19 == io_state_in_6 ? 8'hb5 : _GEN_4632; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4634 = 8'h1a == io_state_in_6 ? 8'ha2 : _GEN_4633; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4635 = 8'h1b == io_state_in_6 ? 8'haf : _GEN_4634; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4636 = 8'h1c == io_state_in_6 ? 8'h8c : _GEN_4635; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4637 = 8'h1d == io_state_in_6 ? 8'h81 : _GEN_4636; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4638 = 8'h1e == io_state_in_6 ? 8'h96 : _GEN_4637; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4639 = 8'h1f == io_state_in_6 ? 8'h9b : _GEN_4638; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4640 = 8'h20 == io_state_in_6 ? 8'hbb : _GEN_4639; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4641 = 8'h21 == io_state_in_6 ? 8'hb6 : _GEN_4640; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4642 = 8'h22 == io_state_in_6 ? 8'ha1 : _GEN_4641; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4643 = 8'h23 == io_state_in_6 ? 8'hac : _GEN_4642; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4644 = 8'h24 == io_state_in_6 ? 8'h8f : _GEN_4643; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4645 = 8'h25 == io_state_in_6 ? 8'h82 : _GEN_4644; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4646 = 8'h26 == io_state_in_6 ? 8'h95 : _GEN_4645; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4647 = 8'h27 == io_state_in_6 ? 8'h98 : _GEN_4646; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4648 = 8'h28 == io_state_in_6 ? 8'hd3 : _GEN_4647; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4649 = 8'h29 == io_state_in_6 ? 8'hde : _GEN_4648; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4650 = 8'h2a == io_state_in_6 ? 8'hc9 : _GEN_4649; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4651 = 8'h2b == io_state_in_6 ? 8'hc4 : _GEN_4650; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4652 = 8'h2c == io_state_in_6 ? 8'he7 : _GEN_4651; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4653 = 8'h2d == io_state_in_6 ? 8'hea : _GEN_4652; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4654 = 8'h2e == io_state_in_6 ? 8'hfd : _GEN_4653; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4655 = 8'h2f == io_state_in_6 ? 8'hf0 : _GEN_4654; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4656 = 8'h30 == io_state_in_6 ? 8'h6b : _GEN_4655; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4657 = 8'h31 == io_state_in_6 ? 8'h66 : _GEN_4656; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4658 = 8'h32 == io_state_in_6 ? 8'h71 : _GEN_4657; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4659 = 8'h33 == io_state_in_6 ? 8'h7c : _GEN_4658; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4660 = 8'h34 == io_state_in_6 ? 8'h5f : _GEN_4659; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4661 = 8'h35 == io_state_in_6 ? 8'h52 : _GEN_4660; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4662 = 8'h36 == io_state_in_6 ? 8'h45 : _GEN_4661; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4663 = 8'h37 == io_state_in_6 ? 8'h48 : _GEN_4662; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4664 = 8'h38 == io_state_in_6 ? 8'h3 : _GEN_4663; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4665 = 8'h39 == io_state_in_6 ? 8'he : _GEN_4664; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4666 = 8'h3a == io_state_in_6 ? 8'h19 : _GEN_4665; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4667 = 8'h3b == io_state_in_6 ? 8'h14 : _GEN_4666; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4668 = 8'h3c == io_state_in_6 ? 8'h37 : _GEN_4667; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4669 = 8'h3d == io_state_in_6 ? 8'h3a : _GEN_4668; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4670 = 8'h3e == io_state_in_6 ? 8'h2d : _GEN_4669; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4671 = 8'h3f == io_state_in_6 ? 8'h20 : _GEN_4670; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4672 = 8'h40 == io_state_in_6 ? 8'h6d : _GEN_4671; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4673 = 8'h41 == io_state_in_6 ? 8'h60 : _GEN_4672; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4674 = 8'h42 == io_state_in_6 ? 8'h77 : _GEN_4673; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4675 = 8'h43 == io_state_in_6 ? 8'h7a : _GEN_4674; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4676 = 8'h44 == io_state_in_6 ? 8'h59 : _GEN_4675; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4677 = 8'h45 == io_state_in_6 ? 8'h54 : _GEN_4676; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4678 = 8'h46 == io_state_in_6 ? 8'h43 : _GEN_4677; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4679 = 8'h47 == io_state_in_6 ? 8'h4e : _GEN_4678; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4680 = 8'h48 == io_state_in_6 ? 8'h5 : _GEN_4679; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4681 = 8'h49 == io_state_in_6 ? 8'h8 : _GEN_4680; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4682 = 8'h4a == io_state_in_6 ? 8'h1f : _GEN_4681; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4683 = 8'h4b == io_state_in_6 ? 8'h12 : _GEN_4682; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4684 = 8'h4c == io_state_in_6 ? 8'h31 : _GEN_4683; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4685 = 8'h4d == io_state_in_6 ? 8'h3c : _GEN_4684; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4686 = 8'h4e == io_state_in_6 ? 8'h2b : _GEN_4685; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4687 = 8'h4f == io_state_in_6 ? 8'h26 : _GEN_4686; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4688 = 8'h50 == io_state_in_6 ? 8'hbd : _GEN_4687; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4689 = 8'h51 == io_state_in_6 ? 8'hb0 : _GEN_4688; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4690 = 8'h52 == io_state_in_6 ? 8'ha7 : _GEN_4689; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4691 = 8'h53 == io_state_in_6 ? 8'haa : _GEN_4690; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4692 = 8'h54 == io_state_in_6 ? 8'h89 : _GEN_4691; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4693 = 8'h55 == io_state_in_6 ? 8'h84 : _GEN_4692; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4694 = 8'h56 == io_state_in_6 ? 8'h93 : _GEN_4693; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4695 = 8'h57 == io_state_in_6 ? 8'h9e : _GEN_4694; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4696 = 8'h58 == io_state_in_6 ? 8'hd5 : _GEN_4695; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4697 = 8'h59 == io_state_in_6 ? 8'hd8 : _GEN_4696; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4698 = 8'h5a == io_state_in_6 ? 8'hcf : _GEN_4697; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4699 = 8'h5b == io_state_in_6 ? 8'hc2 : _GEN_4698; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4700 = 8'h5c == io_state_in_6 ? 8'he1 : _GEN_4699; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4701 = 8'h5d == io_state_in_6 ? 8'hec : _GEN_4700; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4702 = 8'h5e == io_state_in_6 ? 8'hfb : _GEN_4701; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4703 = 8'h5f == io_state_in_6 ? 8'hf6 : _GEN_4702; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4704 = 8'h60 == io_state_in_6 ? 8'hd6 : _GEN_4703; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4705 = 8'h61 == io_state_in_6 ? 8'hdb : _GEN_4704; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4706 = 8'h62 == io_state_in_6 ? 8'hcc : _GEN_4705; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4707 = 8'h63 == io_state_in_6 ? 8'hc1 : _GEN_4706; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4708 = 8'h64 == io_state_in_6 ? 8'he2 : _GEN_4707; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4709 = 8'h65 == io_state_in_6 ? 8'hef : _GEN_4708; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4710 = 8'h66 == io_state_in_6 ? 8'hf8 : _GEN_4709; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4711 = 8'h67 == io_state_in_6 ? 8'hf5 : _GEN_4710; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4712 = 8'h68 == io_state_in_6 ? 8'hbe : _GEN_4711; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4713 = 8'h69 == io_state_in_6 ? 8'hb3 : _GEN_4712; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4714 = 8'h6a == io_state_in_6 ? 8'ha4 : _GEN_4713; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4715 = 8'h6b == io_state_in_6 ? 8'ha9 : _GEN_4714; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4716 = 8'h6c == io_state_in_6 ? 8'h8a : _GEN_4715; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4717 = 8'h6d == io_state_in_6 ? 8'h87 : _GEN_4716; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4718 = 8'h6e == io_state_in_6 ? 8'h90 : _GEN_4717; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4719 = 8'h6f == io_state_in_6 ? 8'h9d : _GEN_4718; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4720 = 8'h70 == io_state_in_6 ? 8'h6 : _GEN_4719; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4721 = 8'h71 == io_state_in_6 ? 8'hb : _GEN_4720; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4722 = 8'h72 == io_state_in_6 ? 8'h1c : _GEN_4721; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4723 = 8'h73 == io_state_in_6 ? 8'h11 : _GEN_4722; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4724 = 8'h74 == io_state_in_6 ? 8'h32 : _GEN_4723; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4725 = 8'h75 == io_state_in_6 ? 8'h3f : _GEN_4724; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4726 = 8'h76 == io_state_in_6 ? 8'h28 : _GEN_4725; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4727 = 8'h77 == io_state_in_6 ? 8'h25 : _GEN_4726; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4728 = 8'h78 == io_state_in_6 ? 8'h6e : _GEN_4727; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4729 = 8'h79 == io_state_in_6 ? 8'h63 : _GEN_4728; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4730 = 8'h7a == io_state_in_6 ? 8'h74 : _GEN_4729; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4731 = 8'h7b == io_state_in_6 ? 8'h79 : _GEN_4730; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4732 = 8'h7c == io_state_in_6 ? 8'h5a : _GEN_4731; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4733 = 8'h7d == io_state_in_6 ? 8'h57 : _GEN_4732; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4734 = 8'h7e == io_state_in_6 ? 8'h40 : _GEN_4733; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4735 = 8'h7f == io_state_in_6 ? 8'h4d : _GEN_4734; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4736 = 8'h80 == io_state_in_6 ? 8'hda : _GEN_4735; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4737 = 8'h81 == io_state_in_6 ? 8'hd7 : _GEN_4736; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4738 = 8'h82 == io_state_in_6 ? 8'hc0 : _GEN_4737; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4739 = 8'h83 == io_state_in_6 ? 8'hcd : _GEN_4738; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4740 = 8'h84 == io_state_in_6 ? 8'hee : _GEN_4739; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4741 = 8'h85 == io_state_in_6 ? 8'he3 : _GEN_4740; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4742 = 8'h86 == io_state_in_6 ? 8'hf4 : _GEN_4741; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4743 = 8'h87 == io_state_in_6 ? 8'hf9 : _GEN_4742; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4744 = 8'h88 == io_state_in_6 ? 8'hb2 : _GEN_4743; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4745 = 8'h89 == io_state_in_6 ? 8'hbf : _GEN_4744; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4746 = 8'h8a == io_state_in_6 ? 8'ha8 : _GEN_4745; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4747 = 8'h8b == io_state_in_6 ? 8'ha5 : _GEN_4746; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4748 = 8'h8c == io_state_in_6 ? 8'h86 : _GEN_4747; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4749 = 8'h8d == io_state_in_6 ? 8'h8b : _GEN_4748; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4750 = 8'h8e == io_state_in_6 ? 8'h9c : _GEN_4749; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4751 = 8'h8f == io_state_in_6 ? 8'h91 : _GEN_4750; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4752 = 8'h90 == io_state_in_6 ? 8'ha : _GEN_4751; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4753 = 8'h91 == io_state_in_6 ? 8'h7 : _GEN_4752; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4754 = 8'h92 == io_state_in_6 ? 8'h10 : _GEN_4753; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4755 = 8'h93 == io_state_in_6 ? 8'h1d : _GEN_4754; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4756 = 8'h94 == io_state_in_6 ? 8'h3e : _GEN_4755; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4757 = 8'h95 == io_state_in_6 ? 8'h33 : _GEN_4756; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4758 = 8'h96 == io_state_in_6 ? 8'h24 : _GEN_4757; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4759 = 8'h97 == io_state_in_6 ? 8'h29 : _GEN_4758; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4760 = 8'h98 == io_state_in_6 ? 8'h62 : _GEN_4759; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4761 = 8'h99 == io_state_in_6 ? 8'h6f : _GEN_4760; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4762 = 8'h9a == io_state_in_6 ? 8'h78 : _GEN_4761; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4763 = 8'h9b == io_state_in_6 ? 8'h75 : _GEN_4762; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4764 = 8'h9c == io_state_in_6 ? 8'h56 : _GEN_4763; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4765 = 8'h9d == io_state_in_6 ? 8'h5b : _GEN_4764; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4766 = 8'h9e == io_state_in_6 ? 8'h4c : _GEN_4765; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4767 = 8'h9f == io_state_in_6 ? 8'h41 : _GEN_4766; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4768 = 8'ha0 == io_state_in_6 ? 8'h61 : _GEN_4767; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4769 = 8'ha1 == io_state_in_6 ? 8'h6c : _GEN_4768; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4770 = 8'ha2 == io_state_in_6 ? 8'h7b : _GEN_4769; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4771 = 8'ha3 == io_state_in_6 ? 8'h76 : _GEN_4770; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4772 = 8'ha4 == io_state_in_6 ? 8'h55 : _GEN_4771; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4773 = 8'ha5 == io_state_in_6 ? 8'h58 : _GEN_4772; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4774 = 8'ha6 == io_state_in_6 ? 8'h4f : _GEN_4773; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4775 = 8'ha7 == io_state_in_6 ? 8'h42 : _GEN_4774; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4776 = 8'ha8 == io_state_in_6 ? 8'h9 : _GEN_4775; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4777 = 8'ha9 == io_state_in_6 ? 8'h4 : _GEN_4776; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4778 = 8'haa == io_state_in_6 ? 8'h13 : _GEN_4777; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4779 = 8'hab == io_state_in_6 ? 8'h1e : _GEN_4778; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4780 = 8'hac == io_state_in_6 ? 8'h3d : _GEN_4779; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4781 = 8'had == io_state_in_6 ? 8'h30 : _GEN_4780; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4782 = 8'hae == io_state_in_6 ? 8'h27 : _GEN_4781; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4783 = 8'haf == io_state_in_6 ? 8'h2a : _GEN_4782; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4784 = 8'hb0 == io_state_in_6 ? 8'hb1 : _GEN_4783; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4785 = 8'hb1 == io_state_in_6 ? 8'hbc : _GEN_4784; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4786 = 8'hb2 == io_state_in_6 ? 8'hab : _GEN_4785; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4787 = 8'hb3 == io_state_in_6 ? 8'ha6 : _GEN_4786; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4788 = 8'hb4 == io_state_in_6 ? 8'h85 : _GEN_4787; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4789 = 8'hb5 == io_state_in_6 ? 8'h88 : _GEN_4788; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4790 = 8'hb6 == io_state_in_6 ? 8'h9f : _GEN_4789; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4791 = 8'hb7 == io_state_in_6 ? 8'h92 : _GEN_4790; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4792 = 8'hb8 == io_state_in_6 ? 8'hd9 : _GEN_4791; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4793 = 8'hb9 == io_state_in_6 ? 8'hd4 : _GEN_4792; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4794 = 8'hba == io_state_in_6 ? 8'hc3 : _GEN_4793; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4795 = 8'hbb == io_state_in_6 ? 8'hce : _GEN_4794; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4796 = 8'hbc == io_state_in_6 ? 8'hed : _GEN_4795; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4797 = 8'hbd == io_state_in_6 ? 8'he0 : _GEN_4796; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4798 = 8'hbe == io_state_in_6 ? 8'hf7 : _GEN_4797; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4799 = 8'hbf == io_state_in_6 ? 8'hfa : _GEN_4798; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4800 = 8'hc0 == io_state_in_6 ? 8'hb7 : _GEN_4799; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4801 = 8'hc1 == io_state_in_6 ? 8'hba : _GEN_4800; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4802 = 8'hc2 == io_state_in_6 ? 8'had : _GEN_4801; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4803 = 8'hc3 == io_state_in_6 ? 8'ha0 : _GEN_4802; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4804 = 8'hc4 == io_state_in_6 ? 8'h83 : _GEN_4803; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4805 = 8'hc5 == io_state_in_6 ? 8'h8e : _GEN_4804; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4806 = 8'hc6 == io_state_in_6 ? 8'h99 : _GEN_4805; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4807 = 8'hc7 == io_state_in_6 ? 8'h94 : _GEN_4806; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4808 = 8'hc8 == io_state_in_6 ? 8'hdf : _GEN_4807; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4809 = 8'hc9 == io_state_in_6 ? 8'hd2 : _GEN_4808; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4810 = 8'hca == io_state_in_6 ? 8'hc5 : _GEN_4809; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4811 = 8'hcb == io_state_in_6 ? 8'hc8 : _GEN_4810; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4812 = 8'hcc == io_state_in_6 ? 8'heb : _GEN_4811; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4813 = 8'hcd == io_state_in_6 ? 8'he6 : _GEN_4812; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4814 = 8'hce == io_state_in_6 ? 8'hf1 : _GEN_4813; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4815 = 8'hcf == io_state_in_6 ? 8'hfc : _GEN_4814; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4816 = 8'hd0 == io_state_in_6 ? 8'h67 : _GEN_4815; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4817 = 8'hd1 == io_state_in_6 ? 8'h6a : _GEN_4816; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4818 = 8'hd2 == io_state_in_6 ? 8'h7d : _GEN_4817; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4819 = 8'hd3 == io_state_in_6 ? 8'h70 : _GEN_4818; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4820 = 8'hd4 == io_state_in_6 ? 8'h53 : _GEN_4819; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4821 = 8'hd5 == io_state_in_6 ? 8'h5e : _GEN_4820; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4822 = 8'hd6 == io_state_in_6 ? 8'h49 : _GEN_4821; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4823 = 8'hd7 == io_state_in_6 ? 8'h44 : _GEN_4822; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4824 = 8'hd8 == io_state_in_6 ? 8'hf : _GEN_4823; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4825 = 8'hd9 == io_state_in_6 ? 8'h2 : _GEN_4824; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4826 = 8'hda == io_state_in_6 ? 8'h15 : _GEN_4825; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4827 = 8'hdb == io_state_in_6 ? 8'h18 : _GEN_4826; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4828 = 8'hdc == io_state_in_6 ? 8'h3b : _GEN_4827; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4829 = 8'hdd == io_state_in_6 ? 8'h36 : _GEN_4828; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4830 = 8'hde == io_state_in_6 ? 8'h21 : _GEN_4829; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4831 = 8'hdf == io_state_in_6 ? 8'h2c : _GEN_4830; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4832 = 8'he0 == io_state_in_6 ? 8'hc : _GEN_4831; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4833 = 8'he1 == io_state_in_6 ? 8'h1 : _GEN_4832; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4834 = 8'he2 == io_state_in_6 ? 8'h16 : _GEN_4833; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4835 = 8'he3 == io_state_in_6 ? 8'h1b : _GEN_4834; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4836 = 8'he4 == io_state_in_6 ? 8'h38 : _GEN_4835; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4837 = 8'he5 == io_state_in_6 ? 8'h35 : _GEN_4836; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4838 = 8'he6 == io_state_in_6 ? 8'h22 : _GEN_4837; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4839 = 8'he7 == io_state_in_6 ? 8'h2f : _GEN_4838; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4840 = 8'he8 == io_state_in_6 ? 8'h64 : _GEN_4839; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4841 = 8'he9 == io_state_in_6 ? 8'h69 : _GEN_4840; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4842 = 8'hea == io_state_in_6 ? 8'h7e : _GEN_4841; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4843 = 8'heb == io_state_in_6 ? 8'h73 : _GEN_4842; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4844 = 8'hec == io_state_in_6 ? 8'h50 : _GEN_4843; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4845 = 8'hed == io_state_in_6 ? 8'h5d : _GEN_4844; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4846 = 8'hee == io_state_in_6 ? 8'h4a : _GEN_4845; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4847 = 8'hef == io_state_in_6 ? 8'h47 : _GEN_4846; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4848 = 8'hf0 == io_state_in_6 ? 8'hdc : _GEN_4847; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4849 = 8'hf1 == io_state_in_6 ? 8'hd1 : _GEN_4848; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4850 = 8'hf2 == io_state_in_6 ? 8'hc6 : _GEN_4849; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4851 = 8'hf3 == io_state_in_6 ? 8'hcb : _GEN_4850; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4852 = 8'hf4 == io_state_in_6 ? 8'he8 : _GEN_4851; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4853 = 8'hf5 == io_state_in_6 ? 8'he5 : _GEN_4852; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4854 = 8'hf6 == io_state_in_6 ? 8'hf2 : _GEN_4853; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4855 = 8'hf7 == io_state_in_6 ? 8'hff : _GEN_4854; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4856 = 8'hf8 == io_state_in_6 ? 8'hb4 : _GEN_4855; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4857 = 8'hf9 == io_state_in_6 ? 8'hb9 : _GEN_4856; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4858 = 8'hfa == io_state_in_6 ? 8'hae : _GEN_4857; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4859 = 8'hfb == io_state_in_6 ? 8'ha3 : _GEN_4858; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4860 = 8'hfc == io_state_in_6 ? 8'h80 : _GEN_4859; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4861 = 8'hfd == io_state_in_6 ? 8'h8d : _GEN_4860; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4862 = 8'hfe == io_state_in_6 ? 8'h9a : _GEN_4861; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _GEN_4863 = 8'hff == io_state_in_6 ? 8'h97 : _GEN_4862; // @[InvMixColumns.scala 131:{65,65}]
  wire [7:0] _tmp_state_4_T_1 = _tmp_state_4_T ^ _GEN_4863; // @[InvMixColumns.scala 131:65]
  wire [7:0] _GEN_4865 = 8'h1 == io_state_in_7 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4866 = 8'h2 == io_state_in_7 ? 8'h12 : _GEN_4865; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4867 = 8'h3 == io_state_in_7 ? 8'h1b : _GEN_4866; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4868 = 8'h4 == io_state_in_7 ? 8'h24 : _GEN_4867; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4869 = 8'h5 == io_state_in_7 ? 8'h2d : _GEN_4868; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4870 = 8'h6 == io_state_in_7 ? 8'h36 : _GEN_4869; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4871 = 8'h7 == io_state_in_7 ? 8'h3f : _GEN_4870; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4872 = 8'h8 == io_state_in_7 ? 8'h48 : _GEN_4871; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4873 = 8'h9 == io_state_in_7 ? 8'h41 : _GEN_4872; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4874 = 8'ha == io_state_in_7 ? 8'h5a : _GEN_4873; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4875 = 8'hb == io_state_in_7 ? 8'h53 : _GEN_4874; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4876 = 8'hc == io_state_in_7 ? 8'h6c : _GEN_4875; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4877 = 8'hd == io_state_in_7 ? 8'h65 : _GEN_4876; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4878 = 8'he == io_state_in_7 ? 8'h7e : _GEN_4877; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4879 = 8'hf == io_state_in_7 ? 8'h77 : _GEN_4878; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4880 = 8'h10 == io_state_in_7 ? 8'h90 : _GEN_4879; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4881 = 8'h11 == io_state_in_7 ? 8'h99 : _GEN_4880; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4882 = 8'h12 == io_state_in_7 ? 8'h82 : _GEN_4881; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4883 = 8'h13 == io_state_in_7 ? 8'h8b : _GEN_4882; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4884 = 8'h14 == io_state_in_7 ? 8'hb4 : _GEN_4883; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4885 = 8'h15 == io_state_in_7 ? 8'hbd : _GEN_4884; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4886 = 8'h16 == io_state_in_7 ? 8'ha6 : _GEN_4885; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4887 = 8'h17 == io_state_in_7 ? 8'haf : _GEN_4886; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4888 = 8'h18 == io_state_in_7 ? 8'hd8 : _GEN_4887; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4889 = 8'h19 == io_state_in_7 ? 8'hd1 : _GEN_4888; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4890 = 8'h1a == io_state_in_7 ? 8'hca : _GEN_4889; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4891 = 8'h1b == io_state_in_7 ? 8'hc3 : _GEN_4890; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4892 = 8'h1c == io_state_in_7 ? 8'hfc : _GEN_4891; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4893 = 8'h1d == io_state_in_7 ? 8'hf5 : _GEN_4892; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4894 = 8'h1e == io_state_in_7 ? 8'hee : _GEN_4893; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4895 = 8'h1f == io_state_in_7 ? 8'he7 : _GEN_4894; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4896 = 8'h20 == io_state_in_7 ? 8'h3b : _GEN_4895; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4897 = 8'h21 == io_state_in_7 ? 8'h32 : _GEN_4896; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4898 = 8'h22 == io_state_in_7 ? 8'h29 : _GEN_4897; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4899 = 8'h23 == io_state_in_7 ? 8'h20 : _GEN_4898; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4900 = 8'h24 == io_state_in_7 ? 8'h1f : _GEN_4899; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4901 = 8'h25 == io_state_in_7 ? 8'h16 : _GEN_4900; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4902 = 8'h26 == io_state_in_7 ? 8'hd : _GEN_4901; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4903 = 8'h27 == io_state_in_7 ? 8'h4 : _GEN_4902; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4904 = 8'h28 == io_state_in_7 ? 8'h73 : _GEN_4903; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4905 = 8'h29 == io_state_in_7 ? 8'h7a : _GEN_4904; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4906 = 8'h2a == io_state_in_7 ? 8'h61 : _GEN_4905; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4907 = 8'h2b == io_state_in_7 ? 8'h68 : _GEN_4906; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4908 = 8'h2c == io_state_in_7 ? 8'h57 : _GEN_4907; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4909 = 8'h2d == io_state_in_7 ? 8'h5e : _GEN_4908; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4910 = 8'h2e == io_state_in_7 ? 8'h45 : _GEN_4909; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4911 = 8'h2f == io_state_in_7 ? 8'h4c : _GEN_4910; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4912 = 8'h30 == io_state_in_7 ? 8'hab : _GEN_4911; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4913 = 8'h31 == io_state_in_7 ? 8'ha2 : _GEN_4912; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4914 = 8'h32 == io_state_in_7 ? 8'hb9 : _GEN_4913; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4915 = 8'h33 == io_state_in_7 ? 8'hb0 : _GEN_4914; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4916 = 8'h34 == io_state_in_7 ? 8'h8f : _GEN_4915; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4917 = 8'h35 == io_state_in_7 ? 8'h86 : _GEN_4916; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4918 = 8'h36 == io_state_in_7 ? 8'h9d : _GEN_4917; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4919 = 8'h37 == io_state_in_7 ? 8'h94 : _GEN_4918; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4920 = 8'h38 == io_state_in_7 ? 8'he3 : _GEN_4919; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4921 = 8'h39 == io_state_in_7 ? 8'hea : _GEN_4920; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4922 = 8'h3a == io_state_in_7 ? 8'hf1 : _GEN_4921; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4923 = 8'h3b == io_state_in_7 ? 8'hf8 : _GEN_4922; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4924 = 8'h3c == io_state_in_7 ? 8'hc7 : _GEN_4923; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4925 = 8'h3d == io_state_in_7 ? 8'hce : _GEN_4924; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4926 = 8'h3e == io_state_in_7 ? 8'hd5 : _GEN_4925; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4927 = 8'h3f == io_state_in_7 ? 8'hdc : _GEN_4926; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4928 = 8'h40 == io_state_in_7 ? 8'h76 : _GEN_4927; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4929 = 8'h41 == io_state_in_7 ? 8'h7f : _GEN_4928; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4930 = 8'h42 == io_state_in_7 ? 8'h64 : _GEN_4929; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4931 = 8'h43 == io_state_in_7 ? 8'h6d : _GEN_4930; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4932 = 8'h44 == io_state_in_7 ? 8'h52 : _GEN_4931; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4933 = 8'h45 == io_state_in_7 ? 8'h5b : _GEN_4932; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4934 = 8'h46 == io_state_in_7 ? 8'h40 : _GEN_4933; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4935 = 8'h47 == io_state_in_7 ? 8'h49 : _GEN_4934; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4936 = 8'h48 == io_state_in_7 ? 8'h3e : _GEN_4935; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4937 = 8'h49 == io_state_in_7 ? 8'h37 : _GEN_4936; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4938 = 8'h4a == io_state_in_7 ? 8'h2c : _GEN_4937; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4939 = 8'h4b == io_state_in_7 ? 8'h25 : _GEN_4938; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4940 = 8'h4c == io_state_in_7 ? 8'h1a : _GEN_4939; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4941 = 8'h4d == io_state_in_7 ? 8'h13 : _GEN_4940; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4942 = 8'h4e == io_state_in_7 ? 8'h8 : _GEN_4941; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4943 = 8'h4f == io_state_in_7 ? 8'h1 : _GEN_4942; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4944 = 8'h50 == io_state_in_7 ? 8'he6 : _GEN_4943; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4945 = 8'h51 == io_state_in_7 ? 8'hef : _GEN_4944; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4946 = 8'h52 == io_state_in_7 ? 8'hf4 : _GEN_4945; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4947 = 8'h53 == io_state_in_7 ? 8'hfd : _GEN_4946; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4948 = 8'h54 == io_state_in_7 ? 8'hc2 : _GEN_4947; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4949 = 8'h55 == io_state_in_7 ? 8'hcb : _GEN_4948; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4950 = 8'h56 == io_state_in_7 ? 8'hd0 : _GEN_4949; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4951 = 8'h57 == io_state_in_7 ? 8'hd9 : _GEN_4950; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4952 = 8'h58 == io_state_in_7 ? 8'hae : _GEN_4951; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4953 = 8'h59 == io_state_in_7 ? 8'ha7 : _GEN_4952; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4954 = 8'h5a == io_state_in_7 ? 8'hbc : _GEN_4953; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4955 = 8'h5b == io_state_in_7 ? 8'hb5 : _GEN_4954; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4956 = 8'h5c == io_state_in_7 ? 8'h8a : _GEN_4955; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4957 = 8'h5d == io_state_in_7 ? 8'h83 : _GEN_4956; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4958 = 8'h5e == io_state_in_7 ? 8'h98 : _GEN_4957; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4959 = 8'h5f == io_state_in_7 ? 8'h91 : _GEN_4958; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4960 = 8'h60 == io_state_in_7 ? 8'h4d : _GEN_4959; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4961 = 8'h61 == io_state_in_7 ? 8'h44 : _GEN_4960; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4962 = 8'h62 == io_state_in_7 ? 8'h5f : _GEN_4961; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4963 = 8'h63 == io_state_in_7 ? 8'h56 : _GEN_4962; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4964 = 8'h64 == io_state_in_7 ? 8'h69 : _GEN_4963; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4965 = 8'h65 == io_state_in_7 ? 8'h60 : _GEN_4964; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4966 = 8'h66 == io_state_in_7 ? 8'h7b : _GEN_4965; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4967 = 8'h67 == io_state_in_7 ? 8'h72 : _GEN_4966; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4968 = 8'h68 == io_state_in_7 ? 8'h5 : _GEN_4967; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4969 = 8'h69 == io_state_in_7 ? 8'hc : _GEN_4968; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4970 = 8'h6a == io_state_in_7 ? 8'h17 : _GEN_4969; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4971 = 8'h6b == io_state_in_7 ? 8'h1e : _GEN_4970; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4972 = 8'h6c == io_state_in_7 ? 8'h21 : _GEN_4971; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4973 = 8'h6d == io_state_in_7 ? 8'h28 : _GEN_4972; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4974 = 8'h6e == io_state_in_7 ? 8'h33 : _GEN_4973; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4975 = 8'h6f == io_state_in_7 ? 8'h3a : _GEN_4974; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4976 = 8'h70 == io_state_in_7 ? 8'hdd : _GEN_4975; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4977 = 8'h71 == io_state_in_7 ? 8'hd4 : _GEN_4976; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4978 = 8'h72 == io_state_in_7 ? 8'hcf : _GEN_4977; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4979 = 8'h73 == io_state_in_7 ? 8'hc6 : _GEN_4978; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4980 = 8'h74 == io_state_in_7 ? 8'hf9 : _GEN_4979; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4981 = 8'h75 == io_state_in_7 ? 8'hf0 : _GEN_4980; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4982 = 8'h76 == io_state_in_7 ? 8'heb : _GEN_4981; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4983 = 8'h77 == io_state_in_7 ? 8'he2 : _GEN_4982; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4984 = 8'h78 == io_state_in_7 ? 8'h95 : _GEN_4983; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4985 = 8'h79 == io_state_in_7 ? 8'h9c : _GEN_4984; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4986 = 8'h7a == io_state_in_7 ? 8'h87 : _GEN_4985; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4987 = 8'h7b == io_state_in_7 ? 8'h8e : _GEN_4986; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4988 = 8'h7c == io_state_in_7 ? 8'hb1 : _GEN_4987; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4989 = 8'h7d == io_state_in_7 ? 8'hb8 : _GEN_4988; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4990 = 8'h7e == io_state_in_7 ? 8'ha3 : _GEN_4989; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4991 = 8'h7f == io_state_in_7 ? 8'haa : _GEN_4990; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4992 = 8'h80 == io_state_in_7 ? 8'hec : _GEN_4991; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4993 = 8'h81 == io_state_in_7 ? 8'he5 : _GEN_4992; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4994 = 8'h82 == io_state_in_7 ? 8'hfe : _GEN_4993; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4995 = 8'h83 == io_state_in_7 ? 8'hf7 : _GEN_4994; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4996 = 8'h84 == io_state_in_7 ? 8'hc8 : _GEN_4995; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4997 = 8'h85 == io_state_in_7 ? 8'hc1 : _GEN_4996; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4998 = 8'h86 == io_state_in_7 ? 8'hda : _GEN_4997; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_4999 = 8'h87 == io_state_in_7 ? 8'hd3 : _GEN_4998; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5000 = 8'h88 == io_state_in_7 ? 8'ha4 : _GEN_4999; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5001 = 8'h89 == io_state_in_7 ? 8'had : _GEN_5000; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5002 = 8'h8a == io_state_in_7 ? 8'hb6 : _GEN_5001; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5003 = 8'h8b == io_state_in_7 ? 8'hbf : _GEN_5002; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5004 = 8'h8c == io_state_in_7 ? 8'h80 : _GEN_5003; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5005 = 8'h8d == io_state_in_7 ? 8'h89 : _GEN_5004; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5006 = 8'h8e == io_state_in_7 ? 8'h92 : _GEN_5005; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5007 = 8'h8f == io_state_in_7 ? 8'h9b : _GEN_5006; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5008 = 8'h90 == io_state_in_7 ? 8'h7c : _GEN_5007; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5009 = 8'h91 == io_state_in_7 ? 8'h75 : _GEN_5008; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5010 = 8'h92 == io_state_in_7 ? 8'h6e : _GEN_5009; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5011 = 8'h93 == io_state_in_7 ? 8'h67 : _GEN_5010; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5012 = 8'h94 == io_state_in_7 ? 8'h58 : _GEN_5011; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5013 = 8'h95 == io_state_in_7 ? 8'h51 : _GEN_5012; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5014 = 8'h96 == io_state_in_7 ? 8'h4a : _GEN_5013; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5015 = 8'h97 == io_state_in_7 ? 8'h43 : _GEN_5014; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5016 = 8'h98 == io_state_in_7 ? 8'h34 : _GEN_5015; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5017 = 8'h99 == io_state_in_7 ? 8'h3d : _GEN_5016; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5018 = 8'h9a == io_state_in_7 ? 8'h26 : _GEN_5017; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5019 = 8'h9b == io_state_in_7 ? 8'h2f : _GEN_5018; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5020 = 8'h9c == io_state_in_7 ? 8'h10 : _GEN_5019; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5021 = 8'h9d == io_state_in_7 ? 8'h19 : _GEN_5020; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5022 = 8'h9e == io_state_in_7 ? 8'h2 : _GEN_5021; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5023 = 8'h9f == io_state_in_7 ? 8'hb : _GEN_5022; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5024 = 8'ha0 == io_state_in_7 ? 8'hd7 : _GEN_5023; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5025 = 8'ha1 == io_state_in_7 ? 8'hde : _GEN_5024; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5026 = 8'ha2 == io_state_in_7 ? 8'hc5 : _GEN_5025; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5027 = 8'ha3 == io_state_in_7 ? 8'hcc : _GEN_5026; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5028 = 8'ha4 == io_state_in_7 ? 8'hf3 : _GEN_5027; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5029 = 8'ha5 == io_state_in_7 ? 8'hfa : _GEN_5028; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5030 = 8'ha6 == io_state_in_7 ? 8'he1 : _GEN_5029; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5031 = 8'ha7 == io_state_in_7 ? 8'he8 : _GEN_5030; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5032 = 8'ha8 == io_state_in_7 ? 8'h9f : _GEN_5031; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5033 = 8'ha9 == io_state_in_7 ? 8'h96 : _GEN_5032; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5034 = 8'haa == io_state_in_7 ? 8'h8d : _GEN_5033; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5035 = 8'hab == io_state_in_7 ? 8'h84 : _GEN_5034; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5036 = 8'hac == io_state_in_7 ? 8'hbb : _GEN_5035; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5037 = 8'had == io_state_in_7 ? 8'hb2 : _GEN_5036; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5038 = 8'hae == io_state_in_7 ? 8'ha9 : _GEN_5037; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5039 = 8'haf == io_state_in_7 ? 8'ha0 : _GEN_5038; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5040 = 8'hb0 == io_state_in_7 ? 8'h47 : _GEN_5039; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5041 = 8'hb1 == io_state_in_7 ? 8'h4e : _GEN_5040; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5042 = 8'hb2 == io_state_in_7 ? 8'h55 : _GEN_5041; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5043 = 8'hb3 == io_state_in_7 ? 8'h5c : _GEN_5042; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5044 = 8'hb4 == io_state_in_7 ? 8'h63 : _GEN_5043; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5045 = 8'hb5 == io_state_in_7 ? 8'h6a : _GEN_5044; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5046 = 8'hb6 == io_state_in_7 ? 8'h71 : _GEN_5045; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5047 = 8'hb7 == io_state_in_7 ? 8'h78 : _GEN_5046; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5048 = 8'hb8 == io_state_in_7 ? 8'hf : _GEN_5047; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5049 = 8'hb9 == io_state_in_7 ? 8'h6 : _GEN_5048; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5050 = 8'hba == io_state_in_7 ? 8'h1d : _GEN_5049; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5051 = 8'hbb == io_state_in_7 ? 8'h14 : _GEN_5050; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5052 = 8'hbc == io_state_in_7 ? 8'h2b : _GEN_5051; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5053 = 8'hbd == io_state_in_7 ? 8'h22 : _GEN_5052; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5054 = 8'hbe == io_state_in_7 ? 8'h39 : _GEN_5053; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5055 = 8'hbf == io_state_in_7 ? 8'h30 : _GEN_5054; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5056 = 8'hc0 == io_state_in_7 ? 8'h9a : _GEN_5055; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5057 = 8'hc1 == io_state_in_7 ? 8'h93 : _GEN_5056; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5058 = 8'hc2 == io_state_in_7 ? 8'h88 : _GEN_5057; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5059 = 8'hc3 == io_state_in_7 ? 8'h81 : _GEN_5058; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5060 = 8'hc4 == io_state_in_7 ? 8'hbe : _GEN_5059; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5061 = 8'hc5 == io_state_in_7 ? 8'hb7 : _GEN_5060; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5062 = 8'hc6 == io_state_in_7 ? 8'hac : _GEN_5061; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5063 = 8'hc7 == io_state_in_7 ? 8'ha5 : _GEN_5062; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5064 = 8'hc8 == io_state_in_7 ? 8'hd2 : _GEN_5063; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5065 = 8'hc9 == io_state_in_7 ? 8'hdb : _GEN_5064; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5066 = 8'hca == io_state_in_7 ? 8'hc0 : _GEN_5065; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5067 = 8'hcb == io_state_in_7 ? 8'hc9 : _GEN_5066; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5068 = 8'hcc == io_state_in_7 ? 8'hf6 : _GEN_5067; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5069 = 8'hcd == io_state_in_7 ? 8'hff : _GEN_5068; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5070 = 8'hce == io_state_in_7 ? 8'he4 : _GEN_5069; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5071 = 8'hcf == io_state_in_7 ? 8'hed : _GEN_5070; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5072 = 8'hd0 == io_state_in_7 ? 8'ha : _GEN_5071; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5073 = 8'hd1 == io_state_in_7 ? 8'h3 : _GEN_5072; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5074 = 8'hd2 == io_state_in_7 ? 8'h18 : _GEN_5073; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5075 = 8'hd3 == io_state_in_7 ? 8'h11 : _GEN_5074; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5076 = 8'hd4 == io_state_in_7 ? 8'h2e : _GEN_5075; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5077 = 8'hd5 == io_state_in_7 ? 8'h27 : _GEN_5076; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5078 = 8'hd6 == io_state_in_7 ? 8'h3c : _GEN_5077; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5079 = 8'hd7 == io_state_in_7 ? 8'h35 : _GEN_5078; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5080 = 8'hd8 == io_state_in_7 ? 8'h42 : _GEN_5079; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5081 = 8'hd9 == io_state_in_7 ? 8'h4b : _GEN_5080; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5082 = 8'hda == io_state_in_7 ? 8'h50 : _GEN_5081; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5083 = 8'hdb == io_state_in_7 ? 8'h59 : _GEN_5082; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5084 = 8'hdc == io_state_in_7 ? 8'h66 : _GEN_5083; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5085 = 8'hdd == io_state_in_7 ? 8'h6f : _GEN_5084; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5086 = 8'hde == io_state_in_7 ? 8'h74 : _GEN_5085; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5087 = 8'hdf == io_state_in_7 ? 8'h7d : _GEN_5086; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5088 = 8'he0 == io_state_in_7 ? 8'ha1 : _GEN_5087; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5089 = 8'he1 == io_state_in_7 ? 8'ha8 : _GEN_5088; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5090 = 8'he2 == io_state_in_7 ? 8'hb3 : _GEN_5089; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5091 = 8'he3 == io_state_in_7 ? 8'hba : _GEN_5090; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5092 = 8'he4 == io_state_in_7 ? 8'h85 : _GEN_5091; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5093 = 8'he5 == io_state_in_7 ? 8'h8c : _GEN_5092; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5094 = 8'he6 == io_state_in_7 ? 8'h97 : _GEN_5093; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5095 = 8'he7 == io_state_in_7 ? 8'h9e : _GEN_5094; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5096 = 8'he8 == io_state_in_7 ? 8'he9 : _GEN_5095; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5097 = 8'he9 == io_state_in_7 ? 8'he0 : _GEN_5096; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5098 = 8'hea == io_state_in_7 ? 8'hfb : _GEN_5097; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5099 = 8'heb == io_state_in_7 ? 8'hf2 : _GEN_5098; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5100 = 8'hec == io_state_in_7 ? 8'hcd : _GEN_5099; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5101 = 8'hed == io_state_in_7 ? 8'hc4 : _GEN_5100; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5102 = 8'hee == io_state_in_7 ? 8'hdf : _GEN_5101; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5103 = 8'hef == io_state_in_7 ? 8'hd6 : _GEN_5102; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5104 = 8'hf0 == io_state_in_7 ? 8'h31 : _GEN_5103; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5105 = 8'hf1 == io_state_in_7 ? 8'h38 : _GEN_5104; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5106 = 8'hf2 == io_state_in_7 ? 8'h23 : _GEN_5105; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5107 = 8'hf3 == io_state_in_7 ? 8'h2a : _GEN_5106; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5108 = 8'hf4 == io_state_in_7 ? 8'h15 : _GEN_5107; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5109 = 8'hf5 == io_state_in_7 ? 8'h1c : _GEN_5108; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5110 = 8'hf6 == io_state_in_7 ? 8'h7 : _GEN_5109; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5111 = 8'hf7 == io_state_in_7 ? 8'he : _GEN_5110; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5112 = 8'hf8 == io_state_in_7 ? 8'h79 : _GEN_5111; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5113 = 8'hf9 == io_state_in_7 ? 8'h70 : _GEN_5112; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5114 = 8'hfa == io_state_in_7 ? 8'h6b : _GEN_5113; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5115 = 8'hfb == io_state_in_7 ? 8'h62 : _GEN_5114; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5116 = 8'hfc == io_state_in_7 ? 8'h5d : _GEN_5115; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5117 = 8'hfd == io_state_in_7 ? 8'h54 : _GEN_5116; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5118 = 8'hfe == io_state_in_7 ? 8'h4f : _GEN_5117; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5119 = 8'hff == io_state_in_7 ? 8'h46 : _GEN_5118; // @[InvMixColumns.scala 131:{89,89}]
  wire [7:0] _GEN_5121 = 8'h1 == io_state_in_4 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5122 = 8'h2 == io_state_in_4 ? 8'h12 : _GEN_5121; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5123 = 8'h3 == io_state_in_4 ? 8'h1b : _GEN_5122; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5124 = 8'h4 == io_state_in_4 ? 8'h24 : _GEN_5123; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5125 = 8'h5 == io_state_in_4 ? 8'h2d : _GEN_5124; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5126 = 8'h6 == io_state_in_4 ? 8'h36 : _GEN_5125; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5127 = 8'h7 == io_state_in_4 ? 8'h3f : _GEN_5126; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5128 = 8'h8 == io_state_in_4 ? 8'h48 : _GEN_5127; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5129 = 8'h9 == io_state_in_4 ? 8'h41 : _GEN_5128; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5130 = 8'ha == io_state_in_4 ? 8'h5a : _GEN_5129; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5131 = 8'hb == io_state_in_4 ? 8'h53 : _GEN_5130; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5132 = 8'hc == io_state_in_4 ? 8'h6c : _GEN_5131; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5133 = 8'hd == io_state_in_4 ? 8'h65 : _GEN_5132; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5134 = 8'he == io_state_in_4 ? 8'h7e : _GEN_5133; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5135 = 8'hf == io_state_in_4 ? 8'h77 : _GEN_5134; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5136 = 8'h10 == io_state_in_4 ? 8'h90 : _GEN_5135; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5137 = 8'h11 == io_state_in_4 ? 8'h99 : _GEN_5136; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5138 = 8'h12 == io_state_in_4 ? 8'h82 : _GEN_5137; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5139 = 8'h13 == io_state_in_4 ? 8'h8b : _GEN_5138; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5140 = 8'h14 == io_state_in_4 ? 8'hb4 : _GEN_5139; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5141 = 8'h15 == io_state_in_4 ? 8'hbd : _GEN_5140; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5142 = 8'h16 == io_state_in_4 ? 8'ha6 : _GEN_5141; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5143 = 8'h17 == io_state_in_4 ? 8'haf : _GEN_5142; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5144 = 8'h18 == io_state_in_4 ? 8'hd8 : _GEN_5143; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5145 = 8'h19 == io_state_in_4 ? 8'hd1 : _GEN_5144; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5146 = 8'h1a == io_state_in_4 ? 8'hca : _GEN_5145; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5147 = 8'h1b == io_state_in_4 ? 8'hc3 : _GEN_5146; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5148 = 8'h1c == io_state_in_4 ? 8'hfc : _GEN_5147; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5149 = 8'h1d == io_state_in_4 ? 8'hf5 : _GEN_5148; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5150 = 8'h1e == io_state_in_4 ? 8'hee : _GEN_5149; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5151 = 8'h1f == io_state_in_4 ? 8'he7 : _GEN_5150; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5152 = 8'h20 == io_state_in_4 ? 8'h3b : _GEN_5151; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5153 = 8'h21 == io_state_in_4 ? 8'h32 : _GEN_5152; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5154 = 8'h22 == io_state_in_4 ? 8'h29 : _GEN_5153; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5155 = 8'h23 == io_state_in_4 ? 8'h20 : _GEN_5154; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5156 = 8'h24 == io_state_in_4 ? 8'h1f : _GEN_5155; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5157 = 8'h25 == io_state_in_4 ? 8'h16 : _GEN_5156; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5158 = 8'h26 == io_state_in_4 ? 8'hd : _GEN_5157; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5159 = 8'h27 == io_state_in_4 ? 8'h4 : _GEN_5158; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5160 = 8'h28 == io_state_in_4 ? 8'h73 : _GEN_5159; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5161 = 8'h29 == io_state_in_4 ? 8'h7a : _GEN_5160; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5162 = 8'h2a == io_state_in_4 ? 8'h61 : _GEN_5161; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5163 = 8'h2b == io_state_in_4 ? 8'h68 : _GEN_5162; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5164 = 8'h2c == io_state_in_4 ? 8'h57 : _GEN_5163; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5165 = 8'h2d == io_state_in_4 ? 8'h5e : _GEN_5164; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5166 = 8'h2e == io_state_in_4 ? 8'h45 : _GEN_5165; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5167 = 8'h2f == io_state_in_4 ? 8'h4c : _GEN_5166; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5168 = 8'h30 == io_state_in_4 ? 8'hab : _GEN_5167; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5169 = 8'h31 == io_state_in_4 ? 8'ha2 : _GEN_5168; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5170 = 8'h32 == io_state_in_4 ? 8'hb9 : _GEN_5169; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5171 = 8'h33 == io_state_in_4 ? 8'hb0 : _GEN_5170; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5172 = 8'h34 == io_state_in_4 ? 8'h8f : _GEN_5171; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5173 = 8'h35 == io_state_in_4 ? 8'h86 : _GEN_5172; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5174 = 8'h36 == io_state_in_4 ? 8'h9d : _GEN_5173; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5175 = 8'h37 == io_state_in_4 ? 8'h94 : _GEN_5174; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5176 = 8'h38 == io_state_in_4 ? 8'he3 : _GEN_5175; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5177 = 8'h39 == io_state_in_4 ? 8'hea : _GEN_5176; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5178 = 8'h3a == io_state_in_4 ? 8'hf1 : _GEN_5177; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5179 = 8'h3b == io_state_in_4 ? 8'hf8 : _GEN_5178; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5180 = 8'h3c == io_state_in_4 ? 8'hc7 : _GEN_5179; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5181 = 8'h3d == io_state_in_4 ? 8'hce : _GEN_5180; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5182 = 8'h3e == io_state_in_4 ? 8'hd5 : _GEN_5181; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5183 = 8'h3f == io_state_in_4 ? 8'hdc : _GEN_5182; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5184 = 8'h40 == io_state_in_4 ? 8'h76 : _GEN_5183; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5185 = 8'h41 == io_state_in_4 ? 8'h7f : _GEN_5184; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5186 = 8'h42 == io_state_in_4 ? 8'h64 : _GEN_5185; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5187 = 8'h43 == io_state_in_4 ? 8'h6d : _GEN_5186; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5188 = 8'h44 == io_state_in_4 ? 8'h52 : _GEN_5187; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5189 = 8'h45 == io_state_in_4 ? 8'h5b : _GEN_5188; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5190 = 8'h46 == io_state_in_4 ? 8'h40 : _GEN_5189; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5191 = 8'h47 == io_state_in_4 ? 8'h49 : _GEN_5190; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5192 = 8'h48 == io_state_in_4 ? 8'h3e : _GEN_5191; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5193 = 8'h49 == io_state_in_4 ? 8'h37 : _GEN_5192; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5194 = 8'h4a == io_state_in_4 ? 8'h2c : _GEN_5193; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5195 = 8'h4b == io_state_in_4 ? 8'h25 : _GEN_5194; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5196 = 8'h4c == io_state_in_4 ? 8'h1a : _GEN_5195; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5197 = 8'h4d == io_state_in_4 ? 8'h13 : _GEN_5196; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5198 = 8'h4e == io_state_in_4 ? 8'h8 : _GEN_5197; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5199 = 8'h4f == io_state_in_4 ? 8'h1 : _GEN_5198; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5200 = 8'h50 == io_state_in_4 ? 8'he6 : _GEN_5199; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5201 = 8'h51 == io_state_in_4 ? 8'hef : _GEN_5200; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5202 = 8'h52 == io_state_in_4 ? 8'hf4 : _GEN_5201; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5203 = 8'h53 == io_state_in_4 ? 8'hfd : _GEN_5202; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5204 = 8'h54 == io_state_in_4 ? 8'hc2 : _GEN_5203; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5205 = 8'h55 == io_state_in_4 ? 8'hcb : _GEN_5204; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5206 = 8'h56 == io_state_in_4 ? 8'hd0 : _GEN_5205; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5207 = 8'h57 == io_state_in_4 ? 8'hd9 : _GEN_5206; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5208 = 8'h58 == io_state_in_4 ? 8'hae : _GEN_5207; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5209 = 8'h59 == io_state_in_4 ? 8'ha7 : _GEN_5208; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5210 = 8'h5a == io_state_in_4 ? 8'hbc : _GEN_5209; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5211 = 8'h5b == io_state_in_4 ? 8'hb5 : _GEN_5210; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5212 = 8'h5c == io_state_in_4 ? 8'h8a : _GEN_5211; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5213 = 8'h5d == io_state_in_4 ? 8'h83 : _GEN_5212; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5214 = 8'h5e == io_state_in_4 ? 8'h98 : _GEN_5213; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5215 = 8'h5f == io_state_in_4 ? 8'h91 : _GEN_5214; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5216 = 8'h60 == io_state_in_4 ? 8'h4d : _GEN_5215; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5217 = 8'h61 == io_state_in_4 ? 8'h44 : _GEN_5216; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5218 = 8'h62 == io_state_in_4 ? 8'h5f : _GEN_5217; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5219 = 8'h63 == io_state_in_4 ? 8'h56 : _GEN_5218; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5220 = 8'h64 == io_state_in_4 ? 8'h69 : _GEN_5219; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5221 = 8'h65 == io_state_in_4 ? 8'h60 : _GEN_5220; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5222 = 8'h66 == io_state_in_4 ? 8'h7b : _GEN_5221; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5223 = 8'h67 == io_state_in_4 ? 8'h72 : _GEN_5222; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5224 = 8'h68 == io_state_in_4 ? 8'h5 : _GEN_5223; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5225 = 8'h69 == io_state_in_4 ? 8'hc : _GEN_5224; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5226 = 8'h6a == io_state_in_4 ? 8'h17 : _GEN_5225; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5227 = 8'h6b == io_state_in_4 ? 8'h1e : _GEN_5226; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5228 = 8'h6c == io_state_in_4 ? 8'h21 : _GEN_5227; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5229 = 8'h6d == io_state_in_4 ? 8'h28 : _GEN_5228; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5230 = 8'h6e == io_state_in_4 ? 8'h33 : _GEN_5229; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5231 = 8'h6f == io_state_in_4 ? 8'h3a : _GEN_5230; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5232 = 8'h70 == io_state_in_4 ? 8'hdd : _GEN_5231; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5233 = 8'h71 == io_state_in_4 ? 8'hd4 : _GEN_5232; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5234 = 8'h72 == io_state_in_4 ? 8'hcf : _GEN_5233; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5235 = 8'h73 == io_state_in_4 ? 8'hc6 : _GEN_5234; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5236 = 8'h74 == io_state_in_4 ? 8'hf9 : _GEN_5235; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5237 = 8'h75 == io_state_in_4 ? 8'hf0 : _GEN_5236; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5238 = 8'h76 == io_state_in_4 ? 8'heb : _GEN_5237; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5239 = 8'h77 == io_state_in_4 ? 8'he2 : _GEN_5238; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5240 = 8'h78 == io_state_in_4 ? 8'h95 : _GEN_5239; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5241 = 8'h79 == io_state_in_4 ? 8'h9c : _GEN_5240; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5242 = 8'h7a == io_state_in_4 ? 8'h87 : _GEN_5241; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5243 = 8'h7b == io_state_in_4 ? 8'h8e : _GEN_5242; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5244 = 8'h7c == io_state_in_4 ? 8'hb1 : _GEN_5243; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5245 = 8'h7d == io_state_in_4 ? 8'hb8 : _GEN_5244; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5246 = 8'h7e == io_state_in_4 ? 8'ha3 : _GEN_5245; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5247 = 8'h7f == io_state_in_4 ? 8'haa : _GEN_5246; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5248 = 8'h80 == io_state_in_4 ? 8'hec : _GEN_5247; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5249 = 8'h81 == io_state_in_4 ? 8'he5 : _GEN_5248; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5250 = 8'h82 == io_state_in_4 ? 8'hfe : _GEN_5249; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5251 = 8'h83 == io_state_in_4 ? 8'hf7 : _GEN_5250; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5252 = 8'h84 == io_state_in_4 ? 8'hc8 : _GEN_5251; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5253 = 8'h85 == io_state_in_4 ? 8'hc1 : _GEN_5252; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5254 = 8'h86 == io_state_in_4 ? 8'hda : _GEN_5253; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5255 = 8'h87 == io_state_in_4 ? 8'hd3 : _GEN_5254; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5256 = 8'h88 == io_state_in_4 ? 8'ha4 : _GEN_5255; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5257 = 8'h89 == io_state_in_4 ? 8'had : _GEN_5256; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5258 = 8'h8a == io_state_in_4 ? 8'hb6 : _GEN_5257; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5259 = 8'h8b == io_state_in_4 ? 8'hbf : _GEN_5258; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5260 = 8'h8c == io_state_in_4 ? 8'h80 : _GEN_5259; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5261 = 8'h8d == io_state_in_4 ? 8'h89 : _GEN_5260; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5262 = 8'h8e == io_state_in_4 ? 8'h92 : _GEN_5261; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5263 = 8'h8f == io_state_in_4 ? 8'h9b : _GEN_5262; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5264 = 8'h90 == io_state_in_4 ? 8'h7c : _GEN_5263; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5265 = 8'h91 == io_state_in_4 ? 8'h75 : _GEN_5264; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5266 = 8'h92 == io_state_in_4 ? 8'h6e : _GEN_5265; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5267 = 8'h93 == io_state_in_4 ? 8'h67 : _GEN_5266; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5268 = 8'h94 == io_state_in_4 ? 8'h58 : _GEN_5267; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5269 = 8'h95 == io_state_in_4 ? 8'h51 : _GEN_5268; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5270 = 8'h96 == io_state_in_4 ? 8'h4a : _GEN_5269; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5271 = 8'h97 == io_state_in_4 ? 8'h43 : _GEN_5270; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5272 = 8'h98 == io_state_in_4 ? 8'h34 : _GEN_5271; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5273 = 8'h99 == io_state_in_4 ? 8'h3d : _GEN_5272; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5274 = 8'h9a == io_state_in_4 ? 8'h26 : _GEN_5273; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5275 = 8'h9b == io_state_in_4 ? 8'h2f : _GEN_5274; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5276 = 8'h9c == io_state_in_4 ? 8'h10 : _GEN_5275; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5277 = 8'h9d == io_state_in_4 ? 8'h19 : _GEN_5276; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5278 = 8'h9e == io_state_in_4 ? 8'h2 : _GEN_5277; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5279 = 8'h9f == io_state_in_4 ? 8'hb : _GEN_5278; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5280 = 8'ha0 == io_state_in_4 ? 8'hd7 : _GEN_5279; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5281 = 8'ha1 == io_state_in_4 ? 8'hde : _GEN_5280; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5282 = 8'ha2 == io_state_in_4 ? 8'hc5 : _GEN_5281; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5283 = 8'ha3 == io_state_in_4 ? 8'hcc : _GEN_5282; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5284 = 8'ha4 == io_state_in_4 ? 8'hf3 : _GEN_5283; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5285 = 8'ha5 == io_state_in_4 ? 8'hfa : _GEN_5284; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5286 = 8'ha6 == io_state_in_4 ? 8'he1 : _GEN_5285; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5287 = 8'ha7 == io_state_in_4 ? 8'he8 : _GEN_5286; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5288 = 8'ha8 == io_state_in_4 ? 8'h9f : _GEN_5287; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5289 = 8'ha9 == io_state_in_4 ? 8'h96 : _GEN_5288; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5290 = 8'haa == io_state_in_4 ? 8'h8d : _GEN_5289; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5291 = 8'hab == io_state_in_4 ? 8'h84 : _GEN_5290; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5292 = 8'hac == io_state_in_4 ? 8'hbb : _GEN_5291; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5293 = 8'had == io_state_in_4 ? 8'hb2 : _GEN_5292; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5294 = 8'hae == io_state_in_4 ? 8'ha9 : _GEN_5293; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5295 = 8'haf == io_state_in_4 ? 8'ha0 : _GEN_5294; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5296 = 8'hb0 == io_state_in_4 ? 8'h47 : _GEN_5295; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5297 = 8'hb1 == io_state_in_4 ? 8'h4e : _GEN_5296; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5298 = 8'hb2 == io_state_in_4 ? 8'h55 : _GEN_5297; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5299 = 8'hb3 == io_state_in_4 ? 8'h5c : _GEN_5298; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5300 = 8'hb4 == io_state_in_4 ? 8'h63 : _GEN_5299; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5301 = 8'hb5 == io_state_in_4 ? 8'h6a : _GEN_5300; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5302 = 8'hb6 == io_state_in_4 ? 8'h71 : _GEN_5301; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5303 = 8'hb7 == io_state_in_4 ? 8'h78 : _GEN_5302; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5304 = 8'hb8 == io_state_in_4 ? 8'hf : _GEN_5303; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5305 = 8'hb9 == io_state_in_4 ? 8'h6 : _GEN_5304; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5306 = 8'hba == io_state_in_4 ? 8'h1d : _GEN_5305; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5307 = 8'hbb == io_state_in_4 ? 8'h14 : _GEN_5306; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5308 = 8'hbc == io_state_in_4 ? 8'h2b : _GEN_5307; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5309 = 8'hbd == io_state_in_4 ? 8'h22 : _GEN_5308; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5310 = 8'hbe == io_state_in_4 ? 8'h39 : _GEN_5309; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5311 = 8'hbf == io_state_in_4 ? 8'h30 : _GEN_5310; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5312 = 8'hc0 == io_state_in_4 ? 8'h9a : _GEN_5311; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5313 = 8'hc1 == io_state_in_4 ? 8'h93 : _GEN_5312; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5314 = 8'hc2 == io_state_in_4 ? 8'h88 : _GEN_5313; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5315 = 8'hc3 == io_state_in_4 ? 8'h81 : _GEN_5314; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5316 = 8'hc4 == io_state_in_4 ? 8'hbe : _GEN_5315; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5317 = 8'hc5 == io_state_in_4 ? 8'hb7 : _GEN_5316; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5318 = 8'hc6 == io_state_in_4 ? 8'hac : _GEN_5317; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5319 = 8'hc7 == io_state_in_4 ? 8'ha5 : _GEN_5318; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5320 = 8'hc8 == io_state_in_4 ? 8'hd2 : _GEN_5319; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5321 = 8'hc9 == io_state_in_4 ? 8'hdb : _GEN_5320; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5322 = 8'hca == io_state_in_4 ? 8'hc0 : _GEN_5321; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5323 = 8'hcb == io_state_in_4 ? 8'hc9 : _GEN_5322; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5324 = 8'hcc == io_state_in_4 ? 8'hf6 : _GEN_5323; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5325 = 8'hcd == io_state_in_4 ? 8'hff : _GEN_5324; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5326 = 8'hce == io_state_in_4 ? 8'he4 : _GEN_5325; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5327 = 8'hcf == io_state_in_4 ? 8'hed : _GEN_5326; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5328 = 8'hd0 == io_state_in_4 ? 8'ha : _GEN_5327; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5329 = 8'hd1 == io_state_in_4 ? 8'h3 : _GEN_5328; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5330 = 8'hd2 == io_state_in_4 ? 8'h18 : _GEN_5329; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5331 = 8'hd3 == io_state_in_4 ? 8'h11 : _GEN_5330; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5332 = 8'hd4 == io_state_in_4 ? 8'h2e : _GEN_5331; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5333 = 8'hd5 == io_state_in_4 ? 8'h27 : _GEN_5332; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5334 = 8'hd6 == io_state_in_4 ? 8'h3c : _GEN_5333; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5335 = 8'hd7 == io_state_in_4 ? 8'h35 : _GEN_5334; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5336 = 8'hd8 == io_state_in_4 ? 8'h42 : _GEN_5335; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5337 = 8'hd9 == io_state_in_4 ? 8'h4b : _GEN_5336; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5338 = 8'hda == io_state_in_4 ? 8'h50 : _GEN_5337; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5339 = 8'hdb == io_state_in_4 ? 8'h59 : _GEN_5338; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5340 = 8'hdc == io_state_in_4 ? 8'h66 : _GEN_5339; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5341 = 8'hdd == io_state_in_4 ? 8'h6f : _GEN_5340; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5342 = 8'hde == io_state_in_4 ? 8'h74 : _GEN_5341; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5343 = 8'hdf == io_state_in_4 ? 8'h7d : _GEN_5342; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5344 = 8'he0 == io_state_in_4 ? 8'ha1 : _GEN_5343; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5345 = 8'he1 == io_state_in_4 ? 8'ha8 : _GEN_5344; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5346 = 8'he2 == io_state_in_4 ? 8'hb3 : _GEN_5345; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5347 = 8'he3 == io_state_in_4 ? 8'hba : _GEN_5346; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5348 = 8'he4 == io_state_in_4 ? 8'h85 : _GEN_5347; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5349 = 8'he5 == io_state_in_4 ? 8'h8c : _GEN_5348; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5350 = 8'he6 == io_state_in_4 ? 8'h97 : _GEN_5349; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5351 = 8'he7 == io_state_in_4 ? 8'h9e : _GEN_5350; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5352 = 8'he8 == io_state_in_4 ? 8'he9 : _GEN_5351; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5353 = 8'he9 == io_state_in_4 ? 8'he0 : _GEN_5352; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5354 = 8'hea == io_state_in_4 ? 8'hfb : _GEN_5353; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5355 = 8'heb == io_state_in_4 ? 8'hf2 : _GEN_5354; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5356 = 8'hec == io_state_in_4 ? 8'hcd : _GEN_5355; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5357 = 8'hed == io_state_in_4 ? 8'hc4 : _GEN_5356; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5358 = 8'hee == io_state_in_4 ? 8'hdf : _GEN_5357; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5359 = 8'hef == io_state_in_4 ? 8'hd6 : _GEN_5358; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5360 = 8'hf0 == io_state_in_4 ? 8'h31 : _GEN_5359; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5361 = 8'hf1 == io_state_in_4 ? 8'h38 : _GEN_5360; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5362 = 8'hf2 == io_state_in_4 ? 8'h23 : _GEN_5361; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5363 = 8'hf3 == io_state_in_4 ? 8'h2a : _GEN_5362; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5364 = 8'hf4 == io_state_in_4 ? 8'h15 : _GEN_5363; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5365 = 8'hf5 == io_state_in_4 ? 8'h1c : _GEN_5364; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5366 = 8'hf6 == io_state_in_4 ? 8'h7 : _GEN_5365; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5367 = 8'hf7 == io_state_in_4 ? 8'he : _GEN_5366; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5368 = 8'hf8 == io_state_in_4 ? 8'h79 : _GEN_5367; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5369 = 8'hf9 == io_state_in_4 ? 8'h70 : _GEN_5368; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5370 = 8'hfa == io_state_in_4 ? 8'h6b : _GEN_5369; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5371 = 8'hfb == io_state_in_4 ? 8'h62 : _GEN_5370; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5372 = 8'hfc == io_state_in_4 ? 8'h5d : _GEN_5371; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5373 = 8'hfd == io_state_in_4 ? 8'h54 : _GEN_5372; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5374 = 8'hfe == io_state_in_4 ? 8'h4f : _GEN_5373; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5375 = 8'hff == io_state_in_4 ? 8'h46 : _GEN_5374; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5377 = 8'h1 == io_state_in_5 ? 8'he : 8'h0; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5378 = 8'h2 == io_state_in_5 ? 8'h1c : _GEN_5377; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5379 = 8'h3 == io_state_in_5 ? 8'h12 : _GEN_5378; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5380 = 8'h4 == io_state_in_5 ? 8'h38 : _GEN_5379; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5381 = 8'h5 == io_state_in_5 ? 8'h36 : _GEN_5380; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5382 = 8'h6 == io_state_in_5 ? 8'h24 : _GEN_5381; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5383 = 8'h7 == io_state_in_5 ? 8'h2a : _GEN_5382; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5384 = 8'h8 == io_state_in_5 ? 8'h70 : _GEN_5383; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5385 = 8'h9 == io_state_in_5 ? 8'h7e : _GEN_5384; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5386 = 8'ha == io_state_in_5 ? 8'h6c : _GEN_5385; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5387 = 8'hb == io_state_in_5 ? 8'h62 : _GEN_5386; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5388 = 8'hc == io_state_in_5 ? 8'h48 : _GEN_5387; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5389 = 8'hd == io_state_in_5 ? 8'h46 : _GEN_5388; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5390 = 8'he == io_state_in_5 ? 8'h54 : _GEN_5389; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5391 = 8'hf == io_state_in_5 ? 8'h5a : _GEN_5390; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5392 = 8'h10 == io_state_in_5 ? 8'he0 : _GEN_5391; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5393 = 8'h11 == io_state_in_5 ? 8'hee : _GEN_5392; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5394 = 8'h12 == io_state_in_5 ? 8'hfc : _GEN_5393; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5395 = 8'h13 == io_state_in_5 ? 8'hf2 : _GEN_5394; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5396 = 8'h14 == io_state_in_5 ? 8'hd8 : _GEN_5395; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5397 = 8'h15 == io_state_in_5 ? 8'hd6 : _GEN_5396; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5398 = 8'h16 == io_state_in_5 ? 8'hc4 : _GEN_5397; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5399 = 8'h17 == io_state_in_5 ? 8'hca : _GEN_5398; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5400 = 8'h18 == io_state_in_5 ? 8'h90 : _GEN_5399; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5401 = 8'h19 == io_state_in_5 ? 8'h9e : _GEN_5400; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5402 = 8'h1a == io_state_in_5 ? 8'h8c : _GEN_5401; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5403 = 8'h1b == io_state_in_5 ? 8'h82 : _GEN_5402; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5404 = 8'h1c == io_state_in_5 ? 8'ha8 : _GEN_5403; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5405 = 8'h1d == io_state_in_5 ? 8'ha6 : _GEN_5404; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5406 = 8'h1e == io_state_in_5 ? 8'hb4 : _GEN_5405; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5407 = 8'h1f == io_state_in_5 ? 8'hba : _GEN_5406; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5408 = 8'h20 == io_state_in_5 ? 8'hdb : _GEN_5407; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5409 = 8'h21 == io_state_in_5 ? 8'hd5 : _GEN_5408; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5410 = 8'h22 == io_state_in_5 ? 8'hc7 : _GEN_5409; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5411 = 8'h23 == io_state_in_5 ? 8'hc9 : _GEN_5410; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5412 = 8'h24 == io_state_in_5 ? 8'he3 : _GEN_5411; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5413 = 8'h25 == io_state_in_5 ? 8'hed : _GEN_5412; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5414 = 8'h26 == io_state_in_5 ? 8'hff : _GEN_5413; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5415 = 8'h27 == io_state_in_5 ? 8'hf1 : _GEN_5414; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5416 = 8'h28 == io_state_in_5 ? 8'hab : _GEN_5415; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5417 = 8'h29 == io_state_in_5 ? 8'ha5 : _GEN_5416; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5418 = 8'h2a == io_state_in_5 ? 8'hb7 : _GEN_5417; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5419 = 8'h2b == io_state_in_5 ? 8'hb9 : _GEN_5418; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5420 = 8'h2c == io_state_in_5 ? 8'h93 : _GEN_5419; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5421 = 8'h2d == io_state_in_5 ? 8'h9d : _GEN_5420; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5422 = 8'h2e == io_state_in_5 ? 8'h8f : _GEN_5421; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5423 = 8'h2f == io_state_in_5 ? 8'h81 : _GEN_5422; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5424 = 8'h30 == io_state_in_5 ? 8'h3b : _GEN_5423; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5425 = 8'h31 == io_state_in_5 ? 8'h35 : _GEN_5424; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5426 = 8'h32 == io_state_in_5 ? 8'h27 : _GEN_5425; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5427 = 8'h33 == io_state_in_5 ? 8'h29 : _GEN_5426; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5428 = 8'h34 == io_state_in_5 ? 8'h3 : _GEN_5427; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5429 = 8'h35 == io_state_in_5 ? 8'hd : _GEN_5428; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5430 = 8'h36 == io_state_in_5 ? 8'h1f : _GEN_5429; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5431 = 8'h37 == io_state_in_5 ? 8'h11 : _GEN_5430; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5432 = 8'h38 == io_state_in_5 ? 8'h4b : _GEN_5431; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5433 = 8'h39 == io_state_in_5 ? 8'h45 : _GEN_5432; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5434 = 8'h3a == io_state_in_5 ? 8'h57 : _GEN_5433; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5435 = 8'h3b == io_state_in_5 ? 8'h59 : _GEN_5434; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5436 = 8'h3c == io_state_in_5 ? 8'h73 : _GEN_5435; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5437 = 8'h3d == io_state_in_5 ? 8'h7d : _GEN_5436; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5438 = 8'h3e == io_state_in_5 ? 8'h6f : _GEN_5437; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5439 = 8'h3f == io_state_in_5 ? 8'h61 : _GEN_5438; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5440 = 8'h40 == io_state_in_5 ? 8'had : _GEN_5439; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5441 = 8'h41 == io_state_in_5 ? 8'ha3 : _GEN_5440; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5442 = 8'h42 == io_state_in_5 ? 8'hb1 : _GEN_5441; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5443 = 8'h43 == io_state_in_5 ? 8'hbf : _GEN_5442; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5444 = 8'h44 == io_state_in_5 ? 8'h95 : _GEN_5443; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5445 = 8'h45 == io_state_in_5 ? 8'h9b : _GEN_5444; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5446 = 8'h46 == io_state_in_5 ? 8'h89 : _GEN_5445; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5447 = 8'h47 == io_state_in_5 ? 8'h87 : _GEN_5446; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5448 = 8'h48 == io_state_in_5 ? 8'hdd : _GEN_5447; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5449 = 8'h49 == io_state_in_5 ? 8'hd3 : _GEN_5448; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5450 = 8'h4a == io_state_in_5 ? 8'hc1 : _GEN_5449; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5451 = 8'h4b == io_state_in_5 ? 8'hcf : _GEN_5450; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5452 = 8'h4c == io_state_in_5 ? 8'he5 : _GEN_5451; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5453 = 8'h4d == io_state_in_5 ? 8'heb : _GEN_5452; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5454 = 8'h4e == io_state_in_5 ? 8'hf9 : _GEN_5453; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5455 = 8'h4f == io_state_in_5 ? 8'hf7 : _GEN_5454; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5456 = 8'h50 == io_state_in_5 ? 8'h4d : _GEN_5455; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5457 = 8'h51 == io_state_in_5 ? 8'h43 : _GEN_5456; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5458 = 8'h52 == io_state_in_5 ? 8'h51 : _GEN_5457; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5459 = 8'h53 == io_state_in_5 ? 8'h5f : _GEN_5458; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5460 = 8'h54 == io_state_in_5 ? 8'h75 : _GEN_5459; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5461 = 8'h55 == io_state_in_5 ? 8'h7b : _GEN_5460; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5462 = 8'h56 == io_state_in_5 ? 8'h69 : _GEN_5461; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5463 = 8'h57 == io_state_in_5 ? 8'h67 : _GEN_5462; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5464 = 8'h58 == io_state_in_5 ? 8'h3d : _GEN_5463; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5465 = 8'h59 == io_state_in_5 ? 8'h33 : _GEN_5464; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5466 = 8'h5a == io_state_in_5 ? 8'h21 : _GEN_5465; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5467 = 8'h5b == io_state_in_5 ? 8'h2f : _GEN_5466; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5468 = 8'h5c == io_state_in_5 ? 8'h5 : _GEN_5467; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5469 = 8'h5d == io_state_in_5 ? 8'hb : _GEN_5468; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5470 = 8'h5e == io_state_in_5 ? 8'h19 : _GEN_5469; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5471 = 8'h5f == io_state_in_5 ? 8'h17 : _GEN_5470; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5472 = 8'h60 == io_state_in_5 ? 8'h76 : _GEN_5471; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5473 = 8'h61 == io_state_in_5 ? 8'h78 : _GEN_5472; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5474 = 8'h62 == io_state_in_5 ? 8'h6a : _GEN_5473; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5475 = 8'h63 == io_state_in_5 ? 8'h64 : _GEN_5474; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5476 = 8'h64 == io_state_in_5 ? 8'h4e : _GEN_5475; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5477 = 8'h65 == io_state_in_5 ? 8'h40 : _GEN_5476; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5478 = 8'h66 == io_state_in_5 ? 8'h52 : _GEN_5477; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5479 = 8'h67 == io_state_in_5 ? 8'h5c : _GEN_5478; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5480 = 8'h68 == io_state_in_5 ? 8'h6 : _GEN_5479; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5481 = 8'h69 == io_state_in_5 ? 8'h8 : _GEN_5480; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5482 = 8'h6a == io_state_in_5 ? 8'h1a : _GEN_5481; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5483 = 8'h6b == io_state_in_5 ? 8'h14 : _GEN_5482; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5484 = 8'h6c == io_state_in_5 ? 8'h3e : _GEN_5483; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5485 = 8'h6d == io_state_in_5 ? 8'h30 : _GEN_5484; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5486 = 8'h6e == io_state_in_5 ? 8'h22 : _GEN_5485; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5487 = 8'h6f == io_state_in_5 ? 8'h2c : _GEN_5486; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5488 = 8'h70 == io_state_in_5 ? 8'h96 : _GEN_5487; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5489 = 8'h71 == io_state_in_5 ? 8'h98 : _GEN_5488; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5490 = 8'h72 == io_state_in_5 ? 8'h8a : _GEN_5489; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5491 = 8'h73 == io_state_in_5 ? 8'h84 : _GEN_5490; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5492 = 8'h74 == io_state_in_5 ? 8'hae : _GEN_5491; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5493 = 8'h75 == io_state_in_5 ? 8'ha0 : _GEN_5492; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5494 = 8'h76 == io_state_in_5 ? 8'hb2 : _GEN_5493; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5495 = 8'h77 == io_state_in_5 ? 8'hbc : _GEN_5494; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5496 = 8'h78 == io_state_in_5 ? 8'he6 : _GEN_5495; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5497 = 8'h79 == io_state_in_5 ? 8'he8 : _GEN_5496; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5498 = 8'h7a == io_state_in_5 ? 8'hfa : _GEN_5497; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5499 = 8'h7b == io_state_in_5 ? 8'hf4 : _GEN_5498; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5500 = 8'h7c == io_state_in_5 ? 8'hde : _GEN_5499; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5501 = 8'h7d == io_state_in_5 ? 8'hd0 : _GEN_5500; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5502 = 8'h7e == io_state_in_5 ? 8'hc2 : _GEN_5501; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5503 = 8'h7f == io_state_in_5 ? 8'hcc : _GEN_5502; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5504 = 8'h80 == io_state_in_5 ? 8'h41 : _GEN_5503; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5505 = 8'h81 == io_state_in_5 ? 8'h4f : _GEN_5504; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5506 = 8'h82 == io_state_in_5 ? 8'h5d : _GEN_5505; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5507 = 8'h83 == io_state_in_5 ? 8'h53 : _GEN_5506; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5508 = 8'h84 == io_state_in_5 ? 8'h79 : _GEN_5507; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5509 = 8'h85 == io_state_in_5 ? 8'h77 : _GEN_5508; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5510 = 8'h86 == io_state_in_5 ? 8'h65 : _GEN_5509; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5511 = 8'h87 == io_state_in_5 ? 8'h6b : _GEN_5510; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5512 = 8'h88 == io_state_in_5 ? 8'h31 : _GEN_5511; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5513 = 8'h89 == io_state_in_5 ? 8'h3f : _GEN_5512; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5514 = 8'h8a == io_state_in_5 ? 8'h2d : _GEN_5513; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5515 = 8'h8b == io_state_in_5 ? 8'h23 : _GEN_5514; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5516 = 8'h8c == io_state_in_5 ? 8'h9 : _GEN_5515; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5517 = 8'h8d == io_state_in_5 ? 8'h7 : _GEN_5516; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5518 = 8'h8e == io_state_in_5 ? 8'h15 : _GEN_5517; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5519 = 8'h8f == io_state_in_5 ? 8'h1b : _GEN_5518; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5520 = 8'h90 == io_state_in_5 ? 8'ha1 : _GEN_5519; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5521 = 8'h91 == io_state_in_5 ? 8'haf : _GEN_5520; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5522 = 8'h92 == io_state_in_5 ? 8'hbd : _GEN_5521; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5523 = 8'h93 == io_state_in_5 ? 8'hb3 : _GEN_5522; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5524 = 8'h94 == io_state_in_5 ? 8'h99 : _GEN_5523; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5525 = 8'h95 == io_state_in_5 ? 8'h97 : _GEN_5524; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5526 = 8'h96 == io_state_in_5 ? 8'h85 : _GEN_5525; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5527 = 8'h97 == io_state_in_5 ? 8'h8b : _GEN_5526; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5528 = 8'h98 == io_state_in_5 ? 8'hd1 : _GEN_5527; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5529 = 8'h99 == io_state_in_5 ? 8'hdf : _GEN_5528; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5530 = 8'h9a == io_state_in_5 ? 8'hcd : _GEN_5529; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5531 = 8'h9b == io_state_in_5 ? 8'hc3 : _GEN_5530; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5532 = 8'h9c == io_state_in_5 ? 8'he9 : _GEN_5531; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5533 = 8'h9d == io_state_in_5 ? 8'he7 : _GEN_5532; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5534 = 8'h9e == io_state_in_5 ? 8'hf5 : _GEN_5533; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5535 = 8'h9f == io_state_in_5 ? 8'hfb : _GEN_5534; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5536 = 8'ha0 == io_state_in_5 ? 8'h9a : _GEN_5535; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5537 = 8'ha1 == io_state_in_5 ? 8'h94 : _GEN_5536; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5538 = 8'ha2 == io_state_in_5 ? 8'h86 : _GEN_5537; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5539 = 8'ha3 == io_state_in_5 ? 8'h88 : _GEN_5538; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5540 = 8'ha4 == io_state_in_5 ? 8'ha2 : _GEN_5539; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5541 = 8'ha5 == io_state_in_5 ? 8'hac : _GEN_5540; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5542 = 8'ha6 == io_state_in_5 ? 8'hbe : _GEN_5541; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5543 = 8'ha7 == io_state_in_5 ? 8'hb0 : _GEN_5542; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5544 = 8'ha8 == io_state_in_5 ? 8'hea : _GEN_5543; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5545 = 8'ha9 == io_state_in_5 ? 8'he4 : _GEN_5544; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5546 = 8'haa == io_state_in_5 ? 8'hf6 : _GEN_5545; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5547 = 8'hab == io_state_in_5 ? 8'hf8 : _GEN_5546; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5548 = 8'hac == io_state_in_5 ? 8'hd2 : _GEN_5547; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5549 = 8'had == io_state_in_5 ? 8'hdc : _GEN_5548; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5550 = 8'hae == io_state_in_5 ? 8'hce : _GEN_5549; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5551 = 8'haf == io_state_in_5 ? 8'hc0 : _GEN_5550; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5552 = 8'hb0 == io_state_in_5 ? 8'h7a : _GEN_5551; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5553 = 8'hb1 == io_state_in_5 ? 8'h74 : _GEN_5552; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5554 = 8'hb2 == io_state_in_5 ? 8'h66 : _GEN_5553; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5555 = 8'hb3 == io_state_in_5 ? 8'h68 : _GEN_5554; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5556 = 8'hb4 == io_state_in_5 ? 8'h42 : _GEN_5555; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5557 = 8'hb5 == io_state_in_5 ? 8'h4c : _GEN_5556; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5558 = 8'hb6 == io_state_in_5 ? 8'h5e : _GEN_5557; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5559 = 8'hb7 == io_state_in_5 ? 8'h50 : _GEN_5558; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5560 = 8'hb8 == io_state_in_5 ? 8'ha : _GEN_5559; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5561 = 8'hb9 == io_state_in_5 ? 8'h4 : _GEN_5560; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5562 = 8'hba == io_state_in_5 ? 8'h16 : _GEN_5561; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5563 = 8'hbb == io_state_in_5 ? 8'h18 : _GEN_5562; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5564 = 8'hbc == io_state_in_5 ? 8'h32 : _GEN_5563; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5565 = 8'hbd == io_state_in_5 ? 8'h3c : _GEN_5564; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5566 = 8'hbe == io_state_in_5 ? 8'h2e : _GEN_5565; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5567 = 8'hbf == io_state_in_5 ? 8'h20 : _GEN_5566; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5568 = 8'hc0 == io_state_in_5 ? 8'hec : _GEN_5567; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5569 = 8'hc1 == io_state_in_5 ? 8'he2 : _GEN_5568; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5570 = 8'hc2 == io_state_in_5 ? 8'hf0 : _GEN_5569; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5571 = 8'hc3 == io_state_in_5 ? 8'hfe : _GEN_5570; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5572 = 8'hc4 == io_state_in_5 ? 8'hd4 : _GEN_5571; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5573 = 8'hc5 == io_state_in_5 ? 8'hda : _GEN_5572; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5574 = 8'hc6 == io_state_in_5 ? 8'hc8 : _GEN_5573; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5575 = 8'hc7 == io_state_in_5 ? 8'hc6 : _GEN_5574; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5576 = 8'hc8 == io_state_in_5 ? 8'h9c : _GEN_5575; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5577 = 8'hc9 == io_state_in_5 ? 8'h92 : _GEN_5576; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5578 = 8'hca == io_state_in_5 ? 8'h80 : _GEN_5577; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5579 = 8'hcb == io_state_in_5 ? 8'h8e : _GEN_5578; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5580 = 8'hcc == io_state_in_5 ? 8'ha4 : _GEN_5579; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5581 = 8'hcd == io_state_in_5 ? 8'haa : _GEN_5580; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5582 = 8'hce == io_state_in_5 ? 8'hb8 : _GEN_5581; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5583 = 8'hcf == io_state_in_5 ? 8'hb6 : _GEN_5582; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5584 = 8'hd0 == io_state_in_5 ? 8'hc : _GEN_5583; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5585 = 8'hd1 == io_state_in_5 ? 8'h2 : _GEN_5584; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5586 = 8'hd2 == io_state_in_5 ? 8'h10 : _GEN_5585; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5587 = 8'hd3 == io_state_in_5 ? 8'h1e : _GEN_5586; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5588 = 8'hd4 == io_state_in_5 ? 8'h34 : _GEN_5587; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5589 = 8'hd5 == io_state_in_5 ? 8'h3a : _GEN_5588; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5590 = 8'hd6 == io_state_in_5 ? 8'h28 : _GEN_5589; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5591 = 8'hd7 == io_state_in_5 ? 8'h26 : _GEN_5590; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5592 = 8'hd8 == io_state_in_5 ? 8'h7c : _GEN_5591; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5593 = 8'hd9 == io_state_in_5 ? 8'h72 : _GEN_5592; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5594 = 8'hda == io_state_in_5 ? 8'h60 : _GEN_5593; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5595 = 8'hdb == io_state_in_5 ? 8'h6e : _GEN_5594; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5596 = 8'hdc == io_state_in_5 ? 8'h44 : _GEN_5595; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5597 = 8'hdd == io_state_in_5 ? 8'h4a : _GEN_5596; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5598 = 8'hde == io_state_in_5 ? 8'h58 : _GEN_5597; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5599 = 8'hdf == io_state_in_5 ? 8'h56 : _GEN_5598; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5600 = 8'he0 == io_state_in_5 ? 8'h37 : _GEN_5599; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5601 = 8'he1 == io_state_in_5 ? 8'h39 : _GEN_5600; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5602 = 8'he2 == io_state_in_5 ? 8'h2b : _GEN_5601; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5603 = 8'he3 == io_state_in_5 ? 8'h25 : _GEN_5602; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5604 = 8'he4 == io_state_in_5 ? 8'hf : _GEN_5603; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5605 = 8'he5 == io_state_in_5 ? 8'h1 : _GEN_5604; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5606 = 8'he6 == io_state_in_5 ? 8'h13 : _GEN_5605; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5607 = 8'he7 == io_state_in_5 ? 8'h1d : _GEN_5606; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5608 = 8'he8 == io_state_in_5 ? 8'h47 : _GEN_5607; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5609 = 8'he9 == io_state_in_5 ? 8'h49 : _GEN_5608; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5610 = 8'hea == io_state_in_5 ? 8'h5b : _GEN_5609; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5611 = 8'heb == io_state_in_5 ? 8'h55 : _GEN_5610; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5612 = 8'hec == io_state_in_5 ? 8'h7f : _GEN_5611; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5613 = 8'hed == io_state_in_5 ? 8'h71 : _GEN_5612; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5614 = 8'hee == io_state_in_5 ? 8'h63 : _GEN_5613; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5615 = 8'hef == io_state_in_5 ? 8'h6d : _GEN_5614; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5616 = 8'hf0 == io_state_in_5 ? 8'hd7 : _GEN_5615; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5617 = 8'hf1 == io_state_in_5 ? 8'hd9 : _GEN_5616; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5618 = 8'hf2 == io_state_in_5 ? 8'hcb : _GEN_5617; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5619 = 8'hf3 == io_state_in_5 ? 8'hc5 : _GEN_5618; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5620 = 8'hf4 == io_state_in_5 ? 8'hef : _GEN_5619; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5621 = 8'hf5 == io_state_in_5 ? 8'he1 : _GEN_5620; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5622 = 8'hf6 == io_state_in_5 ? 8'hf3 : _GEN_5621; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5623 = 8'hf7 == io_state_in_5 ? 8'hfd : _GEN_5622; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5624 = 8'hf8 == io_state_in_5 ? 8'ha7 : _GEN_5623; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5625 = 8'hf9 == io_state_in_5 ? 8'ha9 : _GEN_5624; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5626 = 8'hfa == io_state_in_5 ? 8'hbb : _GEN_5625; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5627 = 8'hfb == io_state_in_5 ? 8'hb5 : _GEN_5626; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5628 = 8'hfc == io_state_in_5 ? 8'h9f : _GEN_5627; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5629 = 8'hfd == io_state_in_5 ? 8'h91 : _GEN_5628; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5630 = 8'hfe == io_state_in_5 ? 8'h83 : _GEN_5629; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _GEN_5631 = 8'hff == io_state_in_5 ? 8'h8d : _GEN_5630; // @[InvMixColumns.scala 132:{41,41}]
  wire [7:0] _tmp_state_5_T = _GEN_5375 ^ _GEN_5631; // @[InvMixColumns.scala 132:41]
  wire [7:0] _GEN_5633 = 8'h1 == io_state_in_6 ? 8'hb : 8'h0; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5634 = 8'h2 == io_state_in_6 ? 8'h16 : _GEN_5633; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5635 = 8'h3 == io_state_in_6 ? 8'h1d : _GEN_5634; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5636 = 8'h4 == io_state_in_6 ? 8'h2c : _GEN_5635; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5637 = 8'h5 == io_state_in_6 ? 8'h27 : _GEN_5636; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5638 = 8'h6 == io_state_in_6 ? 8'h3a : _GEN_5637; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5639 = 8'h7 == io_state_in_6 ? 8'h31 : _GEN_5638; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5640 = 8'h8 == io_state_in_6 ? 8'h58 : _GEN_5639; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5641 = 8'h9 == io_state_in_6 ? 8'h53 : _GEN_5640; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5642 = 8'ha == io_state_in_6 ? 8'h4e : _GEN_5641; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5643 = 8'hb == io_state_in_6 ? 8'h45 : _GEN_5642; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5644 = 8'hc == io_state_in_6 ? 8'h74 : _GEN_5643; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5645 = 8'hd == io_state_in_6 ? 8'h7f : _GEN_5644; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5646 = 8'he == io_state_in_6 ? 8'h62 : _GEN_5645; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5647 = 8'hf == io_state_in_6 ? 8'h69 : _GEN_5646; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5648 = 8'h10 == io_state_in_6 ? 8'hb0 : _GEN_5647; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5649 = 8'h11 == io_state_in_6 ? 8'hbb : _GEN_5648; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5650 = 8'h12 == io_state_in_6 ? 8'ha6 : _GEN_5649; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5651 = 8'h13 == io_state_in_6 ? 8'had : _GEN_5650; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5652 = 8'h14 == io_state_in_6 ? 8'h9c : _GEN_5651; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5653 = 8'h15 == io_state_in_6 ? 8'h97 : _GEN_5652; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5654 = 8'h16 == io_state_in_6 ? 8'h8a : _GEN_5653; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5655 = 8'h17 == io_state_in_6 ? 8'h81 : _GEN_5654; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5656 = 8'h18 == io_state_in_6 ? 8'he8 : _GEN_5655; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5657 = 8'h19 == io_state_in_6 ? 8'he3 : _GEN_5656; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5658 = 8'h1a == io_state_in_6 ? 8'hfe : _GEN_5657; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5659 = 8'h1b == io_state_in_6 ? 8'hf5 : _GEN_5658; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5660 = 8'h1c == io_state_in_6 ? 8'hc4 : _GEN_5659; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5661 = 8'h1d == io_state_in_6 ? 8'hcf : _GEN_5660; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5662 = 8'h1e == io_state_in_6 ? 8'hd2 : _GEN_5661; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5663 = 8'h1f == io_state_in_6 ? 8'hd9 : _GEN_5662; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5664 = 8'h20 == io_state_in_6 ? 8'h7b : _GEN_5663; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5665 = 8'h21 == io_state_in_6 ? 8'h70 : _GEN_5664; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5666 = 8'h22 == io_state_in_6 ? 8'h6d : _GEN_5665; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5667 = 8'h23 == io_state_in_6 ? 8'h66 : _GEN_5666; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5668 = 8'h24 == io_state_in_6 ? 8'h57 : _GEN_5667; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5669 = 8'h25 == io_state_in_6 ? 8'h5c : _GEN_5668; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5670 = 8'h26 == io_state_in_6 ? 8'h41 : _GEN_5669; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5671 = 8'h27 == io_state_in_6 ? 8'h4a : _GEN_5670; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5672 = 8'h28 == io_state_in_6 ? 8'h23 : _GEN_5671; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5673 = 8'h29 == io_state_in_6 ? 8'h28 : _GEN_5672; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5674 = 8'h2a == io_state_in_6 ? 8'h35 : _GEN_5673; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5675 = 8'h2b == io_state_in_6 ? 8'h3e : _GEN_5674; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5676 = 8'h2c == io_state_in_6 ? 8'hf : _GEN_5675; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5677 = 8'h2d == io_state_in_6 ? 8'h4 : _GEN_5676; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5678 = 8'h2e == io_state_in_6 ? 8'h19 : _GEN_5677; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5679 = 8'h2f == io_state_in_6 ? 8'h12 : _GEN_5678; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5680 = 8'h30 == io_state_in_6 ? 8'hcb : _GEN_5679; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5681 = 8'h31 == io_state_in_6 ? 8'hc0 : _GEN_5680; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5682 = 8'h32 == io_state_in_6 ? 8'hdd : _GEN_5681; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5683 = 8'h33 == io_state_in_6 ? 8'hd6 : _GEN_5682; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5684 = 8'h34 == io_state_in_6 ? 8'he7 : _GEN_5683; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5685 = 8'h35 == io_state_in_6 ? 8'hec : _GEN_5684; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5686 = 8'h36 == io_state_in_6 ? 8'hf1 : _GEN_5685; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5687 = 8'h37 == io_state_in_6 ? 8'hfa : _GEN_5686; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5688 = 8'h38 == io_state_in_6 ? 8'h93 : _GEN_5687; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5689 = 8'h39 == io_state_in_6 ? 8'h98 : _GEN_5688; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5690 = 8'h3a == io_state_in_6 ? 8'h85 : _GEN_5689; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5691 = 8'h3b == io_state_in_6 ? 8'h8e : _GEN_5690; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5692 = 8'h3c == io_state_in_6 ? 8'hbf : _GEN_5691; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5693 = 8'h3d == io_state_in_6 ? 8'hb4 : _GEN_5692; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5694 = 8'h3e == io_state_in_6 ? 8'ha9 : _GEN_5693; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5695 = 8'h3f == io_state_in_6 ? 8'ha2 : _GEN_5694; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5696 = 8'h40 == io_state_in_6 ? 8'hf6 : _GEN_5695; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5697 = 8'h41 == io_state_in_6 ? 8'hfd : _GEN_5696; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5698 = 8'h42 == io_state_in_6 ? 8'he0 : _GEN_5697; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5699 = 8'h43 == io_state_in_6 ? 8'heb : _GEN_5698; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5700 = 8'h44 == io_state_in_6 ? 8'hda : _GEN_5699; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5701 = 8'h45 == io_state_in_6 ? 8'hd1 : _GEN_5700; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5702 = 8'h46 == io_state_in_6 ? 8'hcc : _GEN_5701; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5703 = 8'h47 == io_state_in_6 ? 8'hc7 : _GEN_5702; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5704 = 8'h48 == io_state_in_6 ? 8'hae : _GEN_5703; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5705 = 8'h49 == io_state_in_6 ? 8'ha5 : _GEN_5704; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5706 = 8'h4a == io_state_in_6 ? 8'hb8 : _GEN_5705; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5707 = 8'h4b == io_state_in_6 ? 8'hb3 : _GEN_5706; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5708 = 8'h4c == io_state_in_6 ? 8'h82 : _GEN_5707; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5709 = 8'h4d == io_state_in_6 ? 8'h89 : _GEN_5708; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5710 = 8'h4e == io_state_in_6 ? 8'h94 : _GEN_5709; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5711 = 8'h4f == io_state_in_6 ? 8'h9f : _GEN_5710; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5712 = 8'h50 == io_state_in_6 ? 8'h46 : _GEN_5711; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5713 = 8'h51 == io_state_in_6 ? 8'h4d : _GEN_5712; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5714 = 8'h52 == io_state_in_6 ? 8'h50 : _GEN_5713; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5715 = 8'h53 == io_state_in_6 ? 8'h5b : _GEN_5714; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5716 = 8'h54 == io_state_in_6 ? 8'h6a : _GEN_5715; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5717 = 8'h55 == io_state_in_6 ? 8'h61 : _GEN_5716; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5718 = 8'h56 == io_state_in_6 ? 8'h7c : _GEN_5717; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5719 = 8'h57 == io_state_in_6 ? 8'h77 : _GEN_5718; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5720 = 8'h58 == io_state_in_6 ? 8'h1e : _GEN_5719; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5721 = 8'h59 == io_state_in_6 ? 8'h15 : _GEN_5720; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5722 = 8'h5a == io_state_in_6 ? 8'h8 : _GEN_5721; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5723 = 8'h5b == io_state_in_6 ? 8'h3 : _GEN_5722; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5724 = 8'h5c == io_state_in_6 ? 8'h32 : _GEN_5723; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5725 = 8'h5d == io_state_in_6 ? 8'h39 : _GEN_5724; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5726 = 8'h5e == io_state_in_6 ? 8'h24 : _GEN_5725; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5727 = 8'h5f == io_state_in_6 ? 8'h2f : _GEN_5726; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5728 = 8'h60 == io_state_in_6 ? 8'h8d : _GEN_5727; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5729 = 8'h61 == io_state_in_6 ? 8'h86 : _GEN_5728; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5730 = 8'h62 == io_state_in_6 ? 8'h9b : _GEN_5729; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5731 = 8'h63 == io_state_in_6 ? 8'h90 : _GEN_5730; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5732 = 8'h64 == io_state_in_6 ? 8'ha1 : _GEN_5731; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5733 = 8'h65 == io_state_in_6 ? 8'haa : _GEN_5732; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5734 = 8'h66 == io_state_in_6 ? 8'hb7 : _GEN_5733; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5735 = 8'h67 == io_state_in_6 ? 8'hbc : _GEN_5734; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5736 = 8'h68 == io_state_in_6 ? 8'hd5 : _GEN_5735; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5737 = 8'h69 == io_state_in_6 ? 8'hde : _GEN_5736; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5738 = 8'h6a == io_state_in_6 ? 8'hc3 : _GEN_5737; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5739 = 8'h6b == io_state_in_6 ? 8'hc8 : _GEN_5738; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5740 = 8'h6c == io_state_in_6 ? 8'hf9 : _GEN_5739; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5741 = 8'h6d == io_state_in_6 ? 8'hf2 : _GEN_5740; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5742 = 8'h6e == io_state_in_6 ? 8'hef : _GEN_5741; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5743 = 8'h6f == io_state_in_6 ? 8'he4 : _GEN_5742; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5744 = 8'h70 == io_state_in_6 ? 8'h3d : _GEN_5743; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5745 = 8'h71 == io_state_in_6 ? 8'h36 : _GEN_5744; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5746 = 8'h72 == io_state_in_6 ? 8'h2b : _GEN_5745; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5747 = 8'h73 == io_state_in_6 ? 8'h20 : _GEN_5746; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5748 = 8'h74 == io_state_in_6 ? 8'h11 : _GEN_5747; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5749 = 8'h75 == io_state_in_6 ? 8'h1a : _GEN_5748; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5750 = 8'h76 == io_state_in_6 ? 8'h7 : _GEN_5749; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5751 = 8'h77 == io_state_in_6 ? 8'hc : _GEN_5750; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5752 = 8'h78 == io_state_in_6 ? 8'h65 : _GEN_5751; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5753 = 8'h79 == io_state_in_6 ? 8'h6e : _GEN_5752; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5754 = 8'h7a == io_state_in_6 ? 8'h73 : _GEN_5753; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5755 = 8'h7b == io_state_in_6 ? 8'h78 : _GEN_5754; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5756 = 8'h7c == io_state_in_6 ? 8'h49 : _GEN_5755; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5757 = 8'h7d == io_state_in_6 ? 8'h42 : _GEN_5756; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5758 = 8'h7e == io_state_in_6 ? 8'h5f : _GEN_5757; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5759 = 8'h7f == io_state_in_6 ? 8'h54 : _GEN_5758; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5760 = 8'h80 == io_state_in_6 ? 8'hf7 : _GEN_5759; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5761 = 8'h81 == io_state_in_6 ? 8'hfc : _GEN_5760; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5762 = 8'h82 == io_state_in_6 ? 8'he1 : _GEN_5761; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5763 = 8'h83 == io_state_in_6 ? 8'hea : _GEN_5762; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5764 = 8'h84 == io_state_in_6 ? 8'hdb : _GEN_5763; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5765 = 8'h85 == io_state_in_6 ? 8'hd0 : _GEN_5764; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5766 = 8'h86 == io_state_in_6 ? 8'hcd : _GEN_5765; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5767 = 8'h87 == io_state_in_6 ? 8'hc6 : _GEN_5766; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5768 = 8'h88 == io_state_in_6 ? 8'haf : _GEN_5767; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5769 = 8'h89 == io_state_in_6 ? 8'ha4 : _GEN_5768; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5770 = 8'h8a == io_state_in_6 ? 8'hb9 : _GEN_5769; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5771 = 8'h8b == io_state_in_6 ? 8'hb2 : _GEN_5770; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5772 = 8'h8c == io_state_in_6 ? 8'h83 : _GEN_5771; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5773 = 8'h8d == io_state_in_6 ? 8'h88 : _GEN_5772; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5774 = 8'h8e == io_state_in_6 ? 8'h95 : _GEN_5773; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5775 = 8'h8f == io_state_in_6 ? 8'h9e : _GEN_5774; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5776 = 8'h90 == io_state_in_6 ? 8'h47 : _GEN_5775; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5777 = 8'h91 == io_state_in_6 ? 8'h4c : _GEN_5776; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5778 = 8'h92 == io_state_in_6 ? 8'h51 : _GEN_5777; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5779 = 8'h93 == io_state_in_6 ? 8'h5a : _GEN_5778; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5780 = 8'h94 == io_state_in_6 ? 8'h6b : _GEN_5779; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5781 = 8'h95 == io_state_in_6 ? 8'h60 : _GEN_5780; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5782 = 8'h96 == io_state_in_6 ? 8'h7d : _GEN_5781; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5783 = 8'h97 == io_state_in_6 ? 8'h76 : _GEN_5782; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5784 = 8'h98 == io_state_in_6 ? 8'h1f : _GEN_5783; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5785 = 8'h99 == io_state_in_6 ? 8'h14 : _GEN_5784; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5786 = 8'h9a == io_state_in_6 ? 8'h9 : _GEN_5785; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5787 = 8'h9b == io_state_in_6 ? 8'h2 : _GEN_5786; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5788 = 8'h9c == io_state_in_6 ? 8'h33 : _GEN_5787; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5789 = 8'h9d == io_state_in_6 ? 8'h38 : _GEN_5788; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5790 = 8'h9e == io_state_in_6 ? 8'h25 : _GEN_5789; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5791 = 8'h9f == io_state_in_6 ? 8'h2e : _GEN_5790; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5792 = 8'ha0 == io_state_in_6 ? 8'h8c : _GEN_5791; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5793 = 8'ha1 == io_state_in_6 ? 8'h87 : _GEN_5792; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5794 = 8'ha2 == io_state_in_6 ? 8'h9a : _GEN_5793; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5795 = 8'ha3 == io_state_in_6 ? 8'h91 : _GEN_5794; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5796 = 8'ha4 == io_state_in_6 ? 8'ha0 : _GEN_5795; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5797 = 8'ha5 == io_state_in_6 ? 8'hab : _GEN_5796; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5798 = 8'ha6 == io_state_in_6 ? 8'hb6 : _GEN_5797; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5799 = 8'ha7 == io_state_in_6 ? 8'hbd : _GEN_5798; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5800 = 8'ha8 == io_state_in_6 ? 8'hd4 : _GEN_5799; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5801 = 8'ha9 == io_state_in_6 ? 8'hdf : _GEN_5800; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5802 = 8'haa == io_state_in_6 ? 8'hc2 : _GEN_5801; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5803 = 8'hab == io_state_in_6 ? 8'hc9 : _GEN_5802; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5804 = 8'hac == io_state_in_6 ? 8'hf8 : _GEN_5803; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5805 = 8'had == io_state_in_6 ? 8'hf3 : _GEN_5804; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5806 = 8'hae == io_state_in_6 ? 8'hee : _GEN_5805; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5807 = 8'haf == io_state_in_6 ? 8'he5 : _GEN_5806; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5808 = 8'hb0 == io_state_in_6 ? 8'h3c : _GEN_5807; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5809 = 8'hb1 == io_state_in_6 ? 8'h37 : _GEN_5808; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5810 = 8'hb2 == io_state_in_6 ? 8'h2a : _GEN_5809; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5811 = 8'hb3 == io_state_in_6 ? 8'h21 : _GEN_5810; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5812 = 8'hb4 == io_state_in_6 ? 8'h10 : _GEN_5811; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5813 = 8'hb5 == io_state_in_6 ? 8'h1b : _GEN_5812; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5814 = 8'hb6 == io_state_in_6 ? 8'h6 : _GEN_5813; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5815 = 8'hb7 == io_state_in_6 ? 8'hd : _GEN_5814; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5816 = 8'hb8 == io_state_in_6 ? 8'h64 : _GEN_5815; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5817 = 8'hb9 == io_state_in_6 ? 8'h6f : _GEN_5816; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5818 = 8'hba == io_state_in_6 ? 8'h72 : _GEN_5817; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5819 = 8'hbb == io_state_in_6 ? 8'h79 : _GEN_5818; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5820 = 8'hbc == io_state_in_6 ? 8'h48 : _GEN_5819; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5821 = 8'hbd == io_state_in_6 ? 8'h43 : _GEN_5820; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5822 = 8'hbe == io_state_in_6 ? 8'h5e : _GEN_5821; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5823 = 8'hbf == io_state_in_6 ? 8'h55 : _GEN_5822; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5824 = 8'hc0 == io_state_in_6 ? 8'h1 : _GEN_5823; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5825 = 8'hc1 == io_state_in_6 ? 8'ha : _GEN_5824; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5826 = 8'hc2 == io_state_in_6 ? 8'h17 : _GEN_5825; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5827 = 8'hc3 == io_state_in_6 ? 8'h1c : _GEN_5826; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5828 = 8'hc4 == io_state_in_6 ? 8'h2d : _GEN_5827; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5829 = 8'hc5 == io_state_in_6 ? 8'h26 : _GEN_5828; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5830 = 8'hc6 == io_state_in_6 ? 8'h3b : _GEN_5829; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5831 = 8'hc7 == io_state_in_6 ? 8'h30 : _GEN_5830; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5832 = 8'hc8 == io_state_in_6 ? 8'h59 : _GEN_5831; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5833 = 8'hc9 == io_state_in_6 ? 8'h52 : _GEN_5832; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5834 = 8'hca == io_state_in_6 ? 8'h4f : _GEN_5833; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5835 = 8'hcb == io_state_in_6 ? 8'h44 : _GEN_5834; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5836 = 8'hcc == io_state_in_6 ? 8'h75 : _GEN_5835; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5837 = 8'hcd == io_state_in_6 ? 8'h7e : _GEN_5836; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5838 = 8'hce == io_state_in_6 ? 8'h63 : _GEN_5837; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5839 = 8'hcf == io_state_in_6 ? 8'h68 : _GEN_5838; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5840 = 8'hd0 == io_state_in_6 ? 8'hb1 : _GEN_5839; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5841 = 8'hd1 == io_state_in_6 ? 8'hba : _GEN_5840; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5842 = 8'hd2 == io_state_in_6 ? 8'ha7 : _GEN_5841; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5843 = 8'hd3 == io_state_in_6 ? 8'hac : _GEN_5842; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5844 = 8'hd4 == io_state_in_6 ? 8'h9d : _GEN_5843; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5845 = 8'hd5 == io_state_in_6 ? 8'h96 : _GEN_5844; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5846 = 8'hd6 == io_state_in_6 ? 8'h8b : _GEN_5845; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5847 = 8'hd7 == io_state_in_6 ? 8'h80 : _GEN_5846; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5848 = 8'hd8 == io_state_in_6 ? 8'he9 : _GEN_5847; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5849 = 8'hd9 == io_state_in_6 ? 8'he2 : _GEN_5848; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5850 = 8'hda == io_state_in_6 ? 8'hff : _GEN_5849; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5851 = 8'hdb == io_state_in_6 ? 8'hf4 : _GEN_5850; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5852 = 8'hdc == io_state_in_6 ? 8'hc5 : _GEN_5851; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5853 = 8'hdd == io_state_in_6 ? 8'hce : _GEN_5852; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5854 = 8'hde == io_state_in_6 ? 8'hd3 : _GEN_5853; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5855 = 8'hdf == io_state_in_6 ? 8'hd8 : _GEN_5854; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5856 = 8'he0 == io_state_in_6 ? 8'h7a : _GEN_5855; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5857 = 8'he1 == io_state_in_6 ? 8'h71 : _GEN_5856; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5858 = 8'he2 == io_state_in_6 ? 8'h6c : _GEN_5857; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5859 = 8'he3 == io_state_in_6 ? 8'h67 : _GEN_5858; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5860 = 8'he4 == io_state_in_6 ? 8'h56 : _GEN_5859; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5861 = 8'he5 == io_state_in_6 ? 8'h5d : _GEN_5860; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5862 = 8'he6 == io_state_in_6 ? 8'h40 : _GEN_5861; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5863 = 8'he7 == io_state_in_6 ? 8'h4b : _GEN_5862; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5864 = 8'he8 == io_state_in_6 ? 8'h22 : _GEN_5863; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5865 = 8'he9 == io_state_in_6 ? 8'h29 : _GEN_5864; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5866 = 8'hea == io_state_in_6 ? 8'h34 : _GEN_5865; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5867 = 8'heb == io_state_in_6 ? 8'h3f : _GEN_5866; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5868 = 8'hec == io_state_in_6 ? 8'he : _GEN_5867; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5869 = 8'hed == io_state_in_6 ? 8'h5 : _GEN_5868; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5870 = 8'hee == io_state_in_6 ? 8'h18 : _GEN_5869; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5871 = 8'hef == io_state_in_6 ? 8'h13 : _GEN_5870; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5872 = 8'hf0 == io_state_in_6 ? 8'hca : _GEN_5871; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5873 = 8'hf1 == io_state_in_6 ? 8'hc1 : _GEN_5872; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5874 = 8'hf2 == io_state_in_6 ? 8'hdc : _GEN_5873; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5875 = 8'hf3 == io_state_in_6 ? 8'hd7 : _GEN_5874; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5876 = 8'hf4 == io_state_in_6 ? 8'he6 : _GEN_5875; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5877 = 8'hf5 == io_state_in_6 ? 8'hed : _GEN_5876; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5878 = 8'hf6 == io_state_in_6 ? 8'hf0 : _GEN_5877; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5879 = 8'hf7 == io_state_in_6 ? 8'hfb : _GEN_5878; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5880 = 8'hf8 == io_state_in_6 ? 8'h92 : _GEN_5879; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5881 = 8'hf9 == io_state_in_6 ? 8'h99 : _GEN_5880; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5882 = 8'hfa == io_state_in_6 ? 8'h84 : _GEN_5881; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5883 = 8'hfb == io_state_in_6 ? 8'h8f : _GEN_5882; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5884 = 8'hfc == io_state_in_6 ? 8'hbe : _GEN_5883; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5885 = 8'hfd == io_state_in_6 ? 8'hb5 : _GEN_5884; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5886 = 8'hfe == io_state_in_6 ? 8'ha8 : _GEN_5885; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _GEN_5887 = 8'hff == io_state_in_6 ? 8'ha3 : _GEN_5886; // @[InvMixColumns.scala 132:{65,65}]
  wire [7:0] _tmp_state_5_T_1 = _tmp_state_5_T ^ _GEN_5887; // @[InvMixColumns.scala 132:65]
  wire [7:0] _GEN_5889 = 8'h1 == io_state_in_7 ? 8'hd : 8'h0; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5890 = 8'h2 == io_state_in_7 ? 8'h1a : _GEN_5889; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5891 = 8'h3 == io_state_in_7 ? 8'h17 : _GEN_5890; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5892 = 8'h4 == io_state_in_7 ? 8'h34 : _GEN_5891; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5893 = 8'h5 == io_state_in_7 ? 8'h39 : _GEN_5892; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5894 = 8'h6 == io_state_in_7 ? 8'h2e : _GEN_5893; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5895 = 8'h7 == io_state_in_7 ? 8'h23 : _GEN_5894; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5896 = 8'h8 == io_state_in_7 ? 8'h68 : _GEN_5895; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5897 = 8'h9 == io_state_in_7 ? 8'h65 : _GEN_5896; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5898 = 8'ha == io_state_in_7 ? 8'h72 : _GEN_5897; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5899 = 8'hb == io_state_in_7 ? 8'h7f : _GEN_5898; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5900 = 8'hc == io_state_in_7 ? 8'h5c : _GEN_5899; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5901 = 8'hd == io_state_in_7 ? 8'h51 : _GEN_5900; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5902 = 8'he == io_state_in_7 ? 8'h46 : _GEN_5901; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5903 = 8'hf == io_state_in_7 ? 8'h4b : _GEN_5902; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5904 = 8'h10 == io_state_in_7 ? 8'hd0 : _GEN_5903; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5905 = 8'h11 == io_state_in_7 ? 8'hdd : _GEN_5904; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5906 = 8'h12 == io_state_in_7 ? 8'hca : _GEN_5905; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5907 = 8'h13 == io_state_in_7 ? 8'hc7 : _GEN_5906; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5908 = 8'h14 == io_state_in_7 ? 8'he4 : _GEN_5907; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5909 = 8'h15 == io_state_in_7 ? 8'he9 : _GEN_5908; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5910 = 8'h16 == io_state_in_7 ? 8'hfe : _GEN_5909; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5911 = 8'h17 == io_state_in_7 ? 8'hf3 : _GEN_5910; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5912 = 8'h18 == io_state_in_7 ? 8'hb8 : _GEN_5911; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5913 = 8'h19 == io_state_in_7 ? 8'hb5 : _GEN_5912; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5914 = 8'h1a == io_state_in_7 ? 8'ha2 : _GEN_5913; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5915 = 8'h1b == io_state_in_7 ? 8'haf : _GEN_5914; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5916 = 8'h1c == io_state_in_7 ? 8'h8c : _GEN_5915; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5917 = 8'h1d == io_state_in_7 ? 8'h81 : _GEN_5916; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5918 = 8'h1e == io_state_in_7 ? 8'h96 : _GEN_5917; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5919 = 8'h1f == io_state_in_7 ? 8'h9b : _GEN_5918; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5920 = 8'h20 == io_state_in_7 ? 8'hbb : _GEN_5919; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5921 = 8'h21 == io_state_in_7 ? 8'hb6 : _GEN_5920; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5922 = 8'h22 == io_state_in_7 ? 8'ha1 : _GEN_5921; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5923 = 8'h23 == io_state_in_7 ? 8'hac : _GEN_5922; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5924 = 8'h24 == io_state_in_7 ? 8'h8f : _GEN_5923; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5925 = 8'h25 == io_state_in_7 ? 8'h82 : _GEN_5924; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5926 = 8'h26 == io_state_in_7 ? 8'h95 : _GEN_5925; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5927 = 8'h27 == io_state_in_7 ? 8'h98 : _GEN_5926; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5928 = 8'h28 == io_state_in_7 ? 8'hd3 : _GEN_5927; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5929 = 8'h29 == io_state_in_7 ? 8'hde : _GEN_5928; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5930 = 8'h2a == io_state_in_7 ? 8'hc9 : _GEN_5929; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5931 = 8'h2b == io_state_in_7 ? 8'hc4 : _GEN_5930; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5932 = 8'h2c == io_state_in_7 ? 8'he7 : _GEN_5931; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5933 = 8'h2d == io_state_in_7 ? 8'hea : _GEN_5932; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5934 = 8'h2e == io_state_in_7 ? 8'hfd : _GEN_5933; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5935 = 8'h2f == io_state_in_7 ? 8'hf0 : _GEN_5934; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5936 = 8'h30 == io_state_in_7 ? 8'h6b : _GEN_5935; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5937 = 8'h31 == io_state_in_7 ? 8'h66 : _GEN_5936; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5938 = 8'h32 == io_state_in_7 ? 8'h71 : _GEN_5937; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5939 = 8'h33 == io_state_in_7 ? 8'h7c : _GEN_5938; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5940 = 8'h34 == io_state_in_7 ? 8'h5f : _GEN_5939; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5941 = 8'h35 == io_state_in_7 ? 8'h52 : _GEN_5940; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5942 = 8'h36 == io_state_in_7 ? 8'h45 : _GEN_5941; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5943 = 8'h37 == io_state_in_7 ? 8'h48 : _GEN_5942; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5944 = 8'h38 == io_state_in_7 ? 8'h3 : _GEN_5943; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5945 = 8'h39 == io_state_in_7 ? 8'he : _GEN_5944; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5946 = 8'h3a == io_state_in_7 ? 8'h19 : _GEN_5945; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5947 = 8'h3b == io_state_in_7 ? 8'h14 : _GEN_5946; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5948 = 8'h3c == io_state_in_7 ? 8'h37 : _GEN_5947; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5949 = 8'h3d == io_state_in_7 ? 8'h3a : _GEN_5948; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5950 = 8'h3e == io_state_in_7 ? 8'h2d : _GEN_5949; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5951 = 8'h3f == io_state_in_7 ? 8'h20 : _GEN_5950; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5952 = 8'h40 == io_state_in_7 ? 8'h6d : _GEN_5951; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5953 = 8'h41 == io_state_in_7 ? 8'h60 : _GEN_5952; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5954 = 8'h42 == io_state_in_7 ? 8'h77 : _GEN_5953; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5955 = 8'h43 == io_state_in_7 ? 8'h7a : _GEN_5954; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5956 = 8'h44 == io_state_in_7 ? 8'h59 : _GEN_5955; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5957 = 8'h45 == io_state_in_7 ? 8'h54 : _GEN_5956; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5958 = 8'h46 == io_state_in_7 ? 8'h43 : _GEN_5957; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5959 = 8'h47 == io_state_in_7 ? 8'h4e : _GEN_5958; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5960 = 8'h48 == io_state_in_7 ? 8'h5 : _GEN_5959; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5961 = 8'h49 == io_state_in_7 ? 8'h8 : _GEN_5960; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5962 = 8'h4a == io_state_in_7 ? 8'h1f : _GEN_5961; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5963 = 8'h4b == io_state_in_7 ? 8'h12 : _GEN_5962; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5964 = 8'h4c == io_state_in_7 ? 8'h31 : _GEN_5963; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5965 = 8'h4d == io_state_in_7 ? 8'h3c : _GEN_5964; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5966 = 8'h4e == io_state_in_7 ? 8'h2b : _GEN_5965; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5967 = 8'h4f == io_state_in_7 ? 8'h26 : _GEN_5966; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5968 = 8'h50 == io_state_in_7 ? 8'hbd : _GEN_5967; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5969 = 8'h51 == io_state_in_7 ? 8'hb0 : _GEN_5968; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5970 = 8'h52 == io_state_in_7 ? 8'ha7 : _GEN_5969; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5971 = 8'h53 == io_state_in_7 ? 8'haa : _GEN_5970; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5972 = 8'h54 == io_state_in_7 ? 8'h89 : _GEN_5971; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5973 = 8'h55 == io_state_in_7 ? 8'h84 : _GEN_5972; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5974 = 8'h56 == io_state_in_7 ? 8'h93 : _GEN_5973; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5975 = 8'h57 == io_state_in_7 ? 8'h9e : _GEN_5974; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5976 = 8'h58 == io_state_in_7 ? 8'hd5 : _GEN_5975; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5977 = 8'h59 == io_state_in_7 ? 8'hd8 : _GEN_5976; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5978 = 8'h5a == io_state_in_7 ? 8'hcf : _GEN_5977; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5979 = 8'h5b == io_state_in_7 ? 8'hc2 : _GEN_5978; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5980 = 8'h5c == io_state_in_7 ? 8'he1 : _GEN_5979; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5981 = 8'h5d == io_state_in_7 ? 8'hec : _GEN_5980; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5982 = 8'h5e == io_state_in_7 ? 8'hfb : _GEN_5981; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5983 = 8'h5f == io_state_in_7 ? 8'hf6 : _GEN_5982; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5984 = 8'h60 == io_state_in_7 ? 8'hd6 : _GEN_5983; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5985 = 8'h61 == io_state_in_7 ? 8'hdb : _GEN_5984; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5986 = 8'h62 == io_state_in_7 ? 8'hcc : _GEN_5985; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5987 = 8'h63 == io_state_in_7 ? 8'hc1 : _GEN_5986; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5988 = 8'h64 == io_state_in_7 ? 8'he2 : _GEN_5987; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5989 = 8'h65 == io_state_in_7 ? 8'hef : _GEN_5988; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5990 = 8'h66 == io_state_in_7 ? 8'hf8 : _GEN_5989; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5991 = 8'h67 == io_state_in_7 ? 8'hf5 : _GEN_5990; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5992 = 8'h68 == io_state_in_7 ? 8'hbe : _GEN_5991; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5993 = 8'h69 == io_state_in_7 ? 8'hb3 : _GEN_5992; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5994 = 8'h6a == io_state_in_7 ? 8'ha4 : _GEN_5993; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5995 = 8'h6b == io_state_in_7 ? 8'ha9 : _GEN_5994; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5996 = 8'h6c == io_state_in_7 ? 8'h8a : _GEN_5995; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5997 = 8'h6d == io_state_in_7 ? 8'h87 : _GEN_5996; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5998 = 8'h6e == io_state_in_7 ? 8'h90 : _GEN_5997; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_5999 = 8'h6f == io_state_in_7 ? 8'h9d : _GEN_5998; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6000 = 8'h70 == io_state_in_7 ? 8'h6 : _GEN_5999; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6001 = 8'h71 == io_state_in_7 ? 8'hb : _GEN_6000; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6002 = 8'h72 == io_state_in_7 ? 8'h1c : _GEN_6001; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6003 = 8'h73 == io_state_in_7 ? 8'h11 : _GEN_6002; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6004 = 8'h74 == io_state_in_7 ? 8'h32 : _GEN_6003; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6005 = 8'h75 == io_state_in_7 ? 8'h3f : _GEN_6004; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6006 = 8'h76 == io_state_in_7 ? 8'h28 : _GEN_6005; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6007 = 8'h77 == io_state_in_7 ? 8'h25 : _GEN_6006; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6008 = 8'h78 == io_state_in_7 ? 8'h6e : _GEN_6007; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6009 = 8'h79 == io_state_in_7 ? 8'h63 : _GEN_6008; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6010 = 8'h7a == io_state_in_7 ? 8'h74 : _GEN_6009; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6011 = 8'h7b == io_state_in_7 ? 8'h79 : _GEN_6010; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6012 = 8'h7c == io_state_in_7 ? 8'h5a : _GEN_6011; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6013 = 8'h7d == io_state_in_7 ? 8'h57 : _GEN_6012; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6014 = 8'h7e == io_state_in_7 ? 8'h40 : _GEN_6013; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6015 = 8'h7f == io_state_in_7 ? 8'h4d : _GEN_6014; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6016 = 8'h80 == io_state_in_7 ? 8'hda : _GEN_6015; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6017 = 8'h81 == io_state_in_7 ? 8'hd7 : _GEN_6016; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6018 = 8'h82 == io_state_in_7 ? 8'hc0 : _GEN_6017; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6019 = 8'h83 == io_state_in_7 ? 8'hcd : _GEN_6018; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6020 = 8'h84 == io_state_in_7 ? 8'hee : _GEN_6019; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6021 = 8'h85 == io_state_in_7 ? 8'he3 : _GEN_6020; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6022 = 8'h86 == io_state_in_7 ? 8'hf4 : _GEN_6021; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6023 = 8'h87 == io_state_in_7 ? 8'hf9 : _GEN_6022; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6024 = 8'h88 == io_state_in_7 ? 8'hb2 : _GEN_6023; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6025 = 8'h89 == io_state_in_7 ? 8'hbf : _GEN_6024; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6026 = 8'h8a == io_state_in_7 ? 8'ha8 : _GEN_6025; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6027 = 8'h8b == io_state_in_7 ? 8'ha5 : _GEN_6026; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6028 = 8'h8c == io_state_in_7 ? 8'h86 : _GEN_6027; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6029 = 8'h8d == io_state_in_7 ? 8'h8b : _GEN_6028; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6030 = 8'h8e == io_state_in_7 ? 8'h9c : _GEN_6029; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6031 = 8'h8f == io_state_in_7 ? 8'h91 : _GEN_6030; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6032 = 8'h90 == io_state_in_7 ? 8'ha : _GEN_6031; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6033 = 8'h91 == io_state_in_7 ? 8'h7 : _GEN_6032; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6034 = 8'h92 == io_state_in_7 ? 8'h10 : _GEN_6033; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6035 = 8'h93 == io_state_in_7 ? 8'h1d : _GEN_6034; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6036 = 8'h94 == io_state_in_7 ? 8'h3e : _GEN_6035; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6037 = 8'h95 == io_state_in_7 ? 8'h33 : _GEN_6036; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6038 = 8'h96 == io_state_in_7 ? 8'h24 : _GEN_6037; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6039 = 8'h97 == io_state_in_7 ? 8'h29 : _GEN_6038; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6040 = 8'h98 == io_state_in_7 ? 8'h62 : _GEN_6039; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6041 = 8'h99 == io_state_in_7 ? 8'h6f : _GEN_6040; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6042 = 8'h9a == io_state_in_7 ? 8'h78 : _GEN_6041; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6043 = 8'h9b == io_state_in_7 ? 8'h75 : _GEN_6042; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6044 = 8'h9c == io_state_in_7 ? 8'h56 : _GEN_6043; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6045 = 8'h9d == io_state_in_7 ? 8'h5b : _GEN_6044; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6046 = 8'h9e == io_state_in_7 ? 8'h4c : _GEN_6045; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6047 = 8'h9f == io_state_in_7 ? 8'h41 : _GEN_6046; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6048 = 8'ha0 == io_state_in_7 ? 8'h61 : _GEN_6047; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6049 = 8'ha1 == io_state_in_7 ? 8'h6c : _GEN_6048; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6050 = 8'ha2 == io_state_in_7 ? 8'h7b : _GEN_6049; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6051 = 8'ha3 == io_state_in_7 ? 8'h76 : _GEN_6050; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6052 = 8'ha4 == io_state_in_7 ? 8'h55 : _GEN_6051; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6053 = 8'ha5 == io_state_in_7 ? 8'h58 : _GEN_6052; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6054 = 8'ha6 == io_state_in_7 ? 8'h4f : _GEN_6053; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6055 = 8'ha7 == io_state_in_7 ? 8'h42 : _GEN_6054; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6056 = 8'ha8 == io_state_in_7 ? 8'h9 : _GEN_6055; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6057 = 8'ha9 == io_state_in_7 ? 8'h4 : _GEN_6056; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6058 = 8'haa == io_state_in_7 ? 8'h13 : _GEN_6057; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6059 = 8'hab == io_state_in_7 ? 8'h1e : _GEN_6058; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6060 = 8'hac == io_state_in_7 ? 8'h3d : _GEN_6059; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6061 = 8'had == io_state_in_7 ? 8'h30 : _GEN_6060; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6062 = 8'hae == io_state_in_7 ? 8'h27 : _GEN_6061; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6063 = 8'haf == io_state_in_7 ? 8'h2a : _GEN_6062; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6064 = 8'hb0 == io_state_in_7 ? 8'hb1 : _GEN_6063; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6065 = 8'hb1 == io_state_in_7 ? 8'hbc : _GEN_6064; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6066 = 8'hb2 == io_state_in_7 ? 8'hab : _GEN_6065; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6067 = 8'hb3 == io_state_in_7 ? 8'ha6 : _GEN_6066; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6068 = 8'hb4 == io_state_in_7 ? 8'h85 : _GEN_6067; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6069 = 8'hb5 == io_state_in_7 ? 8'h88 : _GEN_6068; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6070 = 8'hb6 == io_state_in_7 ? 8'h9f : _GEN_6069; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6071 = 8'hb7 == io_state_in_7 ? 8'h92 : _GEN_6070; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6072 = 8'hb8 == io_state_in_7 ? 8'hd9 : _GEN_6071; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6073 = 8'hb9 == io_state_in_7 ? 8'hd4 : _GEN_6072; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6074 = 8'hba == io_state_in_7 ? 8'hc3 : _GEN_6073; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6075 = 8'hbb == io_state_in_7 ? 8'hce : _GEN_6074; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6076 = 8'hbc == io_state_in_7 ? 8'hed : _GEN_6075; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6077 = 8'hbd == io_state_in_7 ? 8'he0 : _GEN_6076; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6078 = 8'hbe == io_state_in_7 ? 8'hf7 : _GEN_6077; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6079 = 8'hbf == io_state_in_7 ? 8'hfa : _GEN_6078; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6080 = 8'hc0 == io_state_in_7 ? 8'hb7 : _GEN_6079; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6081 = 8'hc1 == io_state_in_7 ? 8'hba : _GEN_6080; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6082 = 8'hc2 == io_state_in_7 ? 8'had : _GEN_6081; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6083 = 8'hc3 == io_state_in_7 ? 8'ha0 : _GEN_6082; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6084 = 8'hc4 == io_state_in_7 ? 8'h83 : _GEN_6083; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6085 = 8'hc5 == io_state_in_7 ? 8'h8e : _GEN_6084; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6086 = 8'hc6 == io_state_in_7 ? 8'h99 : _GEN_6085; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6087 = 8'hc7 == io_state_in_7 ? 8'h94 : _GEN_6086; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6088 = 8'hc8 == io_state_in_7 ? 8'hdf : _GEN_6087; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6089 = 8'hc9 == io_state_in_7 ? 8'hd2 : _GEN_6088; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6090 = 8'hca == io_state_in_7 ? 8'hc5 : _GEN_6089; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6091 = 8'hcb == io_state_in_7 ? 8'hc8 : _GEN_6090; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6092 = 8'hcc == io_state_in_7 ? 8'heb : _GEN_6091; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6093 = 8'hcd == io_state_in_7 ? 8'he6 : _GEN_6092; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6094 = 8'hce == io_state_in_7 ? 8'hf1 : _GEN_6093; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6095 = 8'hcf == io_state_in_7 ? 8'hfc : _GEN_6094; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6096 = 8'hd0 == io_state_in_7 ? 8'h67 : _GEN_6095; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6097 = 8'hd1 == io_state_in_7 ? 8'h6a : _GEN_6096; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6098 = 8'hd2 == io_state_in_7 ? 8'h7d : _GEN_6097; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6099 = 8'hd3 == io_state_in_7 ? 8'h70 : _GEN_6098; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6100 = 8'hd4 == io_state_in_7 ? 8'h53 : _GEN_6099; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6101 = 8'hd5 == io_state_in_7 ? 8'h5e : _GEN_6100; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6102 = 8'hd6 == io_state_in_7 ? 8'h49 : _GEN_6101; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6103 = 8'hd7 == io_state_in_7 ? 8'h44 : _GEN_6102; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6104 = 8'hd8 == io_state_in_7 ? 8'hf : _GEN_6103; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6105 = 8'hd9 == io_state_in_7 ? 8'h2 : _GEN_6104; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6106 = 8'hda == io_state_in_7 ? 8'h15 : _GEN_6105; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6107 = 8'hdb == io_state_in_7 ? 8'h18 : _GEN_6106; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6108 = 8'hdc == io_state_in_7 ? 8'h3b : _GEN_6107; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6109 = 8'hdd == io_state_in_7 ? 8'h36 : _GEN_6108; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6110 = 8'hde == io_state_in_7 ? 8'h21 : _GEN_6109; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6111 = 8'hdf == io_state_in_7 ? 8'h2c : _GEN_6110; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6112 = 8'he0 == io_state_in_7 ? 8'hc : _GEN_6111; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6113 = 8'he1 == io_state_in_7 ? 8'h1 : _GEN_6112; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6114 = 8'he2 == io_state_in_7 ? 8'h16 : _GEN_6113; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6115 = 8'he3 == io_state_in_7 ? 8'h1b : _GEN_6114; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6116 = 8'he4 == io_state_in_7 ? 8'h38 : _GEN_6115; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6117 = 8'he5 == io_state_in_7 ? 8'h35 : _GEN_6116; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6118 = 8'he6 == io_state_in_7 ? 8'h22 : _GEN_6117; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6119 = 8'he7 == io_state_in_7 ? 8'h2f : _GEN_6118; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6120 = 8'he8 == io_state_in_7 ? 8'h64 : _GEN_6119; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6121 = 8'he9 == io_state_in_7 ? 8'h69 : _GEN_6120; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6122 = 8'hea == io_state_in_7 ? 8'h7e : _GEN_6121; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6123 = 8'heb == io_state_in_7 ? 8'h73 : _GEN_6122; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6124 = 8'hec == io_state_in_7 ? 8'h50 : _GEN_6123; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6125 = 8'hed == io_state_in_7 ? 8'h5d : _GEN_6124; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6126 = 8'hee == io_state_in_7 ? 8'h4a : _GEN_6125; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6127 = 8'hef == io_state_in_7 ? 8'h47 : _GEN_6126; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6128 = 8'hf0 == io_state_in_7 ? 8'hdc : _GEN_6127; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6129 = 8'hf1 == io_state_in_7 ? 8'hd1 : _GEN_6128; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6130 = 8'hf2 == io_state_in_7 ? 8'hc6 : _GEN_6129; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6131 = 8'hf3 == io_state_in_7 ? 8'hcb : _GEN_6130; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6132 = 8'hf4 == io_state_in_7 ? 8'he8 : _GEN_6131; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6133 = 8'hf5 == io_state_in_7 ? 8'he5 : _GEN_6132; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6134 = 8'hf6 == io_state_in_7 ? 8'hf2 : _GEN_6133; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6135 = 8'hf7 == io_state_in_7 ? 8'hff : _GEN_6134; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6136 = 8'hf8 == io_state_in_7 ? 8'hb4 : _GEN_6135; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6137 = 8'hf9 == io_state_in_7 ? 8'hb9 : _GEN_6136; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6138 = 8'hfa == io_state_in_7 ? 8'hae : _GEN_6137; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6139 = 8'hfb == io_state_in_7 ? 8'ha3 : _GEN_6138; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6140 = 8'hfc == io_state_in_7 ? 8'h80 : _GEN_6139; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6141 = 8'hfd == io_state_in_7 ? 8'h8d : _GEN_6140; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6142 = 8'hfe == io_state_in_7 ? 8'h9a : _GEN_6141; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6143 = 8'hff == io_state_in_7 ? 8'h97 : _GEN_6142; // @[InvMixColumns.scala 132:{89,89}]
  wire [7:0] _GEN_6145 = 8'h1 == io_state_in_4 ? 8'hd : 8'h0; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6146 = 8'h2 == io_state_in_4 ? 8'h1a : _GEN_6145; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6147 = 8'h3 == io_state_in_4 ? 8'h17 : _GEN_6146; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6148 = 8'h4 == io_state_in_4 ? 8'h34 : _GEN_6147; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6149 = 8'h5 == io_state_in_4 ? 8'h39 : _GEN_6148; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6150 = 8'h6 == io_state_in_4 ? 8'h2e : _GEN_6149; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6151 = 8'h7 == io_state_in_4 ? 8'h23 : _GEN_6150; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6152 = 8'h8 == io_state_in_4 ? 8'h68 : _GEN_6151; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6153 = 8'h9 == io_state_in_4 ? 8'h65 : _GEN_6152; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6154 = 8'ha == io_state_in_4 ? 8'h72 : _GEN_6153; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6155 = 8'hb == io_state_in_4 ? 8'h7f : _GEN_6154; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6156 = 8'hc == io_state_in_4 ? 8'h5c : _GEN_6155; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6157 = 8'hd == io_state_in_4 ? 8'h51 : _GEN_6156; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6158 = 8'he == io_state_in_4 ? 8'h46 : _GEN_6157; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6159 = 8'hf == io_state_in_4 ? 8'h4b : _GEN_6158; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6160 = 8'h10 == io_state_in_4 ? 8'hd0 : _GEN_6159; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6161 = 8'h11 == io_state_in_4 ? 8'hdd : _GEN_6160; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6162 = 8'h12 == io_state_in_4 ? 8'hca : _GEN_6161; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6163 = 8'h13 == io_state_in_4 ? 8'hc7 : _GEN_6162; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6164 = 8'h14 == io_state_in_4 ? 8'he4 : _GEN_6163; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6165 = 8'h15 == io_state_in_4 ? 8'he9 : _GEN_6164; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6166 = 8'h16 == io_state_in_4 ? 8'hfe : _GEN_6165; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6167 = 8'h17 == io_state_in_4 ? 8'hf3 : _GEN_6166; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6168 = 8'h18 == io_state_in_4 ? 8'hb8 : _GEN_6167; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6169 = 8'h19 == io_state_in_4 ? 8'hb5 : _GEN_6168; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6170 = 8'h1a == io_state_in_4 ? 8'ha2 : _GEN_6169; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6171 = 8'h1b == io_state_in_4 ? 8'haf : _GEN_6170; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6172 = 8'h1c == io_state_in_4 ? 8'h8c : _GEN_6171; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6173 = 8'h1d == io_state_in_4 ? 8'h81 : _GEN_6172; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6174 = 8'h1e == io_state_in_4 ? 8'h96 : _GEN_6173; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6175 = 8'h1f == io_state_in_4 ? 8'h9b : _GEN_6174; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6176 = 8'h20 == io_state_in_4 ? 8'hbb : _GEN_6175; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6177 = 8'h21 == io_state_in_4 ? 8'hb6 : _GEN_6176; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6178 = 8'h22 == io_state_in_4 ? 8'ha1 : _GEN_6177; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6179 = 8'h23 == io_state_in_4 ? 8'hac : _GEN_6178; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6180 = 8'h24 == io_state_in_4 ? 8'h8f : _GEN_6179; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6181 = 8'h25 == io_state_in_4 ? 8'h82 : _GEN_6180; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6182 = 8'h26 == io_state_in_4 ? 8'h95 : _GEN_6181; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6183 = 8'h27 == io_state_in_4 ? 8'h98 : _GEN_6182; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6184 = 8'h28 == io_state_in_4 ? 8'hd3 : _GEN_6183; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6185 = 8'h29 == io_state_in_4 ? 8'hde : _GEN_6184; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6186 = 8'h2a == io_state_in_4 ? 8'hc9 : _GEN_6185; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6187 = 8'h2b == io_state_in_4 ? 8'hc4 : _GEN_6186; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6188 = 8'h2c == io_state_in_4 ? 8'he7 : _GEN_6187; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6189 = 8'h2d == io_state_in_4 ? 8'hea : _GEN_6188; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6190 = 8'h2e == io_state_in_4 ? 8'hfd : _GEN_6189; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6191 = 8'h2f == io_state_in_4 ? 8'hf0 : _GEN_6190; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6192 = 8'h30 == io_state_in_4 ? 8'h6b : _GEN_6191; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6193 = 8'h31 == io_state_in_4 ? 8'h66 : _GEN_6192; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6194 = 8'h32 == io_state_in_4 ? 8'h71 : _GEN_6193; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6195 = 8'h33 == io_state_in_4 ? 8'h7c : _GEN_6194; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6196 = 8'h34 == io_state_in_4 ? 8'h5f : _GEN_6195; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6197 = 8'h35 == io_state_in_4 ? 8'h52 : _GEN_6196; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6198 = 8'h36 == io_state_in_4 ? 8'h45 : _GEN_6197; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6199 = 8'h37 == io_state_in_4 ? 8'h48 : _GEN_6198; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6200 = 8'h38 == io_state_in_4 ? 8'h3 : _GEN_6199; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6201 = 8'h39 == io_state_in_4 ? 8'he : _GEN_6200; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6202 = 8'h3a == io_state_in_4 ? 8'h19 : _GEN_6201; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6203 = 8'h3b == io_state_in_4 ? 8'h14 : _GEN_6202; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6204 = 8'h3c == io_state_in_4 ? 8'h37 : _GEN_6203; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6205 = 8'h3d == io_state_in_4 ? 8'h3a : _GEN_6204; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6206 = 8'h3e == io_state_in_4 ? 8'h2d : _GEN_6205; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6207 = 8'h3f == io_state_in_4 ? 8'h20 : _GEN_6206; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6208 = 8'h40 == io_state_in_4 ? 8'h6d : _GEN_6207; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6209 = 8'h41 == io_state_in_4 ? 8'h60 : _GEN_6208; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6210 = 8'h42 == io_state_in_4 ? 8'h77 : _GEN_6209; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6211 = 8'h43 == io_state_in_4 ? 8'h7a : _GEN_6210; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6212 = 8'h44 == io_state_in_4 ? 8'h59 : _GEN_6211; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6213 = 8'h45 == io_state_in_4 ? 8'h54 : _GEN_6212; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6214 = 8'h46 == io_state_in_4 ? 8'h43 : _GEN_6213; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6215 = 8'h47 == io_state_in_4 ? 8'h4e : _GEN_6214; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6216 = 8'h48 == io_state_in_4 ? 8'h5 : _GEN_6215; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6217 = 8'h49 == io_state_in_4 ? 8'h8 : _GEN_6216; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6218 = 8'h4a == io_state_in_4 ? 8'h1f : _GEN_6217; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6219 = 8'h4b == io_state_in_4 ? 8'h12 : _GEN_6218; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6220 = 8'h4c == io_state_in_4 ? 8'h31 : _GEN_6219; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6221 = 8'h4d == io_state_in_4 ? 8'h3c : _GEN_6220; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6222 = 8'h4e == io_state_in_4 ? 8'h2b : _GEN_6221; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6223 = 8'h4f == io_state_in_4 ? 8'h26 : _GEN_6222; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6224 = 8'h50 == io_state_in_4 ? 8'hbd : _GEN_6223; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6225 = 8'h51 == io_state_in_4 ? 8'hb0 : _GEN_6224; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6226 = 8'h52 == io_state_in_4 ? 8'ha7 : _GEN_6225; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6227 = 8'h53 == io_state_in_4 ? 8'haa : _GEN_6226; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6228 = 8'h54 == io_state_in_4 ? 8'h89 : _GEN_6227; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6229 = 8'h55 == io_state_in_4 ? 8'h84 : _GEN_6228; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6230 = 8'h56 == io_state_in_4 ? 8'h93 : _GEN_6229; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6231 = 8'h57 == io_state_in_4 ? 8'h9e : _GEN_6230; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6232 = 8'h58 == io_state_in_4 ? 8'hd5 : _GEN_6231; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6233 = 8'h59 == io_state_in_4 ? 8'hd8 : _GEN_6232; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6234 = 8'h5a == io_state_in_4 ? 8'hcf : _GEN_6233; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6235 = 8'h5b == io_state_in_4 ? 8'hc2 : _GEN_6234; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6236 = 8'h5c == io_state_in_4 ? 8'he1 : _GEN_6235; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6237 = 8'h5d == io_state_in_4 ? 8'hec : _GEN_6236; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6238 = 8'h5e == io_state_in_4 ? 8'hfb : _GEN_6237; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6239 = 8'h5f == io_state_in_4 ? 8'hf6 : _GEN_6238; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6240 = 8'h60 == io_state_in_4 ? 8'hd6 : _GEN_6239; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6241 = 8'h61 == io_state_in_4 ? 8'hdb : _GEN_6240; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6242 = 8'h62 == io_state_in_4 ? 8'hcc : _GEN_6241; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6243 = 8'h63 == io_state_in_4 ? 8'hc1 : _GEN_6242; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6244 = 8'h64 == io_state_in_4 ? 8'he2 : _GEN_6243; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6245 = 8'h65 == io_state_in_4 ? 8'hef : _GEN_6244; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6246 = 8'h66 == io_state_in_4 ? 8'hf8 : _GEN_6245; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6247 = 8'h67 == io_state_in_4 ? 8'hf5 : _GEN_6246; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6248 = 8'h68 == io_state_in_4 ? 8'hbe : _GEN_6247; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6249 = 8'h69 == io_state_in_4 ? 8'hb3 : _GEN_6248; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6250 = 8'h6a == io_state_in_4 ? 8'ha4 : _GEN_6249; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6251 = 8'h6b == io_state_in_4 ? 8'ha9 : _GEN_6250; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6252 = 8'h6c == io_state_in_4 ? 8'h8a : _GEN_6251; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6253 = 8'h6d == io_state_in_4 ? 8'h87 : _GEN_6252; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6254 = 8'h6e == io_state_in_4 ? 8'h90 : _GEN_6253; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6255 = 8'h6f == io_state_in_4 ? 8'h9d : _GEN_6254; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6256 = 8'h70 == io_state_in_4 ? 8'h6 : _GEN_6255; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6257 = 8'h71 == io_state_in_4 ? 8'hb : _GEN_6256; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6258 = 8'h72 == io_state_in_4 ? 8'h1c : _GEN_6257; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6259 = 8'h73 == io_state_in_4 ? 8'h11 : _GEN_6258; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6260 = 8'h74 == io_state_in_4 ? 8'h32 : _GEN_6259; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6261 = 8'h75 == io_state_in_4 ? 8'h3f : _GEN_6260; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6262 = 8'h76 == io_state_in_4 ? 8'h28 : _GEN_6261; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6263 = 8'h77 == io_state_in_4 ? 8'h25 : _GEN_6262; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6264 = 8'h78 == io_state_in_4 ? 8'h6e : _GEN_6263; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6265 = 8'h79 == io_state_in_4 ? 8'h63 : _GEN_6264; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6266 = 8'h7a == io_state_in_4 ? 8'h74 : _GEN_6265; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6267 = 8'h7b == io_state_in_4 ? 8'h79 : _GEN_6266; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6268 = 8'h7c == io_state_in_4 ? 8'h5a : _GEN_6267; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6269 = 8'h7d == io_state_in_4 ? 8'h57 : _GEN_6268; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6270 = 8'h7e == io_state_in_4 ? 8'h40 : _GEN_6269; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6271 = 8'h7f == io_state_in_4 ? 8'h4d : _GEN_6270; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6272 = 8'h80 == io_state_in_4 ? 8'hda : _GEN_6271; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6273 = 8'h81 == io_state_in_4 ? 8'hd7 : _GEN_6272; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6274 = 8'h82 == io_state_in_4 ? 8'hc0 : _GEN_6273; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6275 = 8'h83 == io_state_in_4 ? 8'hcd : _GEN_6274; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6276 = 8'h84 == io_state_in_4 ? 8'hee : _GEN_6275; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6277 = 8'h85 == io_state_in_4 ? 8'he3 : _GEN_6276; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6278 = 8'h86 == io_state_in_4 ? 8'hf4 : _GEN_6277; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6279 = 8'h87 == io_state_in_4 ? 8'hf9 : _GEN_6278; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6280 = 8'h88 == io_state_in_4 ? 8'hb2 : _GEN_6279; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6281 = 8'h89 == io_state_in_4 ? 8'hbf : _GEN_6280; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6282 = 8'h8a == io_state_in_4 ? 8'ha8 : _GEN_6281; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6283 = 8'h8b == io_state_in_4 ? 8'ha5 : _GEN_6282; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6284 = 8'h8c == io_state_in_4 ? 8'h86 : _GEN_6283; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6285 = 8'h8d == io_state_in_4 ? 8'h8b : _GEN_6284; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6286 = 8'h8e == io_state_in_4 ? 8'h9c : _GEN_6285; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6287 = 8'h8f == io_state_in_4 ? 8'h91 : _GEN_6286; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6288 = 8'h90 == io_state_in_4 ? 8'ha : _GEN_6287; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6289 = 8'h91 == io_state_in_4 ? 8'h7 : _GEN_6288; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6290 = 8'h92 == io_state_in_4 ? 8'h10 : _GEN_6289; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6291 = 8'h93 == io_state_in_4 ? 8'h1d : _GEN_6290; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6292 = 8'h94 == io_state_in_4 ? 8'h3e : _GEN_6291; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6293 = 8'h95 == io_state_in_4 ? 8'h33 : _GEN_6292; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6294 = 8'h96 == io_state_in_4 ? 8'h24 : _GEN_6293; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6295 = 8'h97 == io_state_in_4 ? 8'h29 : _GEN_6294; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6296 = 8'h98 == io_state_in_4 ? 8'h62 : _GEN_6295; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6297 = 8'h99 == io_state_in_4 ? 8'h6f : _GEN_6296; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6298 = 8'h9a == io_state_in_4 ? 8'h78 : _GEN_6297; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6299 = 8'h9b == io_state_in_4 ? 8'h75 : _GEN_6298; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6300 = 8'h9c == io_state_in_4 ? 8'h56 : _GEN_6299; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6301 = 8'h9d == io_state_in_4 ? 8'h5b : _GEN_6300; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6302 = 8'h9e == io_state_in_4 ? 8'h4c : _GEN_6301; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6303 = 8'h9f == io_state_in_4 ? 8'h41 : _GEN_6302; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6304 = 8'ha0 == io_state_in_4 ? 8'h61 : _GEN_6303; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6305 = 8'ha1 == io_state_in_4 ? 8'h6c : _GEN_6304; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6306 = 8'ha2 == io_state_in_4 ? 8'h7b : _GEN_6305; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6307 = 8'ha3 == io_state_in_4 ? 8'h76 : _GEN_6306; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6308 = 8'ha4 == io_state_in_4 ? 8'h55 : _GEN_6307; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6309 = 8'ha5 == io_state_in_4 ? 8'h58 : _GEN_6308; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6310 = 8'ha6 == io_state_in_4 ? 8'h4f : _GEN_6309; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6311 = 8'ha7 == io_state_in_4 ? 8'h42 : _GEN_6310; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6312 = 8'ha8 == io_state_in_4 ? 8'h9 : _GEN_6311; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6313 = 8'ha9 == io_state_in_4 ? 8'h4 : _GEN_6312; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6314 = 8'haa == io_state_in_4 ? 8'h13 : _GEN_6313; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6315 = 8'hab == io_state_in_4 ? 8'h1e : _GEN_6314; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6316 = 8'hac == io_state_in_4 ? 8'h3d : _GEN_6315; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6317 = 8'had == io_state_in_4 ? 8'h30 : _GEN_6316; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6318 = 8'hae == io_state_in_4 ? 8'h27 : _GEN_6317; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6319 = 8'haf == io_state_in_4 ? 8'h2a : _GEN_6318; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6320 = 8'hb0 == io_state_in_4 ? 8'hb1 : _GEN_6319; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6321 = 8'hb1 == io_state_in_4 ? 8'hbc : _GEN_6320; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6322 = 8'hb2 == io_state_in_4 ? 8'hab : _GEN_6321; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6323 = 8'hb3 == io_state_in_4 ? 8'ha6 : _GEN_6322; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6324 = 8'hb4 == io_state_in_4 ? 8'h85 : _GEN_6323; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6325 = 8'hb5 == io_state_in_4 ? 8'h88 : _GEN_6324; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6326 = 8'hb6 == io_state_in_4 ? 8'h9f : _GEN_6325; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6327 = 8'hb7 == io_state_in_4 ? 8'h92 : _GEN_6326; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6328 = 8'hb8 == io_state_in_4 ? 8'hd9 : _GEN_6327; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6329 = 8'hb9 == io_state_in_4 ? 8'hd4 : _GEN_6328; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6330 = 8'hba == io_state_in_4 ? 8'hc3 : _GEN_6329; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6331 = 8'hbb == io_state_in_4 ? 8'hce : _GEN_6330; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6332 = 8'hbc == io_state_in_4 ? 8'hed : _GEN_6331; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6333 = 8'hbd == io_state_in_4 ? 8'he0 : _GEN_6332; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6334 = 8'hbe == io_state_in_4 ? 8'hf7 : _GEN_6333; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6335 = 8'hbf == io_state_in_4 ? 8'hfa : _GEN_6334; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6336 = 8'hc0 == io_state_in_4 ? 8'hb7 : _GEN_6335; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6337 = 8'hc1 == io_state_in_4 ? 8'hba : _GEN_6336; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6338 = 8'hc2 == io_state_in_4 ? 8'had : _GEN_6337; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6339 = 8'hc3 == io_state_in_4 ? 8'ha0 : _GEN_6338; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6340 = 8'hc4 == io_state_in_4 ? 8'h83 : _GEN_6339; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6341 = 8'hc5 == io_state_in_4 ? 8'h8e : _GEN_6340; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6342 = 8'hc6 == io_state_in_4 ? 8'h99 : _GEN_6341; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6343 = 8'hc7 == io_state_in_4 ? 8'h94 : _GEN_6342; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6344 = 8'hc8 == io_state_in_4 ? 8'hdf : _GEN_6343; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6345 = 8'hc9 == io_state_in_4 ? 8'hd2 : _GEN_6344; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6346 = 8'hca == io_state_in_4 ? 8'hc5 : _GEN_6345; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6347 = 8'hcb == io_state_in_4 ? 8'hc8 : _GEN_6346; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6348 = 8'hcc == io_state_in_4 ? 8'heb : _GEN_6347; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6349 = 8'hcd == io_state_in_4 ? 8'he6 : _GEN_6348; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6350 = 8'hce == io_state_in_4 ? 8'hf1 : _GEN_6349; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6351 = 8'hcf == io_state_in_4 ? 8'hfc : _GEN_6350; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6352 = 8'hd0 == io_state_in_4 ? 8'h67 : _GEN_6351; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6353 = 8'hd1 == io_state_in_4 ? 8'h6a : _GEN_6352; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6354 = 8'hd2 == io_state_in_4 ? 8'h7d : _GEN_6353; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6355 = 8'hd3 == io_state_in_4 ? 8'h70 : _GEN_6354; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6356 = 8'hd4 == io_state_in_4 ? 8'h53 : _GEN_6355; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6357 = 8'hd5 == io_state_in_4 ? 8'h5e : _GEN_6356; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6358 = 8'hd6 == io_state_in_4 ? 8'h49 : _GEN_6357; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6359 = 8'hd7 == io_state_in_4 ? 8'h44 : _GEN_6358; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6360 = 8'hd8 == io_state_in_4 ? 8'hf : _GEN_6359; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6361 = 8'hd9 == io_state_in_4 ? 8'h2 : _GEN_6360; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6362 = 8'hda == io_state_in_4 ? 8'h15 : _GEN_6361; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6363 = 8'hdb == io_state_in_4 ? 8'h18 : _GEN_6362; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6364 = 8'hdc == io_state_in_4 ? 8'h3b : _GEN_6363; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6365 = 8'hdd == io_state_in_4 ? 8'h36 : _GEN_6364; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6366 = 8'hde == io_state_in_4 ? 8'h21 : _GEN_6365; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6367 = 8'hdf == io_state_in_4 ? 8'h2c : _GEN_6366; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6368 = 8'he0 == io_state_in_4 ? 8'hc : _GEN_6367; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6369 = 8'he1 == io_state_in_4 ? 8'h1 : _GEN_6368; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6370 = 8'he2 == io_state_in_4 ? 8'h16 : _GEN_6369; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6371 = 8'he3 == io_state_in_4 ? 8'h1b : _GEN_6370; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6372 = 8'he4 == io_state_in_4 ? 8'h38 : _GEN_6371; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6373 = 8'he5 == io_state_in_4 ? 8'h35 : _GEN_6372; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6374 = 8'he6 == io_state_in_4 ? 8'h22 : _GEN_6373; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6375 = 8'he7 == io_state_in_4 ? 8'h2f : _GEN_6374; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6376 = 8'he8 == io_state_in_4 ? 8'h64 : _GEN_6375; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6377 = 8'he9 == io_state_in_4 ? 8'h69 : _GEN_6376; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6378 = 8'hea == io_state_in_4 ? 8'h7e : _GEN_6377; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6379 = 8'heb == io_state_in_4 ? 8'h73 : _GEN_6378; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6380 = 8'hec == io_state_in_4 ? 8'h50 : _GEN_6379; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6381 = 8'hed == io_state_in_4 ? 8'h5d : _GEN_6380; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6382 = 8'hee == io_state_in_4 ? 8'h4a : _GEN_6381; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6383 = 8'hef == io_state_in_4 ? 8'h47 : _GEN_6382; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6384 = 8'hf0 == io_state_in_4 ? 8'hdc : _GEN_6383; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6385 = 8'hf1 == io_state_in_4 ? 8'hd1 : _GEN_6384; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6386 = 8'hf2 == io_state_in_4 ? 8'hc6 : _GEN_6385; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6387 = 8'hf3 == io_state_in_4 ? 8'hcb : _GEN_6386; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6388 = 8'hf4 == io_state_in_4 ? 8'he8 : _GEN_6387; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6389 = 8'hf5 == io_state_in_4 ? 8'he5 : _GEN_6388; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6390 = 8'hf6 == io_state_in_4 ? 8'hf2 : _GEN_6389; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6391 = 8'hf7 == io_state_in_4 ? 8'hff : _GEN_6390; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6392 = 8'hf8 == io_state_in_4 ? 8'hb4 : _GEN_6391; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6393 = 8'hf9 == io_state_in_4 ? 8'hb9 : _GEN_6392; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6394 = 8'hfa == io_state_in_4 ? 8'hae : _GEN_6393; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6395 = 8'hfb == io_state_in_4 ? 8'ha3 : _GEN_6394; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6396 = 8'hfc == io_state_in_4 ? 8'h80 : _GEN_6395; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6397 = 8'hfd == io_state_in_4 ? 8'h8d : _GEN_6396; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6398 = 8'hfe == io_state_in_4 ? 8'h9a : _GEN_6397; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6399 = 8'hff == io_state_in_4 ? 8'h97 : _GEN_6398; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6401 = 8'h1 == io_state_in_5 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6402 = 8'h2 == io_state_in_5 ? 8'h12 : _GEN_6401; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6403 = 8'h3 == io_state_in_5 ? 8'h1b : _GEN_6402; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6404 = 8'h4 == io_state_in_5 ? 8'h24 : _GEN_6403; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6405 = 8'h5 == io_state_in_5 ? 8'h2d : _GEN_6404; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6406 = 8'h6 == io_state_in_5 ? 8'h36 : _GEN_6405; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6407 = 8'h7 == io_state_in_5 ? 8'h3f : _GEN_6406; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6408 = 8'h8 == io_state_in_5 ? 8'h48 : _GEN_6407; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6409 = 8'h9 == io_state_in_5 ? 8'h41 : _GEN_6408; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6410 = 8'ha == io_state_in_5 ? 8'h5a : _GEN_6409; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6411 = 8'hb == io_state_in_5 ? 8'h53 : _GEN_6410; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6412 = 8'hc == io_state_in_5 ? 8'h6c : _GEN_6411; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6413 = 8'hd == io_state_in_5 ? 8'h65 : _GEN_6412; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6414 = 8'he == io_state_in_5 ? 8'h7e : _GEN_6413; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6415 = 8'hf == io_state_in_5 ? 8'h77 : _GEN_6414; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6416 = 8'h10 == io_state_in_5 ? 8'h90 : _GEN_6415; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6417 = 8'h11 == io_state_in_5 ? 8'h99 : _GEN_6416; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6418 = 8'h12 == io_state_in_5 ? 8'h82 : _GEN_6417; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6419 = 8'h13 == io_state_in_5 ? 8'h8b : _GEN_6418; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6420 = 8'h14 == io_state_in_5 ? 8'hb4 : _GEN_6419; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6421 = 8'h15 == io_state_in_5 ? 8'hbd : _GEN_6420; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6422 = 8'h16 == io_state_in_5 ? 8'ha6 : _GEN_6421; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6423 = 8'h17 == io_state_in_5 ? 8'haf : _GEN_6422; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6424 = 8'h18 == io_state_in_5 ? 8'hd8 : _GEN_6423; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6425 = 8'h19 == io_state_in_5 ? 8'hd1 : _GEN_6424; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6426 = 8'h1a == io_state_in_5 ? 8'hca : _GEN_6425; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6427 = 8'h1b == io_state_in_5 ? 8'hc3 : _GEN_6426; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6428 = 8'h1c == io_state_in_5 ? 8'hfc : _GEN_6427; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6429 = 8'h1d == io_state_in_5 ? 8'hf5 : _GEN_6428; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6430 = 8'h1e == io_state_in_5 ? 8'hee : _GEN_6429; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6431 = 8'h1f == io_state_in_5 ? 8'he7 : _GEN_6430; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6432 = 8'h20 == io_state_in_5 ? 8'h3b : _GEN_6431; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6433 = 8'h21 == io_state_in_5 ? 8'h32 : _GEN_6432; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6434 = 8'h22 == io_state_in_5 ? 8'h29 : _GEN_6433; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6435 = 8'h23 == io_state_in_5 ? 8'h20 : _GEN_6434; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6436 = 8'h24 == io_state_in_5 ? 8'h1f : _GEN_6435; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6437 = 8'h25 == io_state_in_5 ? 8'h16 : _GEN_6436; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6438 = 8'h26 == io_state_in_5 ? 8'hd : _GEN_6437; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6439 = 8'h27 == io_state_in_5 ? 8'h4 : _GEN_6438; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6440 = 8'h28 == io_state_in_5 ? 8'h73 : _GEN_6439; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6441 = 8'h29 == io_state_in_5 ? 8'h7a : _GEN_6440; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6442 = 8'h2a == io_state_in_5 ? 8'h61 : _GEN_6441; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6443 = 8'h2b == io_state_in_5 ? 8'h68 : _GEN_6442; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6444 = 8'h2c == io_state_in_5 ? 8'h57 : _GEN_6443; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6445 = 8'h2d == io_state_in_5 ? 8'h5e : _GEN_6444; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6446 = 8'h2e == io_state_in_5 ? 8'h45 : _GEN_6445; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6447 = 8'h2f == io_state_in_5 ? 8'h4c : _GEN_6446; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6448 = 8'h30 == io_state_in_5 ? 8'hab : _GEN_6447; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6449 = 8'h31 == io_state_in_5 ? 8'ha2 : _GEN_6448; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6450 = 8'h32 == io_state_in_5 ? 8'hb9 : _GEN_6449; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6451 = 8'h33 == io_state_in_5 ? 8'hb0 : _GEN_6450; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6452 = 8'h34 == io_state_in_5 ? 8'h8f : _GEN_6451; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6453 = 8'h35 == io_state_in_5 ? 8'h86 : _GEN_6452; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6454 = 8'h36 == io_state_in_5 ? 8'h9d : _GEN_6453; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6455 = 8'h37 == io_state_in_5 ? 8'h94 : _GEN_6454; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6456 = 8'h38 == io_state_in_5 ? 8'he3 : _GEN_6455; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6457 = 8'h39 == io_state_in_5 ? 8'hea : _GEN_6456; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6458 = 8'h3a == io_state_in_5 ? 8'hf1 : _GEN_6457; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6459 = 8'h3b == io_state_in_5 ? 8'hf8 : _GEN_6458; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6460 = 8'h3c == io_state_in_5 ? 8'hc7 : _GEN_6459; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6461 = 8'h3d == io_state_in_5 ? 8'hce : _GEN_6460; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6462 = 8'h3e == io_state_in_5 ? 8'hd5 : _GEN_6461; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6463 = 8'h3f == io_state_in_5 ? 8'hdc : _GEN_6462; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6464 = 8'h40 == io_state_in_5 ? 8'h76 : _GEN_6463; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6465 = 8'h41 == io_state_in_5 ? 8'h7f : _GEN_6464; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6466 = 8'h42 == io_state_in_5 ? 8'h64 : _GEN_6465; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6467 = 8'h43 == io_state_in_5 ? 8'h6d : _GEN_6466; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6468 = 8'h44 == io_state_in_5 ? 8'h52 : _GEN_6467; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6469 = 8'h45 == io_state_in_5 ? 8'h5b : _GEN_6468; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6470 = 8'h46 == io_state_in_5 ? 8'h40 : _GEN_6469; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6471 = 8'h47 == io_state_in_5 ? 8'h49 : _GEN_6470; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6472 = 8'h48 == io_state_in_5 ? 8'h3e : _GEN_6471; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6473 = 8'h49 == io_state_in_5 ? 8'h37 : _GEN_6472; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6474 = 8'h4a == io_state_in_5 ? 8'h2c : _GEN_6473; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6475 = 8'h4b == io_state_in_5 ? 8'h25 : _GEN_6474; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6476 = 8'h4c == io_state_in_5 ? 8'h1a : _GEN_6475; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6477 = 8'h4d == io_state_in_5 ? 8'h13 : _GEN_6476; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6478 = 8'h4e == io_state_in_5 ? 8'h8 : _GEN_6477; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6479 = 8'h4f == io_state_in_5 ? 8'h1 : _GEN_6478; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6480 = 8'h50 == io_state_in_5 ? 8'he6 : _GEN_6479; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6481 = 8'h51 == io_state_in_5 ? 8'hef : _GEN_6480; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6482 = 8'h52 == io_state_in_5 ? 8'hf4 : _GEN_6481; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6483 = 8'h53 == io_state_in_5 ? 8'hfd : _GEN_6482; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6484 = 8'h54 == io_state_in_5 ? 8'hc2 : _GEN_6483; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6485 = 8'h55 == io_state_in_5 ? 8'hcb : _GEN_6484; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6486 = 8'h56 == io_state_in_5 ? 8'hd0 : _GEN_6485; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6487 = 8'h57 == io_state_in_5 ? 8'hd9 : _GEN_6486; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6488 = 8'h58 == io_state_in_5 ? 8'hae : _GEN_6487; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6489 = 8'h59 == io_state_in_5 ? 8'ha7 : _GEN_6488; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6490 = 8'h5a == io_state_in_5 ? 8'hbc : _GEN_6489; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6491 = 8'h5b == io_state_in_5 ? 8'hb5 : _GEN_6490; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6492 = 8'h5c == io_state_in_5 ? 8'h8a : _GEN_6491; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6493 = 8'h5d == io_state_in_5 ? 8'h83 : _GEN_6492; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6494 = 8'h5e == io_state_in_5 ? 8'h98 : _GEN_6493; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6495 = 8'h5f == io_state_in_5 ? 8'h91 : _GEN_6494; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6496 = 8'h60 == io_state_in_5 ? 8'h4d : _GEN_6495; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6497 = 8'h61 == io_state_in_5 ? 8'h44 : _GEN_6496; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6498 = 8'h62 == io_state_in_5 ? 8'h5f : _GEN_6497; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6499 = 8'h63 == io_state_in_5 ? 8'h56 : _GEN_6498; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6500 = 8'h64 == io_state_in_5 ? 8'h69 : _GEN_6499; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6501 = 8'h65 == io_state_in_5 ? 8'h60 : _GEN_6500; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6502 = 8'h66 == io_state_in_5 ? 8'h7b : _GEN_6501; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6503 = 8'h67 == io_state_in_5 ? 8'h72 : _GEN_6502; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6504 = 8'h68 == io_state_in_5 ? 8'h5 : _GEN_6503; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6505 = 8'h69 == io_state_in_5 ? 8'hc : _GEN_6504; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6506 = 8'h6a == io_state_in_5 ? 8'h17 : _GEN_6505; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6507 = 8'h6b == io_state_in_5 ? 8'h1e : _GEN_6506; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6508 = 8'h6c == io_state_in_5 ? 8'h21 : _GEN_6507; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6509 = 8'h6d == io_state_in_5 ? 8'h28 : _GEN_6508; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6510 = 8'h6e == io_state_in_5 ? 8'h33 : _GEN_6509; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6511 = 8'h6f == io_state_in_5 ? 8'h3a : _GEN_6510; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6512 = 8'h70 == io_state_in_5 ? 8'hdd : _GEN_6511; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6513 = 8'h71 == io_state_in_5 ? 8'hd4 : _GEN_6512; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6514 = 8'h72 == io_state_in_5 ? 8'hcf : _GEN_6513; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6515 = 8'h73 == io_state_in_5 ? 8'hc6 : _GEN_6514; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6516 = 8'h74 == io_state_in_5 ? 8'hf9 : _GEN_6515; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6517 = 8'h75 == io_state_in_5 ? 8'hf0 : _GEN_6516; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6518 = 8'h76 == io_state_in_5 ? 8'heb : _GEN_6517; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6519 = 8'h77 == io_state_in_5 ? 8'he2 : _GEN_6518; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6520 = 8'h78 == io_state_in_5 ? 8'h95 : _GEN_6519; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6521 = 8'h79 == io_state_in_5 ? 8'h9c : _GEN_6520; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6522 = 8'h7a == io_state_in_5 ? 8'h87 : _GEN_6521; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6523 = 8'h7b == io_state_in_5 ? 8'h8e : _GEN_6522; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6524 = 8'h7c == io_state_in_5 ? 8'hb1 : _GEN_6523; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6525 = 8'h7d == io_state_in_5 ? 8'hb8 : _GEN_6524; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6526 = 8'h7e == io_state_in_5 ? 8'ha3 : _GEN_6525; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6527 = 8'h7f == io_state_in_5 ? 8'haa : _GEN_6526; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6528 = 8'h80 == io_state_in_5 ? 8'hec : _GEN_6527; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6529 = 8'h81 == io_state_in_5 ? 8'he5 : _GEN_6528; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6530 = 8'h82 == io_state_in_5 ? 8'hfe : _GEN_6529; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6531 = 8'h83 == io_state_in_5 ? 8'hf7 : _GEN_6530; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6532 = 8'h84 == io_state_in_5 ? 8'hc8 : _GEN_6531; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6533 = 8'h85 == io_state_in_5 ? 8'hc1 : _GEN_6532; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6534 = 8'h86 == io_state_in_5 ? 8'hda : _GEN_6533; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6535 = 8'h87 == io_state_in_5 ? 8'hd3 : _GEN_6534; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6536 = 8'h88 == io_state_in_5 ? 8'ha4 : _GEN_6535; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6537 = 8'h89 == io_state_in_5 ? 8'had : _GEN_6536; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6538 = 8'h8a == io_state_in_5 ? 8'hb6 : _GEN_6537; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6539 = 8'h8b == io_state_in_5 ? 8'hbf : _GEN_6538; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6540 = 8'h8c == io_state_in_5 ? 8'h80 : _GEN_6539; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6541 = 8'h8d == io_state_in_5 ? 8'h89 : _GEN_6540; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6542 = 8'h8e == io_state_in_5 ? 8'h92 : _GEN_6541; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6543 = 8'h8f == io_state_in_5 ? 8'h9b : _GEN_6542; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6544 = 8'h90 == io_state_in_5 ? 8'h7c : _GEN_6543; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6545 = 8'h91 == io_state_in_5 ? 8'h75 : _GEN_6544; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6546 = 8'h92 == io_state_in_5 ? 8'h6e : _GEN_6545; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6547 = 8'h93 == io_state_in_5 ? 8'h67 : _GEN_6546; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6548 = 8'h94 == io_state_in_5 ? 8'h58 : _GEN_6547; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6549 = 8'h95 == io_state_in_5 ? 8'h51 : _GEN_6548; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6550 = 8'h96 == io_state_in_5 ? 8'h4a : _GEN_6549; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6551 = 8'h97 == io_state_in_5 ? 8'h43 : _GEN_6550; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6552 = 8'h98 == io_state_in_5 ? 8'h34 : _GEN_6551; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6553 = 8'h99 == io_state_in_5 ? 8'h3d : _GEN_6552; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6554 = 8'h9a == io_state_in_5 ? 8'h26 : _GEN_6553; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6555 = 8'h9b == io_state_in_5 ? 8'h2f : _GEN_6554; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6556 = 8'h9c == io_state_in_5 ? 8'h10 : _GEN_6555; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6557 = 8'h9d == io_state_in_5 ? 8'h19 : _GEN_6556; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6558 = 8'h9e == io_state_in_5 ? 8'h2 : _GEN_6557; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6559 = 8'h9f == io_state_in_5 ? 8'hb : _GEN_6558; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6560 = 8'ha0 == io_state_in_5 ? 8'hd7 : _GEN_6559; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6561 = 8'ha1 == io_state_in_5 ? 8'hde : _GEN_6560; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6562 = 8'ha2 == io_state_in_5 ? 8'hc5 : _GEN_6561; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6563 = 8'ha3 == io_state_in_5 ? 8'hcc : _GEN_6562; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6564 = 8'ha4 == io_state_in_5 ? 8'hf3 : _GEN_6563; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6565 = 8'ha5 == io_state_in_5 ? 8'hfa : _GEN_6564; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6566 = 8'ha6 == io_state_in_5 ? 8'he1 : _GEN_6565; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6567 = 8'ha7 == io_state_in_5 ? 8'he8 : _GEN_6566; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6568 = 8'ha8 == io_state_in_5 ? 8'h9f : _GEN_6567; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6569 = 8'ha9 == io_state_in_5 ? 8'h96 : _GEN_6568; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6570 = 8'haa == io_state_in_5 ? 8'h8d : _GEN_6569; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6571 = 8'hab == io_state_in_5 ? 8'h84 : _GEN_6570; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6572 = 8'hac == io_state_in_5 ? 8'hbb : _GEN_6571; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6573 = 8'had == io_state_in_5 ? 8'hb2 : _GEN_6572; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6574 = 8'hae == io_state_in_5 ? 8'ha9 : _GEN_6573; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6575 = 8'haf == io_state_in_5 ? 8'ha0 : _GEN_6574; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6576 = 8'hb0 == io_state_in_5 ? 8'h47 : _GEN_6575; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6577 = 8'hb1 == io_state_in_5 ? 8'h4e : _GEN_6576; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6578 = 8'hb2 == io_state_in_5 ? 8'h55 : _GEN_6577; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6579 = 8'hb3 == io_state_in_5 ? 8'h5c : _GEN_6578; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6580 = 8'hb4 == io_state_in_5 ? 8'h63 : _GEN_6579; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6581 = 8'hb5 == io_state_in_5 ? 8'h6a : _GEN_6580; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6582 = 8'hb6 == io_state_in_5 ? 8'h71 : _GEN_6581; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6583 = 8'hb7 == io_state_in_5 ? 8'h78 : _GEN_6582; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6584 = 8'hb8 == io_state_in_5 ? 8'hf : _GEN_6583; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6585 = 8'hb9 == io_state_in_5 ? 8'h6 : _GEN_6584; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6586 = 8'hba == io_state_in_5 ? 8'h1d : _GEN_6585; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6587 = 8'hbb == io_state_in_5 ? 8'h14 : _GEN_6586; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6588 = 8'hbc == io_state_in_5 ? 8'h2b : _GEN_6587; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6589 = 8'hbd == io_state_in_5 ? 8'h22 : _GEN_6588; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6590 = 8'hbe == io_state_in_5 ? 8'h39 : _GEN_6589; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6591 = 8'hbf == io_state_in_5 ? 8'h30 : _GEN_6590; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6592 = 8'hc0 == io_state_in_5 ? 8'h9a : _GEN_6591; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6593 = 8'hc1 == io_state_in_5 ? 8'h93 : _GEN_6592; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6594 = 8'hc2 == io_state_in_5 ? 8'h88 : _GEN_6593; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6595 = 8'hc3 == io_state_in_5 ? 8'h81 : _GEN_6594; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6596 = 8'hc4 == io_state_in_5 ? 8'hbe : _GEN_6595; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6597 = 8'hc5 == io_state_in_5 ? 8'hb7 : _GEN_6596; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6598 = 8'hc6 == io_state_in_5 ? 8'hac : _GEN_6597; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6599 = 8'hc7 == io_state_in_5 ? 8'ha5 : _GEN_6598; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6600 = 8'hc8 == io_state_in_5 ? 8'hd2 : _GEN_6599; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6601 = 8'hc9 == io_state_in_5 ? 8'hdb : _GEN_6600; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6602 = 8'hca == io_state_in_5 ? 8'hc0 : _GEN_6601; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6603 = 8'hcb == io_state_in_5 ? 8'hc9 : _GEN_6602; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6604 = 8'hcc == io_state_in_5 ? 8'hf6 : _GEN_6603; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6605 = 8'hcd == io_state_in_5 ? 8'hff : _GEN_6604; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6606 = 8'hce == io_state_in_5 ? 8'he4 : _GEN_6605; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6607 = 8'hcf == io_state_in_5 ? 8'hed : _GEN_6606; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6608 = 8'hd0 == io_state_in_5 ? 8'ha : _GEN_6607; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6609 = 8'hd1 == io_state_in_5 ? 8'h3 : _GEN_6608; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6610 = 8'hd2 == io_state_in_5 ? 8'h18 : _GEN_6609; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6611 = 8'hd3 == io_state_in_5 ? 8'h11 : _GEN_6610; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6612 = 8'hd4 == io_state_in_5 ? 8'h2e : _GEN_6611; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6613 = 8'hd5 == io_state_in_5 ? 8'h27 : _GEN_6612; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6614 = 8'hd6 == io_state_in_5 ? 8'h3c : _GEN_6613; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6615 = 8'hd7 == io_state_in_5 ? 8'h35 : _GEN_6614; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6616 = 8'hd8 == io_state_in_5 ? 8'h42 : _GEN_6615; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6617 = 8'hd9 == io_state_in_5 ? 8'h4b : _GEN_6616; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6618 = 8'hda == io_state_in_5 ? 8'h50 : _GEN_6617; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6619 = 8'hdb == io_state_in_5 ? 8'h59 : _GEN_6618; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6620 = 8'hdc == io_state_in_5 ? 8'h66 : _GEN_6619; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6621 = 8'hdd == io_state_in_5 ? 8'h6f : _GEN_6620; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6622 = 8'hde == io_state_in_5 ? 8'h74 : _GEN_6621; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6623 = 8'hdf == io_state_in_5 ? 8'h7d : _GEN_6622; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6624 = 8'he0 == io_state_in_5 ? 8'ha1 : _GEN_6623; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6625 = 8'he1 == io_state_in_5 ? 8'ha8 : _GEN_6624; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6626 = 8'he2 == io_state_in_5 ? 8'hb3 : _GEN_6625; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6627 = 8'he3 == io_state_in_5 ? 8'hba : _GEN_6626; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6628 = 8'he4 == io_state_in_5 ? 8'h85 : _GEN_6627; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6629 = 8'he5 == io_state_in_5 ? 8'h8c : _GEN_6628; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6630 = 8'he6 == io_state_in_5 ? 8'h97 : _GEN_6629; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6631 = 8'he7 == io_state_in_5 ? 8'h9e : _GEN_6630; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6632 = 8'he8 == io_state_in_5 ? 8'he9 : _GEN_6631; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6633 = 8'he9 == io_state_in_5 ? 8'he0 : _GEN_6632; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6634 = 8'hea == io_state_in_5 ? 8'hfb : _GEN_6633; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6635 = 8'heb == io_state_in_5 ? 8'hf2 : _GEN_6634; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6636 = 8'hec == io_state_in_5 ? 8'hcd : _GEN_6635; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6637 = 8'hed == io_state_in_5 ? 8'hc4 : _GEN_6636; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6638 = 8'hee == io_state_in_5 ? 8'hdf : _GEN_6637; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6639 = 8'hef == io_state_in_5 ? 8'hd6 : _GEN_6638; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6640 = 8'hf0 == io_state_in_5 ? 8'h31 : _GEN_6639; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6641 = 8'hf1 == io_state_in_5 ? 8'h38 : _GEN_6640; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6642 = 8'hf2 == io_state_in_5 ? 8'h23 : _GEN_6641; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6643 = 8'hf3 == io_state_in_5 ? 8'h2a : _GEN_6642; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6644 = 8'hf4 == io_state_in_5 ? 8'h15 : _GEN_6643; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6645 = 8'hf5 == io_state_in_5 ? 8'h1c : _GEN_6644; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6646 = 8'hf6 == io_state_in_5 ? 8'h7 : _GEN_6645; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6647 = 8'hf7 == io_state_in_5 ? 8'he : _GEN_6646; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6648 = 8'hf8 == io_state_in_5 ? 8'h79 : _GEN_6647; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6649 = 8'hf9 == io_state_in_5 ? 8'h70 : _GEN_6648; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6650 = 8'hfa == io_state_in_5 ? 8'h6b : _GEN_6649; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6651 = 8'hfb == io_state_in_5 ? 8'h62 : _GEN_6650; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6652 = 8'hfc == io_state_in_5 ? 8'h5d : _GEN_6651; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6653 = 8'hfd == io_state_in_5 ? 8'h54 : _GEN_6652; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6654 = 8'hfe == io_state_in_5 ? 8'h4f : _GEN_6653; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_6655 = 8'hff == io_state_in_5 ? 8'h46 : _GEN_6654; // @[InvMixColumns.scala 133:{41,41}]
  wire [7:0] _tmp_state_6_T = _GEN_6399 ^ _GEN_6655; // @[InvMixColumns.scala 133:41]
  wire [7:0] _GEN_6657 = 8'h1 == io_state_in_6 ? 8'he : 8'h0; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6658 = 8'h2 == io_state_in_6 ? 8'h1c : _GEN_6657; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6659 = 8'h3 == io_state_in_6 ? 8'h12 : _GEN_6658; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6660 = 8'h4 == io_state_in_6 ? 8'h38 : _GEN_6659; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6661 = 8'h5 == io_state_in_6 ? 8'h36 : _GEN_6660; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6662 = 8'h6 == io_state_in_6 ? 8'h24 : _GEN_6661; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6663 = 8'h7 == io_state_in_6 ? 8'h2a : _GEN_6662; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6664 = 8'h8 == io_state_in_6 ? 8'h70 : _GEN_6663; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6665 = 8'h9 == io_state_in_6 ? 8'h7e : _GEN_6664; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6666 = 8'ha == io_state_in_6 ? 8'h6c : _GEN_6665; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6667 = 8'hb == io_state_in_6 ? 8'h62 : _GEN_6666; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6668 = 8'hc == io_state_in_6 ? 8'h48 : _GEN_6667; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6669 = 8'hd == io_state_in_6 ? 8'h46 : _GEN_6668; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6670 = 8'he == io_state_in_6 ? 8'h54 : _GEN_6669; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6671 = 8'hf == io_state_in_6 ? 8'h5a : _GEN_6670; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6672 = 8'h10 == io_state_in_6 ? 8'he0 : _GEN_6671; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6673 = 8'h11 == io_state_in_6 ? 8'hee : _GEN_6672; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6674 = 8'h12 == io_state_in_6 ? 8'hfc : _GEN_6673; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6675 = 8'h13 == io_state_in_6 ? 8'hf2 : _GEN_6674; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6676 = 8'h14 == io_state_in_6 ? 8'hd8 : _GEN_6675; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6677 = 8'h15 == io_state_in_6 ? 8'hd6 : _GEN_6676; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6678 = 8'h16 == io_state_in_6 ? 8'hc4 : _GEN_6677; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6679 = 8'h17 == io_state_in_6 ? 8'hca : _GEN_6678; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6680 = 8'h18 == io_state_in_6 ? 8'h90 : _GEN_6679; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6681 = 8'h19 == io_state_in_6 ? 8'h9e : _GEN_6680; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6682 = 8'h1a == io_state_in_6 ? 8'h8c : _GEN_6681; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6683 = 8'h1b == io_state_in_6 ? 8'h82 : _GEN_6682; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6684 = 8'h1c == io_state_in_6 ? 8'ha8 : _GEN_6683; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6685 = 8'h1d == io_state_in_6 ? 8'ha6 : _GEN_6684; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6686 = 8'h1e == io_state_in_6 ? 8'hb4 : _GEN_6685; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6687 = 8'h1f == io_state_in_6 ? 8'hba : _GEN_6686; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6688 = 8'h20 == io_state_in_6 ? 8'hdb : _GEN_6687; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6689 = 8'h21 == io_state_in_6 ? 8'hd5 : _GEN_6688; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6690 = 8'h22 == io_state_in_6 ? 8'hc7 : _GEN_6689; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6691 = 8'h23 == io_state_in_6 ? 8'hc9 : _GEN_6690; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6692 = 8'h24 == io_state_in_6 ? 8'he3 : _GEN_6691; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6693 = 8'h25 == io_state_in_6 ? 8'hed : _GEN_6692; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6694 = 8'h26 == io_state_in_6 ? 8'hff : _GEN_6693; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6695 = 8'h27 == io_state_in_6 ? 8'hf1 : _GEN_6694; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6696 = 8'h28 == io_state_in_6 ? 8'hab : _GEN_6695; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6697 = 8'h29 == io_state_in_6 ? 8'ha5 : _GEN_6696; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6698 = 8'h2a == io_state_in_6 ? 8'hb7 : _GEN_6697; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6699 = 8'h2b == io_state_in_6 ? 8'hb9 : _GEN_6698; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6700 = 8'h2c == io_state_in_6 ? 8'h93 : _GEN_6699; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6701 = 8'h2d == io_state_in_6 ? 8'h9d : _GEN_6700; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6702 = 8'h2e == io_state_in_6 ? 8'h8f : _GEN_6701; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6703 = 8'h2f == io_state_in_6 ? 8'h81 : _GEN_6702; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6704 = 8'h30 == io_state_in_6 ? 8'h3b : _GEN_6703; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6705 = 8'h31 == io_state_in_6 ? 8'h35 : _GEN_6704; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6706 = 8'h32 == io_state_in_6 ? 8'h27 : _GEN_6705; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6707 = 8'h33 == io_state_in_6 ? 8'h29 : _GEN_6706; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6708 = 8'h34 == io_state_in_6 ? 8'h3 : _GEN_6707; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6709 = 8'h35 == io_state_in_6 ? 8'hd : _GEN_6708; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6710 = 8'h36 == io_state_in_6 ? 8'h1f : _GEN_6709; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6711 = 8'h37 == io_state_in_6 ? 8'h11 : _GEN_6710; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6712 = 8'h38 == io_state_in_6 ? 8'h4b : _GEN_6711; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6713 = 8'h39 == io_state_in_6 ? 8'h45 : _GEN_6712; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6714 = 8'h3a == io_state_in_6 ? 8'h57 : _GEN_6713; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6715 = 8'h3b == io_state_in_6 ? 8'h59 : _GEN_6714; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6716 = 8'h3c == io_state_in_6 ? 8'h73 : _GEN_6715; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6717 = 8'h3d == io_state_in_6 ? 8'h7d : _GEN_6716; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6718 = 8'h3e == io_state_in_6 ? 8'h6f : _GEN_6717; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6719 = 8'h3f == io_state_in_6 ? 8'h61 : _GEN_6718; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6720 = 8'h40 == io_state_in_6 ? 8'had : _GEN_6719; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6721 = 8'h41 == io_state_in_6 ? 8'ha3 : _GEN_6720; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6722 = 8'h42 == io_state_in_6 ? 8'hb1 : _GEN_6721; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6723 = 8'h43 == io_state_in_6 ? 8'hbf : _GEN_6722; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6724 = 8'h44 == io_state_in_6 ? 8'h95 : _GEN_6723; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6725 = 8'h45 == io_state_in_6 ? 8'h9b : _GEN_6724; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6726 = 8'h46 == io_state_in_6 ? 8'h89 : _GEN_6725; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6727 = 8'h47 == io_state_in_6 ? 8'h87 : _GEN_6726; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6728 = 8'h48 == io_state_in_6 ? 8'hdd : _GEN_6727; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6729 = 8'h49 == io_state_in_6 ? 8'hd3 : _GEN_6728; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6730 = 8'h4a == io_state_in_6 ? 8'hc1 : _GEN_6729; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6731 = 8'h4b == io_state_in_6 ? 8'hcf : _GEN_6730; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6732 = 8'h4c == io_state_in_6 ? 8'he5 : _GEN_6731; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6733 = 8'h4d == io_state_in_6 ? 8'heb : _GEN_6732; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6734 = 8'h4e == io_state_in_6 ? 8'hf9 : _GEN_6733; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6735 = 8'h4f == io_state_in_6 ? 8'hf7 : _GEN_6734; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6736 = 8'h50 == io_state_in_6 ? 8'h4d : _GEN_6735; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6737 = 8'h51 == io_state_in_6 ? 8'h43 : _GEN_6736; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6738 = 8'h52 == io_state_in_6 ? 8'h51 : _GEN_6737; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6739 = 8'h53 == io_state_in_6 ? 8'h5f : _GEN_6738; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6740 = 8'h54 == io_state_in_6 ? 8'h75 : _GEN_6739; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6741 = 8'h55 == io_state_in_6 ? 8'h7b : _GEN_6740; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6742 = 8'h56 == io_state_in_6 ? 8'h69 : _GEN_6741; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6743 = 8'h57 == io_state_in_6 ? 8'h67 : _GEN_6742; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6744 = 8'h58 == io_state_in_6 ? 8'h3d : _GEN_6743; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6745 = 8'h59 == io_state_in_6 ? 8'h33 : _GEN_6744; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6746 = 8'h5a == io_state_in_6 ? 8'h21 : _GEN_6745; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6747 = 8'h5b == io_state_in_6 ? 8'h2f : _GEN_6746; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6748 = 8'h5c == io_state_in_6 ? 8'h5 : _GEN_6747; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6749 = 8'h5d == io_state_in_6 ? 8'hb : _GEN_6748; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6750 = 8'h5e == io_state_in_6 ? 8'h19 : _GEN_6749; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6751 = 8'h5f == io_state_in_6 ? 8'h17 : _GEN_6750; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6752 = 8'h60 == io_state_in_6 ? 8'h76 : _GEN_6751; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6753 = 8'h61 == io_state_in_6 ? 8'h78 : _GEN_6752; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6754 = 8'h62 == io_state_in_6 ? 8'h6a : _GEN_6753; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6755 = 8'h63 == io_state_in_6 ? 8'h64 : _GEN_6754; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6756 = 8'h64 == io_state_in_6 ? 8'h4e : _GEN_6755; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6757 = 8'h65 == io_state_in_6 ? 8'h40 : _GEN_6756; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6758 = 8'h66 == io_state_in_6 ? 8'h52 : _GEN_6757; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6759 = 8'h67 == io_state_in_6 ? 8'h5c : _GEN_6758; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6760 = 8'h68 == io_state_in_6 ? 8'h6 : _GEN_6759; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6761 = 8'h69 == io_state_in_6 ? 8'h8 : _GEN_6760; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6762 = 8'h6a == io_state_in_6 ? 8'h1a : _GEN_6761; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6763 = 8'h6b == io_state_in_6 ? 8'h14 : _GEN_6762; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6764 = 8'h6c == io_state_in_6 ? 8'h3e : _GEN_6763; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6765 = 8'h6d == io_state_in_6 ? 8'h30 : _GEN_6764; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6766 = 8'h6e == io_state_in_6 ? 8'h22 : _GEN_6765; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6767 = 8'h6f == io_state_in_6 ? 8'h2c : _GEN_6766; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6768 = 8'h70 == io_state_in_6 ? 8'h96 : _GEN_6767; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6769 = 8'h71 == io_state_in_6 ? 8'h98 : _GEN_6768; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6770 = 8'h72 == io_state_in_6 ? 8'h8a : _GEN_6769; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6771 = 8'h73 == io_state_in_6 ? 8'h84 : _GEN_6770; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6772 = 8'h74 == io_state_in_6 ? 8'hae : _GEN_6771; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6773 = 8'h75 == io_state_in_6 ? 8'ha0 : _GEN_6772; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6774 = 8'h76 == io_state_in_6 ? 8'hb2 : _GEN_6773; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6775 = 8'h77 == io_state_in_6 ? 8'hbc : _GEN_6774; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6776 = 8'h78 == io_state_in_6 ? 8'he6 : _GEN_6775; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6777 = 8'h79 == io_state_in_6 ? 8'he8 : _GEN_6776; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6778 = 8'h7a == io_state_in_6 ? 8'hfa : _GEN_6777; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6779 = 8'h7b == io_state_in_6 ? 8'hf4 : _GEN_6778; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6780 = 8'h7c == io_state_in_6 ? 8'hde : _GEN_6779; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6781 = 8'h7d == io_state_in_6 ? 8'hd0 : _GEN_6780; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6782 = 8'h7e == io_state_in_6 ? 8'hc2 : _GEN_6781; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6783 = 8'h7f == io_state_in_6 ? 8'hcc : _GEN_6782; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6784 = 8'h80 == io_state_in_6 ? 8'h41 : _GEN_6783; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6785 = 8'h81 == io_state_in_6 ? 8'h4f : _GEN_6784; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6786 = 8'h82 == io_state_in_6 ? 8'h5d : _GEN_6785; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6787 = 8'h83 == io_state_in_6 ? 8'h53 : _GEN_6786; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6788 = 8'h84 == io_state_in_6 ? 8'h79 : _GEN_6787; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6789 = 8'h85 == io_state_in_6 ? 8'h77 : _GEN_6788; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6790 = 8'h86 == io_state_in_6 ? 8'h65 : _GEN_6789; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6791 = 8'h87 == io_state_in_6 ? 8'h6b : _GEN_6790; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6792 = 8'h88 == io_state_in_6 ? 8'h31 : _GEN_6791; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6793 = 8'h89 == io_state_in_6 ? 8'h3f : _GEN_6792; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6794 = 8'h8a == io_state_in_6 ? 8'h2d : _GEN_6793; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6795 = 8'h8b == io_state_in_6 ? 8'h23 : _GEN_6794; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6796 = 8'h8c == io_state_in_6 ? 8'h9 : _GEN_6795; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6797 = 8'h8d == io_state_in_6 ? 8'h7 : _GEN_6796; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6798 = 8'h8e == io_state_in_6 ? 8'h15 : _GEN_6797; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6799 = 8'h8f == io_state_in_6 ? 8'h1b : _GEN_6798; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6800 = 8'h90 == io_state_in_6 ? 8'ha1 : _GEN_6799; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6801 = 8'h91 == io_state_in_6 ? 8'haf : _GEN_6800; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6802 = 8'h92 == io_state_in_6 ? 8'hbd : _GEN_6801; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6803 = 8'h93 == io_state_in_6 ? 8'hb3 : _GEN_6802; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6804 = 8'h94 == io_state_in_6 ? 8'h99 : _GEN_6803; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6805 = 8'h95 == io_state_in_6 ? 8'h97 : _GEN_6804; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6806 = 8'h96 == io_state_in_6 ? 8'h85 : _GEN_6805; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6807 = 8'h97 == io_state_in_6 ? 8'h8b : _GEN_6806; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6808 = 8'h98 == io_state_in_6 ? 8'hd1 : _GEN_6807; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6809 = 8'h99 == io_state_in_6 ? 8'hdf : _GEN_6808; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6810 = 8'h9a == io_state_in_6 ? 8'hcd : _GEN_6809; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6811 = 8'h9b == io_state_in_6 ? 8'hc3 : _GEN_6810; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6812 = 8'h9c == io_state_in_6 ? 8'he9 : _GEN_6811; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6813 = 8'h9d == io_state_in_6 ? 8'he7 : _GEN_6812; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6814 = 8'h9e == io_state_in_6 ? 8'hf5 : _GEN_6813; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6815 = 8'h9f == io_state_in_6 ? 8'hfb : _GEN_6814; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6816 = 8'ha0 == io_state_in_6 ? 8'h9a : _GEN_6815; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6817 = 8'ha1 == io_state_in_6 ? 8'h94 : _GEN_6816; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6818 = 8'ha2 == io_state_in_6 ? 8'h86 : _GEN_6817; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6819 = 8'ha3 == io_state_in_6 ? 8'h88 : _GEN_6818; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6820 = 8'ha4 == io_state_in_6 ? 8'ha2 : _GEN_6819; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6821 = 8'ha5 == io_state_in_6 ? 8'hac : _GEN_6820; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6822 = 8'ha6 == io_state_in_6 ? 8'hbe : _GEN_6821; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6823 = 8'ha7 == io_state_in_6 ? 8'hb0 : _GEN_6822; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6824 = 8'ha8 == io_state_in_6 ? 8'hea : _GEN_6823; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6825 = 8'ha9 == io_state_in_6 ? 8'he4 : _GEN_6824; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6826 = 8'haa == io_state_in_6 ? 8'hf6 : _GEN_6825; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6827 = 8'hab == io_state_in_6 ? 8'hf8 : _GEN_6826; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6828 = 8'hac == io_state_in_6 ? 8'hd2 : _GEN_6827; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6829 = 8'had == io_state_in_6 ? 8'hdc : _GEN_6828; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6830 = 8'hae == io_state_in_6 ? 8'hce : _GEN_6829; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6831 = 8'haf == io_state_in_6 ? 8'hc0 : _GEN_6830; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6832 = 8'hb0 == io_state_in_6 ? 8'h7a : _GEN_6831; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6833 = 8'hb1 == io_state_in_6 ? 8'h74 : _GEN_6832; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6834 = 8'hb2 == io_state_in_6 ? 8'h66 : _GEN_6833; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6835 = 8'hb3 == io_state_in_6 ? 8'h68 : _GEN_6834; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6836 = 8'hb4 == io_state_in_6 ? 8'h42 : _GEN_6835; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6837 = 8'hb5 == io_state_in_6 ? 8'h4c : _GEN_6836; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6838 = 8'hb6 == io_state_in_6 ? 8'h5e : _GEN_6837; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6839 = 8'hb7 == io_state_in_6 ? 8'h50 : _GEN_6838; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6840 = 8'hb8 == io_state_in_6 ? 8'ha : _GEN_6839; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6841 = 8'hb9 == io_state_in_6 ? 8'h4 : _GEN_6840; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6842 = 8'hba == io_state_in_6 ? 8'h16 : _GEN_6841; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6843 = 8'hbb == io_state_in_6 ? 8'h18 : _GEN_6842; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6844 = 8'hbc == io_state_in_6 ? 8'h32 : _GEN_6843; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6845 = 8'hbd == io_state_in_6 ? 8'h3c : _GEN_6844; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6846 = 8'hbe == io_state_in_6 ? 8'h2e : _GEN_6845; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6847 = 8'hbf == io_state_in_6 ? 8'h20 : _GEN_6846; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6848 = 8'hc0 == io_state_in_6 ? 8'hec : _GEN_6847; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6849 = 8'hc1 == io_state_in_6 ? 8'he2 : _GEN_6848; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6850 = 8'hc2 == io_state_in_6 ? 8'hf0 : _GEN_6849; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6851 = 8'hc3 == io_state_in_6 ? 8'hfe : _GEN_6850; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6852 = 8'hc4 == io_state_in_6 ? 8'hd4 : _GEN_6851; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6853 = 8'hc5 == io_state_in_6 ? 8'hda : _GEN_6852; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6854 = 8'hc6 == io_state_in_6 ? 8'hc8 : _GEN_6853; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6855 = 8'hc7 == io_state_in_6 ? 8'hc6 : _GEN_6854; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6856 = 8'hc8 == io_state_in_6 ? 8'h9c : _GEN_6855; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6857 = 8'hc9 == io_state_in_6 ? 8'h92 : _GEN_6856; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6858 = 8'hca == io_state_in_6 ? 8'h80 : _GEN_6857; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6859 = 8'hcb == io_state_in_6 ? 8'h8e : _GEN_6858; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6860 = 8'hcc == io_state_in_6 ? 8'ha4 : _GEN_6859; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6861 = 8'hcd == io_state_in_6 ? 8'haa : _GEN_6860; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6862 = 8'hce == io_state_in_6 ? 8'hb8 : _GEN_6861; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6863 = 8'hcf == io_state_in_6 ? 8'hb6 : _GEN_6862; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6864 = 8'hd0 == io_state_in_6 ? 8'hc : _GEN_6863; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6865 = 8'hd1 == io_state_in_6 ? 8'h2 : _GEN_6864; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6866 = 8'hd2 == io_state_in_6 ? 8'h10 : _GEN_6865; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6867 = 8'hd3 == io_state_in_6 ? 8'h1e : _GEN_6866; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6868 = 8'hd4 == io_state_in_6 ? 8'h34 : _GEN_6867; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6869 = 8'hd5 == io_state_in_6 ? 8'h3a : _GEN_6868; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6870 = 8'hd6 == io_state_in_6 ? 8'h28 : _GEN_6869; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6871 = 8'hd7 == io_state_in_6 ? 8'h26 : _GEN_6870; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6872 = 8'hd8 == io_state_in_6 ? 8'h7c : _GEN_6871; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6873 = 8'hd9 == io_state_in_6 ? 8'h72 : _GEN_6872; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6874 = 8'hda == io_state_in_6 ? 8'h60 : _GEN_6873; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6875 = 8'hdb == io_state_in_6 ? 8'h6e : _GEN_6874; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6876 = 8'hdc == io_state_in_6 ? 8'h44 : _GEN_6875; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6877 = 8'hdd == io_state_in_6 ? 8'h4a : _GEN_6876; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6878 = 8'hde == io_state_in_6 ? 8'h58 : _GEN_6877; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6879 = 8'hdf == io_state_in_6 ? 8'h56 : _GEN_6878; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6880 = 8'he0 == io_state_in_6 ? 8'h37 : _GEN_6879; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6881 = 8'he1 == io_state_in_6 ? 8'h39 : _GEN_6880; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6882 = 8'he2 == io_state_in_6 ? 8'h2b : _GEN_6881; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6883 = 8'he3 == io_state_in_6 ? 8'h25 : _GEN_6882; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6884 = 8'he4 == io_state_in_6 ? 8'hf : _GEN_6883; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6885 = 8'he5 == io_state_in_6 ? 8'h1 : _GEN_6884; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6886 = 8'he6 == io_state_in_6 ? 8'h13 : _GEN_6885; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6887 = 8'he7 == io_state_in_6 ? 8'h1d : _GEN_6886; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6888 = 8'he8 == io_state_in_6 ? 8'h47 : _GEN_6887; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6889 = 8'he9 == io_state_in_6 ? 8'h49 : _GEN_6888; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6890 = 8'hea == io_state_in_6 ? 8'h5b : _GEN_6889; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6891 = 8'heb == io_state_in_6 ? 8'h55 : _GEN_6890; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6892 = 8'hec == io_state_in_6 ? 8'h7f : _GEN_6891; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6893 = 8'hed == io_state_in_6 ? 8'h71 : _GEN_6892; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6894 = 8'hee == io_state_in_6 ? 8'h63 : _GEN_6893; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6895 = 8'hef == io_state_in_6 ? 8'h6d : _GEN_6894; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6896 = 8'hf0 == io_state_in_6 ? 8'hd7 : _GEN_6895; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6897 = 8'hf1 == io_state_in_6 ? 8'hd9 : _GEN_6896; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6898 = 8'hf2 == io_state_in_6 ? 8'hcb : _GEN_6897; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6899 = 8'hf3 == io_state_in_6 ? 8'hc5 : _GEN_6898; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6900 = 8'hf4 == io_state_in_6 ? 8'hef : _GEN_6899; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6901 = 8'hf5 == io_state_in_6 ? 8'he1 : _GEN_6900; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6902 = 8'hf6 == io_state_in_6 ? 8'hf3 : _GEN_6901; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6903 = 8'hf7 == io_state_in_6 ? 8'hfd : _GEN_6902; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6904 = 8'hf8 == io_state_in_6 ? 8'ha7 : _GEN_6903; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6905 = 8'hf9 == io_state_in_6 ? 8'ha9 : _GEN_6904; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6906 = 8'hfa == io_state_in_6 ? 8'hbb : _GEN_6905; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6907 = 8'hfb == io_state_in_6 ? 8'hb5 : _GEN_6906; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6908 = 8'hfc == io_state_in_6 ? 8'h9f : _GEN_6907; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6909 = 8'hfd == io_state_in_6 ? 8'h91 : _GEN_6908; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6910 = 8'hfe == io_state_in_6 ? 8'h83 : _GEN_6909; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _GEN_6911 = 8'hff == io_state_in_6 ? 8'h8d : _GEN_6910; // @[InvMixColumns.scala 133:{65,65}]
  wire [7:0] _tmp_state_6_T_1 = _tmp_state_6_T ^ _GEN_6911; // @[InvMixColumns.scala 133:65]
  wire [7:0] _GEN_6913 = 8'h1 == io_state_in_7 ? 8'hb : 8'h0; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6914 = 8'h2 == io_state_in_7 ? 8'h16 : _GEN_6913; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6915 = 8'h3 == io_state_in_7 ? 8'h1d : _GEN_6914; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6916 = 8'h4 == io_state_in_7 ? 8'h2c : _GEN_6915; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6917 = 8'h5 == io_state_in_7 ? 8'h27 : _GEN_6916; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6918 = 8'h6 == io_state_in_7 ? 8'h3a : _GEN_6917; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6919 = 8'h7 == io_state_in_7 ? 8'h31 : _GEN_6918; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6920 = 8'h8 == io_state_in_7 ? 8'h58 : _GEN_6919; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6921 = 8'h9 == io_state_in_7 ? 8'h53 : _GEN_6920; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6922 = 8'ha == io_state_in_7 ? 8'h4e : _GEN_6921; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6923 = 8'hb == io_state_in_7 ? 8'h45 : _GEN_6922; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6924 = 8'hc == io_state_in_7 ? 8'h74 : _GEN_6923; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6925 = 8'hd == io_state_in_7 ? 8'h7f : _GEN_6924; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6926 = 8'he == io_state_in_7 ? 8'h62 : _GEN_6925; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6927 = 8'hf == io_state_in_7 ? 8'h69 : _GEN_6926; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6928 = 8'h10 == io_state_in_7 ? 8'hb0 : _GEN_6927; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6929 = 8'h11 == io_state_in_7 ? 8'hbb : _GEN_6928; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6930 = 8'h12 == io_state_in_7 ? 8'ha6 : _GEN_6929; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6931 = 8'h13 == io_state_in_7 ? 8'had : _GEN_6930; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6932 = 8'h14 == io_state_in_7 ? 8'h9c : _GEN_6931; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6933 = 8'h15 == io_state_in_7 ? 8'h97 : _GEN_6932; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6934 = 8'h16 == io_state_in_7 ? 8'h8a : _GEN_6933; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6935 = 8'h17 == io_state_in_7 ? 8'h81 : _GEN_6934; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6936 = 8'h18 == io_state_in_7 ? 8'he8 : _GEN_6935; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6937 = 8'h19 == io_state_in_7 ? 8'he3 : _GEN_6936; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6938 = 8'h1a == io_state_in_7 ? 8'hfe : _GEN_6937; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6939 = 8'h1b == io_state_in_7 ? 8'hf5 : _GEN_6938; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6940 = 8'h1c == io_state_in_7 ? 8'hc4 : _GEN_6939; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6941 = 8'h1d == io_state_in_7 ? 8'hcf : _GEN_6940; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6942 = 8'h1e == io_state_in_7 ? 8'hd2 : _GEN_6941; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6943 = 8'h1f == io_state_in_7 ? 8'hd9 : _GEN_6942; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6944 = 8'h20 == io_state_in_7 ? 8'h7b : _GEN_6943; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6945 = 8'h21 == io_state_in_7 ? 8'h70 : _GEN_6944; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6946 = 8'h22 == io_state_in_7 ? 8'h6d : _GEN_6945; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6947 = 8'h23 == io_state_in_7 ? 8'h66 : _GEN_6946; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6948 = 8'h24 == io_state_in_7 ? 8'h57 : _GEN_6947; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6949 = 8'h25 == io_state_in_7 ? 8'h5c : _GEN_6948; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6950 = 8'h26 == io_state_in_7 ? 8'h41 : _GEN_6949; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6951 = 8'h27 == io_state_in_7 ? 8'h4a : _GEN_6950; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6952 = 8'h28 == io_state_in_7 ? 8'h23 : _GEN_6951; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6953 = 8'h29 == io_state_in_7 ? 8'h28 : _GEN_6952; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6954 = 8'h2a == io_state_in_7 ? 8'h35 : _GEN_6953; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6955 = 8'h2b == io_state_in_7 ? 8'h3e : _GEN_6954; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6956 = 8'h2c == io_state_in_7 ? 8'hf : _GEN_6955; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6957 = 8'h2d == io_state_in_7 ? 8'h4 : _GEN_6956; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6958 = 8'h2e == io_state_in_7 ? 8'h19 : _GEN_6957; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6959 = 8'h2f == io_state_in_7 ? 8'h12 : _GEN_6958; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6960 = 8'h30 == io_state_in_7 ? 8'hcb : _GEN_6959; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6961 = 8'h31 == io_state_in_7 ? 8'hc0 : _GEN_6960; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6962 = 8'h32 == io_state_in_7 ? 8'hdd : _GEN_6961; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6963 = 8'h33 == io_state_in_7 ? 8'hd6 : _GEN_6962; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6964 = 8'h34 == io_state_in_7 ? 8'he7 : _GEN_6963; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6965 = 8'h35 == io_state_in_7 ? 8'hec : _GEN_6964; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6966 = 8'h36 == io_state_in_7 ? 8'hf1 : _GEN_6965; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6967 = 8'h37 == io_state_in_7 ? 8'hfa : _GEN_6966; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6968 = 8'h38 == io_state_in_7 ? 8'h93 : _GEN_6967; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6969 = 8'h39 == io_state_in_7 ? 8'h98 : _GEN_6968; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6970 = 8'h3a == io_state_in_7 ? 8'h85 : _GEN_6969; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6971 = 8'h3b == io_state_in_7 ? 8'h8e : _GEN_6970; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6972 = 8'h3c == io_state_in_7 ? 8'hbf : _GEN_6971; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6973 = 8'h3d == io_state_in_7 ? 8'hb4 : _GEN_6972; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6974 = 8'h3e == io_state_in_7 ? 8'ha9 : _GEN_6973; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6975 = 8'h3f == io_state_in_7 ? 8'ha2 : _GEN_6974; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6976 = 8'h40 == io_state_in_7 ? 8'hf6 : _GEN_6975; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6977 = 8'h41 == io_state_in_7 ? 8'hfd : _GEN_6976; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6978 = 8'h42 == io_state_in_7 ? 8'he0 : _GEN_6977; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6979 = 8'h43 == io_state_in_7 ? 8'heb : _GEN_6978; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6980 = 8'h44 == io_state_in_7 ? 8'hda : _GEN_6979; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6981 = 8'h45 == io_state_in_7 ? 8'hd1 : _GEN_6980; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6982 = 8'h46 == io_state_in_7 ? 8'hcc : _GEN_6981; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6983 = 8'h47 == io_state_in_7 ? 8'hc7 : _GEN_6982; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6984 = 8'h48 == io_state_in_7 ? 8'hae : _GEN_6983; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6985 = 8'h49 == io_state_in_7 ? 8'ha5 : _GEN_6984; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6986 = 8'h4a == io_state_in_7 ? 8'hb8 : _GEN_6985; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6987 = 8'h4b == io_state_in_7 ? 8'hb3 : _GEN_6986; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6988 = 8'h4c == io_state_in_7 ? 8'h82 : _GEN_6987; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6989 = 8'h4d == io_state_in_7 ? 8'h89 : _GEN_6988; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6990 = 8'h4e == io_state_in_7 ? 8'h94 : _GEN_6989; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6991 = 8'h4f == io_state_in_7 ? 8'h9f : _GEN_6990; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6992 = 8'h50 == io_state_in_7 ? 8'h46 : _GEN_6991; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6993 = 8'h51 == io_state_in_7 ? 8'h4d : _GEN_6992; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6994 = 8'h52 == io_state_in_7 ? 8'h50 : _GEN_6993; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6995 = 8'h53 == io_state_in_7 ? 8'h5b : _GEN_6994; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6996 = 8'h54 == io_state_in_7 ? 8'h6a : _GEN_6995; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6997 = 8'h55 == io_state_in_7 ? 8'h61 : _GEN_6996; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6998 = 8'h56 == io_state_in_7 ? 8'h7c : _GEN_6997; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_6999 = 8'h57 == io_state_in_7 ? 8'h77 : _GEN_6998; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7000 = 8'h58 == io_state_in_7 ? 8'h1e : _GEN_6999; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7001 = 8'h59 == io_state_in_7 ? 8'h15 : _GEN_7000; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7002 = 8'h5a == io_state_in_7 ? 8'h8 : _GEN_7001; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7003 = 8'h5b == io_state_in_7 ? 8'h3 : _GEN_7002; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7004 = 8'h5c == io_state_in_7 ? 8'h32 : _GEN_7003; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7005 = 8'h5d == io_state_in_7 ? 8'h39 : _GEN_7004; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7006 = 8'h5e == io_state_in_7 ? 8'h24 : _GEN_7005; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7007 = 8'h5f == io_state_in_7 ? 8'h2f : _GEN_7006; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7008 = 8'h60 == io_state_in_7 ? 8'h8d : _GEN_7007; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7009 = 8'h61 == io_state_in_7 ? 8'h86 : _GEN_7008; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7010 = 8'h62 == io_state_in_7 ? 8'h9b : _GEN_7009; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7011 = 8'h63 == io_state_in_7 ? 8'h90 : _GEN_7010; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7012 = 8'h64 == io_state_in_7 ? 8'ha1 : _GEN_7011; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7013 = 8'h65 == io_state_in_7 ? 8'haa : _GEN_7012; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7014 = 8'h66 == io_state_in_7 ? 8'hb7 : _GEN_7013; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7015 = 8'h67 == io_state_in_7 ? 8'hbc : _GEN_7014; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7016 = 8'h68 == io_state_in_7 ? 8'hd5 : _GEN_7015; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7017 = 8'h69 == io_state_in_7 ? 8'hde : _GEN_7016; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7018 = 8'h6a == io_state_in_7 ? 8'hc3 : _GEN_7017; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7019 = 8'h6b == io_state_in_7 ? 8'hc8 : _GEN_7018; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7020 = 8'h6c == io_state_in_7 ? 8'hf9 : _GEN_7019; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7021 = 8'h6d == io_state_in_7 ? 8'hf2 : _GEN_7020; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7022 = 8'h6e == io_state_in_7 ? 8'hef : _GEN_7021; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7023 = 8'h6f == io_state_in_7 ? 8'he4 : _GEN_7022; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7024 = 8'h70 == io_state_in_7 ? 8'h3d : _GEN_7023; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7025 = 8'h71 == io_state_in_7 ? 8'h36 : _GEN_7024; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7026 = 8'h72 == io_state_in_7 ? 8'h2b : _GEN_7025; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7027 = 8'h73 == io_state_in_7 ? 8'h20 : _GEN_7026; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7028 = 8'h74 == io_state_in_7 ? 8'h11 : _GEN_7027; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7029 = 8'h75 == io_state_in_7 ? 8'h1a : _GEN_7028; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7030 = 8'h76 == io_state_in_7 ? 8'h7 : _GEN_7029; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7031 = 8'h77 == io_state_in_7 ? 8'hc : _GEN_7030; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7032 = 8'h78 == io_state_in_7 ? 8'h65 : _GEN_7031; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7033 = 8'h79 == io_state_in_7 ? 8'h6e : _GEN_7032; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7034 = 8'h7a == io_state_in_7 ? 8'h73 : _GEN_7033; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7035 = 8'h7b == io_state_in_7 ? 8'h78 : _GEN_7034; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7036 = 8'h7c == io_state_in_7 ? 8'h49 : _GEN_7035; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7037 = 8'h7d == io_state_in_7 ? 8'h42 : _GEN_7036; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7038 = 8'h7e == io_state_in_7 ? 8'h5f : _GEN_7037; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7039 = 8'h7f == io_state_in_7 ? 8'h54 : _GEN_7038; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7040 = 8'h80 == io_state_in_7 ? 8'hf7 : _GEN_7039; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7041 = 8'h81 == io_state_in_7 ? 8'hfc : _GEN_7040; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7042 = 8'h82 == io_state_in_7 ? 8'he1 : _GEN_7041; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7043 = 8'h83 == io_state_in_7 ? 8'hea : _GEN_7042; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7044 = 8'h84 == io_state_in_7 ? 8'hdb : _GEN_7043; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7045 = 8'h85 == io_state_in_7 ? 8'hd0 : _GEN_7044; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7046 = 8'h86 == io_state_in_7 ? 8'hcd : _GEN_7045; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7047 = 8'h87 == io_state_in_7 ? 8'hc6 : _GEN_7046; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7048 = 8'h88 == io_state_in_7 ? 8'haf : _GEN_7047; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7049 = 8'h89 == io_state_in_7 ? 8'ha4 : _GEN_7048; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7050 = 8'h8a == io_state_in_7 ? 8'hb9 : _GEN_7049; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7051 = 8'h8b == io_state_in_7 ? 8'hb2 : _GEN_7050; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7052 = 8'h8c == io_state_in_7 ? 8'h83 : _GEN_7051; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7053 = 8'h8d == io_state_in_7 ? 8'h88 : _GEN_7052; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7054 = 8'h8e == io_state_in_7 ? 8'h95 : _GEN_7053; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7055 = 8'h8f == io_state_in_7 ? 8'h9e : _GEN_7054; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7056 = 8'h90 == io_state_in_7 ? 8'h47 : _GEN_7055; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7057 = 8'h91 == io_state_in_7 ? 8'h4c : _GEN_7056; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7058 = 8'h92 == io_state_in_7 ? 8'h51 : _GEN_7057; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7059 = 8'h93 == io_state_in_7 ? 8'h5a : _GEN_7058; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7060 = 8'h94 == io_state_in_7 ? 8'h6b : _GEN_7059; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7061 = 8'h95 == io_state_in_7 ? 8'h60 : _GEN_7060; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7062 = 8'h96 == io_state_in_7 ? 8'h7d : _GEN_7061; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7063 = 8'h97 == io_state_in_7 ? 8'h76 : _GEN_7062; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7064 = 8'h98 == io_state_in_7 ? 8'h1f : _GEN_7063; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7065 = 8'h99 == io_state_in_7 ? 8'h14 : _GEN_7064; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7066 = 8'h9a == io_state_in_7 ? 8'h9 : _GEN_7065; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7067 = 8'h9b == io_state_in_7 ? 8'h2 : _GEN_7066; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7068 = 8'h9c == io_state_in_7 ? 8'h33 : _GEN_7067; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7069 = 8'h9d == io_state_in_7 ? 8'h38 : _GEN_7068; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7070 = 8'h9e == io_state_in_7 ? 8'h25 : _GEN_7069; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7071 = 8'h9f == io_state_in_7 ? 8'h2e : _GEN_7070; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7072 = 8'ha0 == io_state_in_7 ? 8'h8c : _GEN_7071; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7073 = 8'ha1 == io_state_in_7 ? 8'h87 : _GEN_7072; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7074 = 8'ha2 == io_state_in_7 ? 8'h9a : _GEN_7073; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7075 = 8'ha3 == io_state_in_7 ? 8'h91 : _GEN_7074; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7076 = 8'ha4 == io_state_in_7 ? 8'ha0 : _GEN_7075; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7077 = 8'ha5 == io_state_in_7 ? 8'hab : _GEN_7076; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7078 = 8'ha6 == io_state_in_7 ? 8'hb6 : _GEN_7077; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7079 = 8'ha7 == io_state_in_7 ? 8'hbd : _GEN_7078; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7080 = 8'ha8 == io_state_in_7 ? 8'hd4 : _GEN_7079; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7081 = 8'ha9 == io_state_in_7 ? 8'hdf : _GEN_7080; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7082 = 8'haa == io_state_in_7 ? 8'hc2 : _GEN_7081; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7083 = 8'hab == io_state_in_7 ? 8'hc9 : _GEN_7082; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7084 = 8'hac == io_state_in_7 ? 8'hf8 : _GEN_7083; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7085 = 8'had == io_state_in_7 ? 8'hf3 : _GEN_7084; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7086 = 8'hae == io_state_in_7 ? 8'hee : _GEN_7085; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7087 = 8'haf == io_state_in_7 ? 8'he5 : _GEN_7086; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7088 = 8'hb0 == io_state_in_7 ? 8'h3c : _GEN_7087; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7089 = 8'hb1 == io_state_in_7 ? 8'h37 : _GEN_7088; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7090 = 8'hb2 == io_state_in_7 ? 8'h2a : _GEN_7089; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7091 = 8'hb3 == io_state_in_7 ? 8'h21 : _GEN_7090; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7092 = 8'hb4 == io_state_in_7 ? 8'h10 : _GEN_7091; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7093 = 8'hb5 == io_state_in_7 ? 8'h1b : _GEN_7092; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7094 = 8'hb6 == io_state_in_7 ? 8'h6 : _GEN_7093; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7095 = 8'hb7 == io_state_in_7 ? 8'hd : _GEN_7094; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7096 = 8'hb8 == io_state_in_7 ? 8'h64 : _GEN_7095; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7097 = 8'hb9 == io_state_in_7 ? 8'h6f : _GEN_7096; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7098 = 8'hba == io_state_in_7 ? 8'h72 : _GEN_7097; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7099 = 8'hbb == io_state_in_7 ? 8'h79 : _GEN_7098; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7100 = 8'hbc == io_state_in_7 ? 8'h48 : _GEN_7099; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7101 = 8'hbd == io_state_in_7 ? 8'h43 : _GEN_7100; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7102 = 8'hbe == io_state_in_7 ? 8'h5e : _GEN_7101; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7103 = 8'hbf == io_state_in_7 ? 8'h55 : _GEN_7102; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7104 = 8'hc0 == io_state_in_7 ? 8'h1 : _GEN_7103; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7105 = 8'hc1 == io_state_in_7 ? 8'ha : _GEN_7104; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7106 = 8'hc2 == io_state_in_7 ? 8'h17 : _GEN_7105; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7107 = 8'hc3 == io_state_in_7 ? 8'h1c : _GEN_7106; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7108 = 8'hc4 == io_state_in_7 ? 8'h2d : _GEN_7107; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7109 = 8'hc5 == io_state_in_7 ? 8'h26 : _GEN_7108; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7110 = 8'hc6 == io_state_in_7 ? 8'h3b : _GEN_7109; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7111 = 8'hc7 == io_state_in_7 ? 8'h30 : _GEN_7110; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7112 = 8'hc8 == io_state_in_7 ? 8'h59 : _GEN_7111; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7113 = 8'hc9 == io_state_in_7 ? 8'h52 : _GEN_7112; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7114 = 8'hca == io_state_in_7 ? 8'h4f : _GEN_7113; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7115 = 8'hcb == io_state_in_7 ? 8'h44 : _GEN_7114; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7116 = 8'hcc == io_state_in_7 ? 8'h75 : _GEN_7115; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7117 = 8'hcd == io_state_in_7 ? 8'h7e : _GEN_7116; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7118 = 8'hce == io_state_in_7 ? 8'h63 : _GEN_7117; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7119 = 8'hcf == io_state_in_7 ? 8'h68 : _GEN_7118; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7120 = 8'hd0 == io_state_in_7 ? 8'hb1 : _GEN_7119; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7121 = 8'hd1 == io_state_in_7 ? 8'hba : _GEN_7120; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7122 = 8'hd2 == io_state_in_7 ? 8'ha7 : _GEN_7121; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7123 = 8'hd3 == io_state_in_7 ? 8'hac : _GEN_7122; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7124 = 8'hd4 == io_state_in_7 ? 8'h9d : _GEN_7123; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7125 = 8'hd5 == io_state_in_7 ? 8'h96 : _GEN_7124; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7126 = 8'hd6 == io_state_in_7 ? 8'h8b : _GEN_7125; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7127 = 8'hd7 == io_state_in_7 ? 8'h80 : _GEN_7126; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7128 = 8'hd8 == io_state_in_7 ? 8'he9 : _GEN_7127; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7129 = 8'hd9 == io_state_in_7 ? 8'he2 : _GEN_7128; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7130 = 8'hda == io_state_in_7 ? 8'hff : _GEN_7129; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7131 = 8'hdb == io_state_in_7 ? 8'hf4 : _GEN_7130; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7132 = 8'hdc == io_state_in_7 ? 8'hc5 : _GEN_7131; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7133 = 8'hdd == io_state_in_7 ? 8'hce : _GEN_7132; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7134 = 8'hde == io_state_in_7 ? 8'hd3 : _GEN_7133; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7135 = 8'hdf == io_state_in_7 ? 8'hd8 : _GEN_7134; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7136 = 8'he0 == io_state_in_7 ? 8'h7a : _GEN_7135; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7137 = 8'he1 == io_state_in_7 ? 8'h71 : _GEN_7136; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7138 = 8'he2 == io_state_in_7 ? 8'h6c : _GEN_7137; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7139 = 8'he3 == io_state_in_7 ? 8'h67 : _GEN_7138; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7140 = 8'he4 == io_state_in_7 ? 8'h56 : _GEN_7139; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7141 = 8'he5 == io_state_in_7 ? 8'h5d : _GEN_7140; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7142 = 8'he6 == io_state_in_7 ? 8'h40 : _GEN_7141; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7143 = 8'he7 == io_state_in_7 ? 8'h4b : _GEN_7142; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7144 = 8'he8 == io_state_in_7 ? 8'h22 : _GEN_7143; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7145 = 8'he9 == io_state_in_7 ? 8'h29 : _GEN_7144; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7146 = 8'hea == io_state_in_7 ? 8'h34 : _GEN_7145; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7147 = 8'heb == io_state_in_7 ? 8'h3f : _GEN_7146; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7148 = 8'hec == io_state_in_7 ? 8'he : _GEN_7147; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7149 = 8'hed == io_state_in_7 ? 8'h5 : _GEN_7148; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7150 = 8'hee == io_state_in_7 ? 8'h18 : _GEN_7149; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7151 = 8'hef == io_state_in_7 ? 8'h13 : _GEN_7150; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7152 = 8'hf0 == io_state_in_7 ? 8'hca : _GEN_7151; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7153 = 8'hf1 == io_state_in_7 ? 8'hc1 : _GEN_7152; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7154 = 8'hf2 == io_state_in_7 ? 8'hdc : _GEN_7153; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7155 = 8'hf3 == io_state_in_7 ? 8'hd7 : _GEN_7154; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7156 = 8'hf4 == io_state_in_7 ? 8'he6 : _GEN_7155; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7157 = 8'hf5 == io_state_in_7 ? 8'hed : _GEN_7156; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7158 = 8'hf6 == io_state_in_7 ? 8'hf0 : _GEN_7157; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7159 = 8'hf7 == io_state_in_7 ? 8'hfb : _GEN_7158; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7160 = 8'hf8 == io_state_in_7 ? 8'h92 : _GEN_7159; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7161 = 8'hf9 == io_state_in_7 ? 8'h99 : _GEN_7160; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7162 = 8'hfa == io_state_in_7 ? 8'h84 : _GEN_7161; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7163 = 8'hfb == io_state_in_7 ? 8'h8f : _GEN_7162; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7164 = 8'hfc == io_state_in_7 ? 8'hbe : _GEN_7163; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7165 = 8'hfd == io_state_in_7 ? 8'hb5 : _GEN_7164; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7166 = 8'hfe == io_state_in_7 ? 8'ha8 : _GEN_7165; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7167 = 8'hff == io_state_in_7 ? 8'ha3 : _GEN_7166; // @[InvMixColumns.scala 133:{89,89}]
  wire [7:0] _GEN_7169 = 8'h1 == io_state_in_4 ? 8'hb : 8'h0; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7170 = 8'h2 == io_state_in_4 ? 8'h16 : _GEN_7169; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7171 = 8'h3 == io_state_in_4 ? 8'h1d : _GEN_7170; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7172 = 8'h4 == io_state_in_4 ? 8'h2c : _GEN_7171; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7173 = 8'h5 == io_state_in_4 ? 8'h27 : _GEN_7172; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7174 = 8'h6 == io_state_in_4 ? 8'h3a : _GEN_7173; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7175 = 8'h7 == io_state_in_4 ? 8'h31 : _GEN_7174; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7176 = 8'h8 == io_state_in_4 ? 8'h58 : _GEN_7175; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7177 = 8'h9 == io_state_in_4 ? 8'h53 : _GEN_7176; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7178 = 8'ha == io_state_in_4 ? 8'h4e : _GEN_7177; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7179 = 8'hb == io_state_in_4 ? 8'h45 : _GEN_7178; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7180 = 8'hc == io_state_in_4 ? 8'h74 : _GEN_7179; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7181 = 8'hd == io_state_in_4 ? 8'h7f : _GEN_7180; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7182 = 8'he == io_state_in_4 ? 8'h62 : _GEN_7181; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7183 = 8'hf == io_state_in_4 ? 8'h69 : _GEN_7182; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7184 = 8'h10 == io_state_in_4 ? 8'hb0 : _GEN_7183; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7185 = 8'h11 == io_state_in_4 ? 8'hbb : _GEN_7184; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7186 = 8'h12 == io_state_in_4 ? 8'ha6 : _GEN_7185; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7187 = 8'h13 == io_state_in_4 ? 8'had : _GEN_7186; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7188 = 8'h14 == io_state_in_4 ? 8'h9c : _GEN_7187; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7189 = 8'h15 == io_state_in_4 ? 8'h97 : _GEN_7188; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7190 = 8'h16 == io_state_in_4 ? 8'h8a : _GEN_7189; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7191 = 8'h17 == io_state_in_4 ? 8'h81 : _GEN_7190; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7192 = 8'h18 == io_state_in_4 ? 8'he8 : _GEN_7191; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7193 = 8'h19 == io_state_in_4 ? 8'he3 : _GEN_7192; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7194 = 8'h1a == io_state_in_4 ? 8'hfe : _GEN_7193; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7195 = 8'h1b == io_state_in_4 ? 8'hf5 : _GEN_7194; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7196 = 8'h1c == io_state_in_4 ? 8'hc4 : _GEN_7195; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7197 = 8'h1d == io_state_in_4 ? 8'hcf : _GEN_7196; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7198 = 8'h1e == io_state_in_4 ? 8'hd2 : _GEN_7197; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7199 = 8'h1f == io_state_in_4 ? 8'hd9 : _GEN_7198; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7200 = 8'h20 == io_state_in_4 ? 8'h7b : _GEN_7199; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7201 = 8'h21 == io_state_in_4 ? 8'h70 : _GEN_7200; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7202 = 8'h22 == io_state_in_4 ? 8'h6d : _GEN_7201; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7203 = 8'h23 == io_state_in_4 ? 8'h66 : _GEN_7202; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7204 = 8'h24 == io_state_in_4 ? 8'h57 : _GEN_7203; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7205 = 8'h25 == io_state_in_4 ? 8'h5c : _GEN_7204; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7206 = 8'h26 == io_state_in_4 ? 8'h41 : _GEN_7205; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7207 = 8'h27 == io_state_in_4 ? 8'h4a : _GEN_7206; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7208 = 8'h28 == io_state_in_4 ? 8'h23 : _GEN_7207; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7209 = 8'h29 == io_state_in_4 ? 8'h28 : _GEN_7208; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7210 = 8'h2a == io_state_in_4 ? 8'h35 : _GEN_7209; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7211 = 8'h2b == io_state_in_4 ? 8'h3e : _GEN_7210; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7212 = 8'h2c == io_state_in_4 ? 8'hf : _GEN_7211; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7213 = 8'h2d == io_state_in_4 ? 8'h4 : _GEN_7212; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7214 = 8'h2e == io_state_in_4 ? 8'h19 : _GEN_7213; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7215 = 8'h2f == io_state_in_4 ? 8'h12 : _GEN_7214; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7216 = 8'h30 == io_state_in_4 ? 8'hcb : _GEN_7215; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7217 = 8'h31 == io_state_in_4 ? 8'hc0 : _GEN_7216; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7218 = 8'h32 == io_state_in_4 ? 8'hdd : _GEN_7217; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7219 = 8'h33 == io_state_in_4 ? 8'hd6 : _GEN_7218; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7220 = 8'h34 == io_state_in_4 ? 8'he7 : _GEN_7219; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7221 = 8'h35 == io_state_in_4 ? 8'hec : _GEN_7220; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7222 = 8'h36 == io_state_in_4 ? 8'hf1 : _GEN_7221; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7223 = 8'h37 == io_state_in_4 ? 8'hfa : _GEN_7222; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7224 = 8'h38 == io_state_in_4 ? 8'h93 : _GEN_7223; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7225 = 8'h39 == io_state_in_4 ? 8'h98 : _GEN_7224; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7226 = 8'h3a == io_state_in_4 ? 8'h85 : _GEN_7225; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7227 = 8'h3b == io_state_in_4 ? 8'h8e : _GEN_7226; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7228 = 8'h3c == io_state_in_4 ? 8'hbf : _GEN_7227; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7229 = 8'h3d == io_state_in_4 ? 8'hb4 : _GEN_7228; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7230 = 8'h3e == io_state_in_4 ? 8'ha9 : _GEN_7229; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7231 = 8'h3f == io_state_in_4 ? 8'ha2 : _GEN_7230; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7232 = 8'h40 == io_state_in_4 ? 8'hf6 : _GEN_7231; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7233 = 8'h41 == io_state_in_4 ? 8'hfd : _GEN_7232; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7234 = 8'h42 == io_state_in_4 ? 8'he0 : _GEN_7233; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7235 = 8'h43 == io_state_in_4 ? 8'heb : _GEN_7234; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7236 = 8'h44 == io_state_in_4 ? 8'hda : _GEN_7235; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7237 = 8'h45 == io_state_in_4 ? 8'hd1 : _GEN_7236; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7238 = 8'h46 == io_state_in_4 ? 8'hcc : _GEN_7237; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7239 = 8'h47 == io_state_in_4 ? 8'hc7 : _GEN_7238; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7240 = 8'h48 == io_state_in_4 ? 8'hae : _GEN_7239; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7241 = 8'h49 == io_state_in_4 ? 8'ha5 : _GEN_7240; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7242 = 8'h4a == io_state_in_4 ? 8'hb8 : _GEN_7241; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7243 = 8'h4b == io_state_in_4 ? 8'hb3 : _GEN_7242; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7244 = 8'h4c == io_state_in_4 ? 8'h82 : _GEN_7243; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7245 = 8'h4d == io_state_in_4 ? 8'h89 : _GEN_7244; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7246 = 8'h4e == io_state_in_4 ? 8'h94 : _GEN_7245; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7247 = 8'h4f == io_state_in_4 ? 8'h9f : _GEN_7246; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7248 = 8'h50 == io_state_in_4 ? 8'h46 : _GEN_7247; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7249 = 8'h51 == io_state_in_4 ? 8'h4d : _GEN_7248; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7250 = 8'h52 == io_state_in_4 ? 8'h50 : _GEN_7249; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7251 = 8'h53 == io_state_in_4 ? 8'h5b : _GEN_7250; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7252 = 8'h54 == io_state_in_4 ? 8'h6a : _GEN_7251; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7253 = 8'h55 == io_state_in_4 ? 8'h61 : _GEN_7252; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7254 = 8'h56 == io_state_in_4 ? 8'h7c : _GEN_7253; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7255 = 8'h57 == io_state_in_4 ? 8'h77 : _GEN_7254; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7256 = 8'h58 == io_state_in_4 ? 8'h1e : _GEN_7255; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7257 = 8'h59 == io_state_in_4 ? 8'h15 : _GEN_7256; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7258 = 8'h5a == io_state_in_4 ? 8'h8 : _GEN_7257; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7259 = 8'h5b == io_state_in_4 ? 8'h3 : _GEN_7258; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7260 = 8'h5c == io_state_in_4 ? 8'h32 : _GEN_7259; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7261 = 8'h5d == io_state_in_4 ? 8'h39 : _GEN_7260; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7262 = 8'h5e == io_state_in_4 ? 8'h24 : _GEN_7261; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7263 = 8'h5f == io_state_in_4 ? 8'h2f : _GEN_7262; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7264 = 8'h60 == io_state_in_4 ? 8'h8d : _GEN_7263; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7265 = 8'h61 == io_state_in_4 ? 8'h86 : _GEN_7264; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7266 = 8'h62 == io_state_in_4 ? 8'h9b : _GEN_7265; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7267 = 8'h63 == io_state_in_4 ? 8'h90 : _GEN_7266; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7268 = 8'h64 == io_state_in_4 ? 8'ha1 : _GEN_7267; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7269 = 8'h65 == io_state_in_4 ? 8'haa : _GEN_7268; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7270 = 8'h66 == io_state_in_4 ? 8'hb7 : _GEN_7269; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7271 = 8'h67 == io_state_in_4 ? 8'hbc : _GEN_7270; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7272 = 8'h68 == io_state_in_4 ? 8'hd5 : _GEN_7271; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7273 = 8'h69 == io_state_in_4 ? 8'hde : _GEN_7272; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7274 = 8'h6a == io_state_in_4 ? 8'hc3 : _GEN_7273; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7275 = 8'h6b == io_state_in_4 ? 8'hc8 : _GEN_7274; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7276 = 8'h6c == io_state_in_4 ? 8'hf9 : _GEN_7275; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7277 = 8'h6d == io_state_in_4 ? 8'hf2 : _GEN_7276; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7278 = 8'h6e == io_state_in_4 ? 8'hef : _GEN_7277; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7279 = 8'h6f == io_state_in_4 ? 8'he4 : _GEN_7278; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7280 = 8'h70 == io_state_in_4 ? 8'h3d : _GEN_7279; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7281 = 8'h71 == io_state_in_4 ? 8'h36 : _GEN_7280; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7282 = 8'h72 == io_state_in_4 ? 8'h2b : _GEN_7281; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7283 = 8'h73 == io_state_in_4 ? 8'h20 : _GEN_7282; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7284 = 8'h74 == io_state_in_4 ? 8'h11 : _GEN_7283; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7285 = 8'h75 == io_state_in_4 ? 8'h1a : _GEN_7284; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7286 = 8'h76 == io_state_in_4 ? 8'h7 : _GEN_7285; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7287 = 8'h77 == io_state_in_4 ? 8'hc : _GEN_7286; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7288 = 8'h78 == io_state_in_4 ? 8'h65 : _GEN_7287; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7289 = 8'h79 == io_state_in_4 ? 8'h6e : _GEN_7288; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7290 = 8'h7a == io_state_in_4 ? 8'h73 : _GEN_7289; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7291 = 8'h7b == io_state_in_4 ? 8'h78 : _GEN_7290; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7292 = 8'h7c == io_state_in_4 ? 8'h49 : _GEN_7291; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7293 = 8'h7d == io_state_in_4 ? 8'h42 : _GEN_7292; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7294 = 8'h7e == io_state_in_4 ? 8'h5f : _GEN_7293; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7295 = 8'h7f == io_state_in_4 ? 8'h54 : _GEN_7294; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7296 = 8'h80 == io_state_in_4 ? 8'hf7 : _GEN_7295; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7297 = 8'h81 == io_state_in_4 ? 8'hfc : _GEN_7296; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7298 = 8'h82 == io_state_in_4 ? 8'he1 : _GEN_7297; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7299 = 8'h83 == io_state_in_4 ? 8'hea : _GEN_7298; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7300 = 8'h84 == io_state_in_4 ? 8'hdb : _GEN_7299; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7301 = 8'h85 == io_state_in_4 ? 8'hd0 : _GEN_7300; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7302 = 8'h86 == io_state_in_4 ? 8'hcd : _GEN_7301; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7303 = 8'h87 == io_state_in_4 ? 8'hc6 : _GEN_7302; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7304 = 8'h88 == io_state_in_4 ? 8'haf : _GEN_7303; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7305 = 8'h89 == io_state_in_4 ? 8'ha4 : _GEN_7304; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7306 = 8'h8a == io_state_in_4 ? 8'hb9 : _GEN_7305; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7307 = 8'h8b == io_state_in_4 ? 8'hb2 : _GEN_7306; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7308 = 8'h8c == io_state_in_4 ? 8'h83 : _GEN_7307; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7309 = 8'h8d == io_state_in_4 ? 8'h88 : _GEN_7308; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7310 = 8'h8e == io_state_in_4 ? 8'h95 : _GEN_7309; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7311 = 8'h8f == io_state_in_4 ? 8'h9e : _GEN_7310; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7312 = 8'h90 == io_state_in_4 ? 8'h47 : _GEN_7311; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7313 = 8'h91 == io_state_in_4 ? 8'h4c : _GEN_7312; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7314 = 8'h92 == io_state_in_4 ? 8'h51 : _GEN_7313; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7315 = 8'h93 == io_state_in_4 ? 8'h5a : _GEN_7314; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7316 = 8'h94 == io_state_in_4 ? 8'h6b : _GEN_7315; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7317 = 8'h95 == io_state_in_4 ? 8'h60 : _GEN_7316; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7318 = 8'h96 == io_state_in_4 ? 8'h7d : _GEN_7317; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7319 = 8'h97 == io_state_in_4 ? 8'h76 : _GEN_7318; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7320 = 8'h98 == io_state_in_4 ? 8'h1f : _GEN_7319; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7321 = 8'h99 == io_state_in_4 ? 8'h14 : _GEN_7320; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7322 = 8'h9a == io_state_in_4 ? 8'h9 : _GEN_7321; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7323 = 8'h9b == io_state_in_4 ? 8'h2 : _GEN_7322; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7324 = 8'h9c == io_state_in_4 ? 8'h33 : _GEN_7323; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7325 = 8'h9d == io_state_in_4 ? 8'h38 : _GEN_7324; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7326 = 8'h9e == io_state_in_4 ? 8'h25 : _GEN_7325; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7327 = 8'h9f == io_state_in_4 ? 8'h2e : _GEN_7326; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7328 = 8'ha0 == io_state_in_4 ? 8'h8c : _GEN_7327; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7329 = 8'ha1 == io_state_in_4 ? 8'h87 : _GEN_7328; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7330 = 8'ha2 == io_state_in_4 ? 8'h9a : _GEN_7329; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7331 = 8'ha3 == io_state_in_4 ? 8'h91 : _GEN_7330; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7332 = 8'ha4 == io_state_in_4 ? 8'ha0 : _GEN_7331; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7333 = 8'ha5 == io_state_in_4 ? 8'hab : _GEN_7332; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7334 = 8'ha6 == io_state_in_4 ? 8'hb6 : _GEN_7333; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7335 = 8'ha7 == io_state_in_4 ? 8'hbd : _GEN_7334; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7336 = 8'ha8 == io_state_in_4 ? 8'hd4 : _GEN_7335; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7337 = 8'ha9 == io_state_in_4 ? 8'hdf : _GEN_7336; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7338 = 8'haa == io_state_in_4 ? 8'hc2 : _GEN_7337; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7339 = 8'hab == io_state_in_4 ? 8'hc9 : _GEN_7338; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7340 = 8'hac == io_state_in_4 ? 8'hf8 : _GEN_7339; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7341 = 8'had == io_state_in_4 ? 8'hf3 : _GEN_7340; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7342 = 8'hae == io_state_in_4 ? 8'hee : _GEN_7341; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7343 = 8'haf == io_state_in_4 ? 8'he5 : _GEN_7342; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7344 = 8'hb0 == io_state_in_4 ? 8'h3c : _GEN_7343; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7345 = 8'hb1 == io_state_in_4 ? 8'h37 : _GEN_7344; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7346 = 8'hb2 == io_state_in_4 ? 8'h2a : _GEN_7345; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7347 = 8'hb3 == io_state_in_4 ? 8'h21 : _GEN_7346; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7348 = 8'hb4 == io_state_in_4 ? 8'h10 : _GEN_7347; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7349 = 8'hb5 == io_state_in_4 ? 8'h1b : _GEN_7348; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7350 = 8'hb6 == io_state_in_4 ? 8'h6 : _GEN_7349; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7351 = 8'hb7 == io_state_in_4 ? 8'hd : _GEN_7350; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7352 = 8'hb8 == io_state_in_4 ? 8'h64 : _GEN_7351; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7353 = 8'hb9 == io_state_in_4 ? 8'h6f : _GEN_7352; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7354 = 8'hba == io_state_in_4 ? 8'h72 : _GEN_7353; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7355 = 8'hbb == io_state_in_4 ? 8'h79 : _GEN_7354; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7356 = 8'hbc == io_state_in_4 ? 8'h48 : _GEN_7355; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7357 = 8'hbd == io_state_in_4 ? 8'h43 : _GEN_7356; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7358 = 8'hbe == io_state_in_4 ? 8'h5e : _GEN_7357; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7359 = 8'hbf == io_state_in_4 ? 8'h55 : _GEN_7358; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7360 = 8'hc0 == io_state_in_4 ? 8'h1 : _GEN_7359; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7361 = 8'hc1 == io_state_in_4 ? 8'ha : _GEN_7360; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7362 = 8'hc2 == io_state_in_4 ? 8'h17 : _GEN_7361; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7363 = 8'hc3 == io_state_in_4 ? 8'h1c : _GEN_7362; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7364 = 8'hc4 == io_state_in_4 ? 8'h2d : _GEN_7363; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7365 = 8'hc5 == io_state_in_4 ? 8'h26 : _GEN_7364; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7366 = 8'hc6 == io_state_in_4 ? 8'h3b : _GEN_7365; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7367 = 8'hc7 == io_state_in_4 ? 8'h30 : _GEN_7366; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7368 = 8'hc8 == io_state_in_4 ? 8'h59 : _GEN_7367; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7369 = 8'hc9 == io_state_in_4 ? 8'h52 : _GEN_7368; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7370 = 8'hca == io_state_in_4 ? 8'h4f : _GEN_7369; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7371 = 8'hcb == io_state_in_4 ? 8'h44 : _GEN_7370; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7372 = 8'hcc == io_state_in_4 ? 8'h75 : _GEN_7371; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7373 = 8'hcd == io_state_in_4 ? 8'h7e : _GEN_7372; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7374 = 8'hce == io_state_in_4 ? 8'h63 : _GEN_7373; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7375 = 8'hcf == io_state_in_4 ? 8'h68 : _GEN_7374; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7376 = 8'hd0 == io_state_in_4 ? 8'hb1 : _GEN_7375; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7377 = 8'hd1 == io_state_in_4 ? 8'hba : _GEN_7376; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7378 = 8'hd2 == io_state_in_4 ? 8'ha7 : _GEN_7377; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7379 = 8'hd3 == io_state_in_4 ? 8'hac : _GEN_7378; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7380 = 8'hd4 == io_state_in_4 ? 8'h9d : _GEN_7379; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7381 = 8'hd5 == io_state_in_4 ? 8'h96 : _GEN_7380; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7382 = 8'hd6 == io_state_in_4 ? 8'h8b : _GEN_7381; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7383 = 8'hd7 == io_state_in_4 ? 8'h80 : _GEN_7382; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7384 = 8'hd8 == io_state_in_4 ? 8'he9 : _GEN_7383; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7385 = 8'hd9 == io_state_in_4 ? 8'he2 : _GEN_7384; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7386 = 8'hda == io_state_in_4 ? 8'hff : _GEN_7385; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7387 = 8'hdb == io_state_in_4 ? 8'hf4 : _GEN_7386; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7388 = 8'hdc == io_state_in_4 ? 8'hc5 : _GEN_7387; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7389 = 8'hdd == io_state_in_4 ? 8'hce : _GEN_7388; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7390 = 8'hde == io_state_in_4 ? 8'hd3 : _GEN_7389; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7391 = 8'hdf == io_state_in_4 ? 8'hd8 : _GEN_7390; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7392 = 8'he0 == io_state_in_4 ? 8'h7a : _GEN_7391; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7393 = 8'he1 == io_state_in_4 ? 8'h71 : _GEN_7392; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7394 = 8'he2 == io_state_in_4 ? 8'h6c : _GEN_7393; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7395 = 8'he3 == io_state_in_4 ? 8'h67 : _GEN_7394; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7396 = 8'he4 == io_state_in_4 ? 8'h56 : _GEN_7395; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7397 = 8'he5 == io_state_in_4 ? 8'h5d : _GEN_7396; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7398 = 8'he6 == io_state_in_4 ? 8'h40 : _GEN_7397; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7399 = 8'he7 == io_state_in_4 ? 8'h4b : _GEN_7398; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7400 = 8'he8 == io_state_in_4 ? 8'h22 : _GEN_7399; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7401 = 8'he9 == io_state_in_4 ? 8'h29 : _GEN_7400; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7402 = 8'hea == io_state_in_4 ? 8'h34 : _GEN_7401; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7403 = 8'heb == io_state_in_4 ? 8'h3f : _GEN_7402; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7404 = 8'hec == io_state_in_4 ? 8'he : _GEN_7403; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7405 = 8'hed == io_state_in_4 ? 8'h5 : _GEN_7404; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7406 = 8'hee == io_state_in_4 ? 8'h18 : _GEN_7405; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7407 = 8'hef == io_state_in_4 ? 8'h13 : _GEN_7406; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7408 = 8'hf0 == io_state_in_4 ? 8'hca : _GEN_7407; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7409 = 8'hf1 == io_state_in_4 ? 8'hc1 : _GEN_7408; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7410 = 8'hf2 == io_state_in_4 ? 8'hdc : _GEN_7409; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7411 = 8'hf3 == io_state_in_4 ? 8'hd7 : _GEN_7410; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7412 = 8'hf4 == io_state_in_4 ? 8'he6 : _GEN_7411; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7413 = 8'hf5 == io_state_in_4 ? 8'hed : _GEN_7412; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7414 = 8'hf6 == io_state_in_4 ? 8'hf0 : _GEN_7413; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7415 = 8'hf7 == io_state_in_4 ? 8'hfb : _GEN_7414; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7416 = 8'hf8 == io_state_in_4 ? 8'h92 : _GEN_7415; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7417 = 8'hf9 == io_state_in_4 ? 8'h99 : _GEN_7416; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7418 = 8'hfa == io_state_in_4 ? 8'h84 : _GEN_7417; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7419 = 8'hfb == io_state_in_4 ? 8'h8f : _GEN_7418; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7420 = 8'hfc == io_state_in_4 ? 8'hbe : _GEN_7419; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7421 = 8'hfd == io_state_in_4 ? 8'hb5 : _GEN_7420; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7422 = 8'hfe == io_state_in_4 ? 8'ha8 : _GEN_7421; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7423 = 8'hff == io_state_in_4 ? 8'ha3 : _GEN_7422; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7425 = 8'h1 == io_state_in_5 ? 8'hd : 8'h0; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7426 = 8'h2 == io_state_in_5 ? 8'h1a : _GEN_7425; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7427 = 8'h3 == io_state_in_5 ? 8'h17 : _GEN_7426; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7428 = 8'h4 == io_state_in_5 ? 8'h34 : _GEN_7427; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7429 = 8'h5 == io_state_in_5 ? 8'h39 : _GEN_7428; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7430 = 8'h6 == io_state_in_5 ? 8'h2e : _GEN_7429; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7431 = 8'h7 == io_state_in_5 ? 8'h23 : _GEN_7430; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7432 = 8'h8 == io_state_in_5 ? 8'h68 : _GEN_7431; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7433 = 8'h9 == io_state_in_5 ? 8'h65 : _GEN_7432; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7434 = 8'ha == io_state_in_5 ? 8'h72 : _GEN_7433; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7435 = 8'hb == io_state_in_5 ? 8'h7f : _GEN_7434; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7436 = 8'hc == io_state_in_5 ? 8'h5c : _GEN_7435; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7437 = 8'hd == io_state_in_5 ? 8'h51 : _GEN_7436; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7438 = 8'he == io_state_in_5 ? 8'h46 : _GEN_7437; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7439 = 8'hf == io_state_in_5 ? 8'h4b : _GEN_7438; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7440 = 8'h10 == io_state_in_5 ? 8'hd0 : _GEN_7439; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7441 = 8'h11 == io_state_in_5 ? 8'hdd : _GEN_7440; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7442 = 8'h12 == io_state_in_5 ? 8'hca : _GEN_7441; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7443 = 8'h13 == io_state_in_5 ? 8'hc7 : _GEN_7442; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7444 = 8'h14 == io_state_in_5 ? 8'he4 : _GEN_7443; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7445 = 8'h15 == io_state_in_5 ? 8'he9 : _GEN_7444; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7446 = 8'h16 == io_state_in_5 ? 8'hfe : _GEN_7445; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7447 = 8'h17 == io_state_in_5 ? 8'hf3 : _GEN_7446; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7448 = 8'h18 == io_state_in_5 ? 8'hb8 : _GEN_7447; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7449 = 8'h19 == io_state_in_5 ? 8'hb5 : _GEN_7448; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7450 = 8'h1a == io_state_in_5 ? 8'ha2 : _GEN_7449; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7451 = 8'h1b == io_state_in_5 ? 8'haf : _GEN_7450; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7452 = 8'h1c == io_state_in_5 ? 8'h8c : _GEN_7451; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7453 = 8'h1d == io_state_in_5 ? 8'h81 : _GEN_7452; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7454 = 8'h1e == io_state_in_5 ? 8'h96 : _GEN_7453; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7455 = 8'h1f == io_state_in_5 ? 8'h9b : _GEN_7454; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7456 = 8'h20 == io_state_in_5 ? 8'hbb : _GEN_7455; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7457 = 8'h21 == io_state_in_5 ? 8'hb6 : _GEN_7456; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7458 = 8'h22 == io_state_in_5 ? 8'ha1 : _GEN_7457; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7459 = 8'h23 == io_state_in_5 ? 8'hac : _GEN_7458; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7460 = 8'h24 == io_state_in_5 ? 8'h8f : _GEN_7459; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7461 = 8'h25 == io_state_in_5 ? 8'h82 : _GEN_7460; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7462 = 8'h26 == io_state_in_5 ? 8'h95 : _GEN_7461; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7463 = 8'h27 == io_state_in_5 ? 8'h98 : _GEN_7462; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7464 = 8'h28 == io_state_in_5 ? 8'hd3 : _GEN_7463; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7465 = 8'h29 == io_state_in_5 ? 8'hde : _GEN_7464; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7466 = 8'h2a == io_state_in_5 ? 8'hc9 : _GEN_7465; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7467 = 8'h2b == io_state_in_5 ? 8'hc4 : _GEN_7466; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7468 = 8'h2c == io_state_in_5 ? 8'he7 : _GEN_7467; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7469 = 8'h2d == io_state_in_5 ? 8'hea : _GEN_7468; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7470 = 8'h2e == io_state_in_5 ? 8'hfd : _GEN_7469; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7471 = 8'h2f == io_state_in_5 ? 8'hf0 : _GEN_7470; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7472 = 8'h30 == io_state_in_5 ? 8'h6b : _GEN_7471; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7473 = 8'h31 == io_state_in_5 ? 8'h66 : _GEN_7472; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7474 = 8'h32 == io_state_in_5 ? 8'h71 : _GEN_7473; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7475 = 8'h33 == io_state_in_5 ? 8'h7c : _GEN_7474; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7476 = 8'h34 == io_state_in_5 ? 8'h5f : _GEN_7475; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7477 = 8'h35 == io_state_in_5 ? 8'h52 : _GEN_7476; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7478 = 8'h36 == io_state_in_5 ? 8'h45 : _GEN_7477; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7479 = 8'h37 == io_state_in_5 ? 8'h48 : _GEN_7478; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7480 = 8'h38 == io_state_in_5 ? 8'h3 : _GEN_7479; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7481 = 8'h39 == io_state_in_5 ? 8'he : _GEN_7480; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7482 = 8'h3a == io_state_in_5 ? 8'h19 : _GEN_7481; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7483 = 8'h3b == io_state_in_5 ? 8'h14 : _GEN_7482; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7484 = 8'h3c == io_state_in_5 ? 8'h37 : _GEN_7483; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7485 = 8'h3d == io_state_in_5 ? 8'h3a : _GEN_7484; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7486 = 8'h3e == io_state_in_5 ? 8'h2d : _GEN_7485; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7487 = 8'h3f == io_state_in_5 ? 8'h20 : _GEN_7486; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7488 = 8'h40 == io_state_in_5 ? 8'h6d : _GEN_7487; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7489 = 8'h41 == io_state_in_5 ? 8'h60 : _GEN_7488; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7490 = 8'h42 == io_state_in_5 ? 8'h77 : _GEN_7489; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7491 = 8'h43 == io_state_in_5 ? 8'h7a : _GEN_7490; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7492 = 8'h44 == io_state_in_5 ? 8'h59 : _GEN_7491; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7493 = 8'h45 == io_state_in_5 ? 8'h54 : _GEN_7492; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7494 = 8'h46 == io_state_in_5 ? 8'h43 : _GEN_7493; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7495 = 8'h47 == io_state_in_5 ? 8'h4e : _GEN_7494; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7496 = 8'h48 == io_state_in_5 ? 8'h5 : _GEN_7495; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7497 = 8'h49 == io_state_in_5 ? 8'h8 : _GEN_7496; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7498 = 8'h4a == io_state_in_5 ? 8'h1f : _GEN_7497; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7499 = 8'h4b == io_state_in_5 ? 8'h12 : _GEN_7498; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7500 = 8'h4c == io_state_in_5 ? 8'h31 : _GEN_7499; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7501 = 8'h4d == io_state_in_5 ? 8'h3c : _GEN_7500; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7502 = 8'h4e == io_state_in_5 ? 8'h2b : _GEN_7501; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7503 = 8'h4f == io_state_in_5 ? 8'h26 : _GEN_7502; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7504 = 8'h50 == io_state_in_5 ? 8'hbd : _GEN_7503; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7505 = 8'h51 == io_state_in_5 ? 8'hb0 : _GEN_7504; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7506 = 8'h52 == io_state_in_5 ? 8'ha7 : _GEN_7505; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7507 = 8'h53 == io_state_in_5 ? 8'haa : _GEN_7506; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7508 = 8'h54 == io_state_in_5 ? 8'h89 : _GEN_7507; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7509 = 8'h55 == io_state_in_5 ? 8'h84 : _GEN_7508; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7510 = 8'h56 == io_state_in_5 ? 8'h93 : _GEN_7509; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7511 = 8'h57 == io_state_in_5 ? 8'h9e : _GEN_7510; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7512 = 8'h58 == io_state_in_5 ? 8'hd5 : _GEN_7511; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7513 = 8'h59 == io_state_in_5 ? 8'hd8 : _GEN_7512; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7514 = 8'h5a == io_state_in_5 ? 8'hcf : _GEN_7513; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7515 = 8'h5b == io_state_in_5 ? 8'hc2 : _GEN_7514; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7516 = 8'h5c == io_state_in_5 ? 8'he1 : _GEN_7515; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7517 = 8'h5d == io_state_in_5 ? 8'hec : _GEN_7516; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7518 = 8'h5e == io_state_in_5 ? 8'hfb : _GEN_7517; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7519 = 8'h5f == io_state_in_5 ? 8'hf6 : _GEN_7518; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7520 = 8'h60 == io_state_in_5 ? 8'hd6 : _GEN_7519; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7521 = 8'h61 == io_state_in_5 ? 8'hdb : _GEN_7520; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7522 = 8'h62 == io_state_in_5 ? 8'hcc : _GEN_7521; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7523 = 8'h63 == io_state_in_5 ? 8'hc1 : _GEN_7522; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7524 = 8'h64 == io_state_in_5 ? 8'he2 : _GEN_7523; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7525 = 8'h65 == io_state_in_5 ? 8'hef : _GEN_7524; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7526 = 8'h66 == io_state_in_5 ? 8'hf8 : _GEN_7525; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7527 = 8'h67 == io_state_in_5 ? 8'hf5 : _GEN_7526; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7528 = 8'h68 == io_state_in_5 ? 8'hbe : _GEN_7527; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7529 = 8'h69 == io_state_in_5 ? 8'hb3 : _GEN_7528; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7530 = 8'h6a == io_state_in_5 ? 8'ha4 : _GEN_7529; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7531 = 8'h6b == io_state_in_5 ? 8'ha9 : _GEN_7530; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7532 = 8'h6c == io_state_in_5 ? 8'h8a : _GEN_7531; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7533 = 8'h6d == io_state_in_5 ? 8'h87 : _GEN_7532; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7534 = 8'h6e == io_state_in_5 ? 8'h90 : _GEN_7533; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7535 = 8'h6f == io_state_in_5 ? 8'h9d : _GEN_7534; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7536 = 8'h70 == io_state_in_5 ? 8'h6 : _GEN_7535; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7537 = 8'h71 == io_state_in_5 ? 8'hb : _GEN_7536; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7538 = 8'h72 == io_state_in_5 ? 8'h1c : _GEN_7537; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7539 = 8'h73 == io_state_in_5 ? 8'h11 : _GEN_7538; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7540 = 8'h74 == io_state_in_5 ? 8'h32 : _GEN_7539; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7541 = 8'h75 == io_state_in_5 ? 8'h3f : _GEN_7540; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7542 = 8'h76 == io_state_in_5 ? 8'h28 : _GEN_7541; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7543 = 8'h77 == io_state_in_5 ? 8'h25 : _GEN_7542; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7544 = 8'h78 == io_state_in_5 ? 8'h6e : _GEN_7543; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7545 = 8'h79 == io_state_in_5 ? 8'h63 : _GEN_7544; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7546 = 8'h7a == io_state_in_5 ? 8'h74 : _GEN_7545; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7547 = 8'h7b == io_state_in_5 ? 8'h79 : _GEN_7546; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7548 = 8'h7c == io_state_in_5 ? 8'h5a : _GEN_7547; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7549 = 8'h7d == io_state_in_5 ? 8'h57 : _GEN_7548; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7550 = 8'h7e == io_state_in_5 ? 8'h40 : _GEN_7549; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7551 = 8'h7f == io_state_in_5 ? 8'h4d : _GEN_7550; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7552 = 8'h80 == io_state_in_5 ? 8'hda : _GEN_7551; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7553 = 8'h81 == io_state_in_5 ? 8'hd7 : _GEN_7552; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7554 = 8'h82 == io_state_in_5 ? 8'hc0 : _GEN_7553; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7555 = 8'h83 == io_state_in_5 ? 8'hcd : _GEN_7554; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7556 = 8'h84 == io_state_in_5 ? 8'hee : _GEN_7555; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7557 = 8'h85 == io_state_in_5 ? 8'he3 : _GEN_7556; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7558 = 8'h86 == io_state_in_5 ? 8'hf4 : _GEN_7557; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7559 = 8'h87 == io_state_in_5 ? 8'hf9 : _GEN_7558; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7560 = 8'h88 == io_state_in_5 ? 8'hb2 : _GEN_7559; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7561 = 8'h89 == io_state_in_5 ? 8'hbf : _GEN_7560; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7562 = 8'h8a == io_state_in_5 ? 8'ha8 : _GEN_7561; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7563 = 8'h8b == io_state_in_5 ? 8'ha5 : _GEN_7562; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7564 = 8'h8c == io_state_in_5 ? 8'h86 : _GEN_7563; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7565 = 8'h8d == io_state_in_5 ? 8'h8b : _GEN_7564; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7566 = 8'h8e == io_state_in_5 ? 8'h9c : _GEN_7565; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7567 = 8'h8f == io_state_in_5 ? 8'h91 : _GEN_7566; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7568 = 8'h90 == io_state_in_5 ? 8'ha : _GEN_7567; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7569 = 8'h91 == io_state_in_5 ? 8'h7 : _GEN_7568; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7570 = 8'h92 == io_state_in_5 ? 8'h10 : _GEN_7569; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7571 = 8'h93 == io_state_in_5 ? 8'h1d : _GEN_7570; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7572 = 8'h94 == io_state_in_5 ? 8'h3e : _GEN_7571; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7573 = 8'h95 == io_state_in_5 ? 8'h33 : _GEN_7572; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7574 = 8'h96 == io_state_in_5 ? 8'h24 : _GEN_7573; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7575 = 8'h97 == io_state_in_5 ? 8'h29 : _GEN_7574; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7576 = 8'h98 == io_state_in_5 ? 8'h62 : _GEN_7575; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7577 = 8'h99 == io_state_in_5 ? 8'h6f : _GEN_7576; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7578 = 8'h9a == io_state_in_5 ? 8'h78 : _GEN_7577; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7579 = 8'h9b == io_state_in_5 ? 8'h75 : _GEN_7578; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7580 = 8'h9c == io_state_in_5 ? 8'h56 : _GEN_7579; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7581 = 8'h9d == io_state_in_5 ? 8'h5b : _GEN_7580; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7582 = 8'h9e == io_state_in_5 ? 8'h4c : _GEN_7581; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7583 = 8'h9f == io_state_in_5 ? 8'h41 : _GEN_7582; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7584 = 8'ha0 == io_state_in_5 ? 8'h61 : _GEN_7583; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7585 = 8'ha1 == io_state_in_5 ? 8'h6c : _GEN_7584; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7586 = 8'ha2 == io_state_in_5 ? 8'h7b : _GEN_7585; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7587 = 8'ha3 == io_state_in_5 ? 8'h76 : _GEN_7586; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7588 = 8'ha4 == io_state_in_5 ? 8'h55 : _GEN_7587; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7589 = 8'ha5 == io_state_in_5 ? 8'h58 : _GEN_7588; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7590 = 8'ha6 == io_state_in_5 ? 8'h4f : _GEN_7589; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7591 = 8'ha7 == io_state_in_5 ? 8'h42 : _GEN_7590; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7592 = 8'ha8 == io_state_in_5 ? 8'h9 : _GEN_7591; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7593 = 8'ha9 == io_state_in_5 ? 8'h4 : _GEN_7592; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7594 = 8'haa == io_state_in_5 ? 8'h13 : _GEN_7593; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7595 = 8'hab == io_state_in_5 ? 8'h1e : _GEN_7594; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7596 = 8'hac == io_state_in_5 ? 8'h3d : _GEN_7595; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7597 = 8'had == io_state_in_5 ? 8'h30 : _GEN_7596; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7598 = 8'hae == io_state_in_5 ? 8'h27 : _GEN_7597; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7599 = 8'haf == io_state_in_5 ? 8'h2a : _GEN_7598; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7600 = 8'hb0 == io_state_in_5 ? 8'hb1 : _GEN_7599; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7601 = 8'hb1 == io_state_in_5 ? 8'hbc : _GEN_7600; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7602 = 8'hb2 == io_state_in_5 ? 8'hab : _GEN_7601; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7603 = 8'hb3 == io_state_in_5 ? 8'ha6 : _GEN_7602; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7604 = 8'hb4 == io_state_in_5 ? 8'h85 : _GEN_7603; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7605 = 8'hb5 == io_state_in_5 ? 8'h88 : _GEN_7604; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7606 = 8'hb6 == io_state_in_5 ? 8'h9f : _GEN_7605; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7607 = 8'hb7 == io_state_in_5 ? 8'h92 : _GEN_7606; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7608 = 8'hb8 == io_state_in_5 ? 8'hd9 : _GEN_7607; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7609 = 8'hb9 == io_state_in_5 ? 8'hd4 : _GEN_7608; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7610 = 8'hba == io_state_in_5 ? 8'hc3 : _GEN_7609; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7611 = 8'hbb == io_state_in_5 ? 8'hce : _GEN_7610; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7612 = 8'hbc == io_state_in_5 ? 8'hed : _GEN_7611; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7613 = 8'hbd == io_state_in_5 ? 8'he0 : _GEN_7612; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7614 = 8'hbe == io_state_in_5 ? 8'hf7 : _GEN_7613; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7615 = 8'hbf == io_state_in_5 ? 8'hfa : _GEN_7614; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7616 = 8'hc0 == io_state_in_5 ? 8'hb7 : _GEN_7615; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7617 = 8'hc1 == io_state_in_5 ? 8'hba : _GEN_7616; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7618 = 8'hc2 == io_state_in_5 ? 8'had : _GEN_7617; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7619 = 8'hc3 == io_state_in_5 ? 8'ha0 : _GEN_7618; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7620 = 8'hc4 == io_state_in_5 ? 8'h83 : _GEN_7619; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7621 = 8'hc5 == io_state_in_5 ? 8'h8e : _GEN_7620; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7622 = 8'hc6 == io_state_in_5 ? 8'h99 : _GEN_7621; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7623 = 8'hc7 == io_state_in_5 ? 8'h94 : _GEN_7622; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7624 = 8'hc8 == io_state_in_5 ? 8'hdf : _GEN_7623; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7625 = 8'hc9 == io_state_in_5 ? 8'hd2 : _GEN_7624; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7626 = 8'hca == io_state_in_5 ? 8'hc5 : _GEN_7625; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7627 = 8'hcb == io_state_in_5 ? 8'hc8 : _GEN_7626; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7628 = 8'hcc == io_state_in_5 ? 8'heb : _GEN_7627; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7629 = 8'hcd == io_state_in_5 ? 8'he6 : _GEN_7628; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7630 = 8'hce == io_state_in_5 ? 8'hf1 : _GEN_7629; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7631 = 8'hcf == io_state_in_5 ? 8'hfc : _GEN_7630; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7632 = 8'hd0 == io_state_in_5 ? 8'h67 : _GEN_7631; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7633 = 8'hd1 == io_state_in_5 ? 8'h6a : _GEN_7632; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7634 = 8'hd2 == io_state_in_5 ? 8'h7d : _GEN_7633; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7635 = 8'hd3 == io_state_in_5 ? 8'h70 : _GEN_7634; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7636 = 8'hd4 == io_state_in_5 ? 8'h53 : _GEN_7635; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7637 = 8'hd5 == io_state_in_5 ? 8'h5e : _GEN_7636; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7638 = 8'hd6 == io_state_in_5 ? 8'h49 : _GEN_7637; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7639 = 8'hd7 == io_state_in_5 ? 8'h44 : _GEN_7638; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7640 = 8'hd8 == io_state_in_5 ? 8'hf : _GEN_7639; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7641 = 8'hd9 == io_state_in_5 ? 8'h2 : _GEN_7640; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7642 = 8'hda == io_state_in_5 ? 8'h15 : _GEN_7641; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7643 = 8'hdb == io_state_in_5 ? 8'h18 : _GEN_7642; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7644 = 8'hdc == io_state_in_5 ? 8'h3b : _GEN_7643; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7645 = 8'hdd == io_state_in_5 ? 8'h36 : _GEN_7644; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7646 = 8'hde == io_state_in_5 ? 8'h21 : _GEN_7645; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7647 = 8'hdf == io_state_in_5 ? 8'h2c : _GEN_7646; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7648 = 8'he0 == io_state_in_5 ? 8'hc : _GEN_7647; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7649 = 8'he1 == io_state_in_5 ? 8'h1 : _GEN_7648; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7650 = 8'he2 == io_state_in_5 ? 8'h16 : _GEN_7649; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7651 = 8'he3 == io_state_in_5 ? 8'h1b : _GEN_7650; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7652 = 8'he4 == io_state_in_5 ? 8'h38 : _GEN_7651; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7653 = 8'he5 == io_state_in_5 ? 8'h35 : _GEN_7652; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7654 = 8'he6 == io_state_in_5 ? 8'h22 : _GEN_7653; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7655 = 8'he7 == io_state_in_5 ? 8'h2f : _GEN_7654; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7656 = 8'he8 == io_state_in_5 ? 8'h64 : _GEN_7655; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7657 = 8'he9 == io_state_in_5 ? 8'h69 : _GEN_7656; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7658 = 8'hea == io_state_in_5 ? 8'h7e : _GEN_7657; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7659 = 8'heb == io_state_in_5 ? 8'h73 : _GEN_7658; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7660 = 8'hec == io_state_in_5 ? 8'h50 : _GEN_7659; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7661 = 8'hed == io_state_in_5 ? 8'h5d : _GEN_7660; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7662 = 8'hee == io_state_in_5 ? 8'h4a : _GEN_7661; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7663 = 8'hef == io_state_in_5 ? 8'h47 : _GEN_7662; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7664 = 8'hf0 == io_state_in_5 ? 8'hdc : _GEN_7663; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7665 = 8'hf1 == io_state_in_5 ? 8'hd1 : _GEN_7664; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7666 = 8'hf2 == io_state_in_5 ? 8'hc6 : _GEN_7665; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7667 = 8'hf3 == io_state_in_5 ? 8'hcb : _GEN_7666; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7668 = 8'hf4 == io_state_in_5 ? 8'he8 : _GEN_7667; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7669 = 8'hf5 == io_state_in_5 ? 8'he5 : _GEN_7668; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7670 = 8'hf6 == io_state_in_5 ? 8'hf2 : _GEN_7669; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7671 = 8'hf7 == io_state_in_5 ? 8'hff : _GEN_7670; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7672 = 8'hf8 == io_state_in_5 ? 8'hb4 : _GEN_7671; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7673 = 8'hf9 == io_state_in_5 ? 8'hb9 : _GEN_7672; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7674 = 8'hfa == io_state_in_5 ? 8'hae : _GEN_7673; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7675 = 8'hfb == io_state_in_5 ? 8'ha3 : _GEN_7674; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7676 = 8'hfc == io_state_in_5 ? 8'h80 : _GEN_7675; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7677 = 8'hfd == io_state_in_5 ? 8'h8d : _GEN_7676; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7678 = 8'hfe == io_state_in_5 ? 8'h9a : _GEN_7677; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _GEN_7679 = 8'hff == io_state_in_5 ? 8'h97 : _GEN_7678; // @[InvMixColumns.scala 134:{41,41}]
  wire [7:0] _tmp_state_7_T = _GEN_7423 ^ _GEN_7679; // @[InvMixColumns.scala 134:41]
  wire [7:0] _GEN_7681 = 8'h1 == io_state_in_6 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7682 = 8'h2 == io_state_in_6 ? 8'h12 : _GEN_7681; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7683 = 8'h3 == io_state_in_6 ? 8'h1b : _GEN_7682; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7684 = 8'h4 == io_state_in_6 ? 8'h24 : _GEN_7683; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7685 = 8'h5 == io_state_in_6 ? 8'h2d : _GEN_7684; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7686 = 8'h6 == io_state_in_6 ? 8'h36 : _GEN_7685; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7687 = 8'h7 == io_state_in_6 ? 8'h3f : _GEN_7686; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7688 = 8'h8 == io_state_in_6 ? 8'h48 : _GEN_7687; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7689 = 8'h9 == io_state_in_6 ? 8'h41 : _GEN_7688; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7690 = 8'ha == io_state_in_6 ? 8'h5a : _GEN_7689; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7691 = 8'hb == io_state_in_6 ? 8'h53 : _GEN_7690; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7692 = 8'hc == io_state_in_6 ? 8'h6c : _GEN_7691; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7693 = 8'hd == io_state_in_6 ? 8'h65 : _GEN_7692; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7694 = 8'he == io_state_in_6 ? 8'h7e : _GEN_7693; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7695 = 8'hf == io_state_in_6 ? 8'h77 : _GEN_7694; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7696 = 8'h10 == io_state_in_6 ? 8'h90 : _GEN_7695; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7697 = 8'h11 == io_state_in_6 ? 8'h99 : _GEN_7696; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7698 = 8'h12 == io_state_in_6 ? 8'h82 : _GEN_7697; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7699 = 8'h13 == io_state_in_6 ? 8'h8b : _GEN_7698; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7700 = 8'h14 == io_state_in_6 ? 8'hb4 : _GEN_7699; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7701 = 8'h15 == io_state_in_6 ? 8'hbd : _GEN_7700; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7702 = 8'h16 == io_state_in_6 ? 8'ha6 : _GEN_7701; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7703 = 8'h17 == io_state_in_6 ? 8'haf : _GEN_7702; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7704 = 8'h18 == io_state_in_6 ? 8'hd8 : _GEN_7703; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7705 = 8'h19 == io_state_in_6 ? 8'hd1 : _GEN_7704; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7706 = 8'h1a == io_state_in_6 ? 8'hca : _GEN_7705; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7707 = 8'h1b == io_state_in_6 ? 8'hc3 : _GEN_7706; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7708 = 8'h1c == io_state_in_6 ? 8'hfc : _GEN_7707; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7709 = 8'h1d == io_state_in_6 ? 8'hf5 : _GEN_7708; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7710 = 8'h1e == io_state_in_6 ? 8'hee : _GEN_7709; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7711 = 8'h1f == io_state_in_6 ? 8'he7 : _GEN_7710; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7712 = 8'h20 == io_state_in_6 ? 8'h3b : _GEN_7711; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7713 = 8'h21 == io_state_in_6 ? 8'h32 : _GEN_7712; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7714 = 8'h22 == io_state_in_6 ? 8'h29 : _GEN_7713; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7715 = 8'h23 == io_state_in_6 ? 8'h20 : _GEN_7714; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7716 = 8'h24 == io_state_in_6 ? 8'h1f : _GEN_7715; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7717 = 8'h25 == io_state_in_6 ? 8'h16 : _GEN_7716; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7718 = 8'h26 == io_state_in_6 ? 8'hd : _GEN_7717; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7719 = 8'h27 == io_state_in_6 ? 8'h4 : _GEN_7718; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7720 = 8'h28 == io_state_in_6 ? 8'h73 : _GEN_7719; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7721 = 8'h29 == io_state_in_6 ? 8'h7a : _GEN_7720; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7722 = 8'h2a == io_state_in_6 ? 8'h61 : _GEN_7721; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7723 = 8'h2b == io_state_in_6 ? 8'h68 : _GEN_7722; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7724 = 8'h2c == io_state_in_6 ? 8'h57 : _GEN_7723; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7725 = 8'h2d == io_state_in_6 ? 8'h5e : _GEN_7724; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7726 = 8'h2e == io_state_in_6 ? 8'h45 : _GEN_7725; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7727 = 8'h2f == io_state_in_6 ? 8'h4c : _GEN_7726; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7728 = 8'h30 == io_state_in_6 ? 8'hab : _GEN_7727; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7729 = 8'h31 == io_state_in_6 ? 8'ha2 : _GEN_7728; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7730 = 8'h32 == io_state_in_6 ? 8'hb9 : _GEN_7729; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7731 = 8'h33 == io_state_in_6 ? 8'hb0 : _GEN_7730; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7732 = 8'h34 == io_state_in_6 ? 8'h8f : _GEN_7731; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7733 = 8'h35 == io_state_in_6 ? 8'h86 : _GEN_7732; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7734 = 8'h36 == io_state_in_6 ? 8'h9d : _GEN_7733; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7735 = 8'h37 == io_state_in_6 ? 8'h94 : _GEN_7734; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7736 = 8'h38 == io_state_in_6 ? 8'he3 : _GEN_7735; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7737 = 8'h39 == io_state_in_6 ? 8'hea : _GEN_7736; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7738 = 8'h3a == io_state_in_6 ? 8'hf1 : _GEN_7737; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7739 = 8'h3b == io_state_in_6 ? 8'hf8 : _GEN_7738; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7740 = 8'h3c == io_state_in_6 ? 8'hc7 : _GEN_7739; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7741 = 8'h3d == io_state_in_6 ? 8'hce : _GEN_7740; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7742 = 8'h3e == io_state_in_6 ? 8'hd5 : _GEN_7741; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7743 = 8'h3f == io_state_in_6 ? 8'hdc : _GEN_7742; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7744 = 8'h40 == io_state_in_6 ? 8'h76 : _GEN_7743; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7745 = 8'h41 == io_state_in_6 ? 8'h7f : _GEN_7744; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7746 = 8'h42 == io_state_in_6 ? 8'h64 : _GEN_7745; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7747 = 8'h43 == io_state_in_6 ? 8'h6d : _GEN_7746; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7748 = 8'h44 == io_state_in_6 ? 8'h52 : _GEN_7747; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7749 = 8'h45 == io_state_in_6 ? 8'h5b : _GEN_7748; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7750 = 8'h46 == io_state_in_6 ? 8'h40 : _GEN_7749; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7751 = 8'h47 == io_state_in_6 ? 8'h49 : _GEN_7750; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7752 = 8'h48 == io_state_in_6 ? 8'h3e : _GEN_7751; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7753 = 8'h49 == io_state_in_6 ? 8'h37 : _GEN_7752; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7754 = 8'h4a == io_state_in_6 ? 8'h2c : _GEN_7753; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7755 = 8'h4b == io_state_in_6 ? 8'h25 : _GEN_7754; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7756 = 8'h4c == io_state_in_6 ? 8'h1a : _GEN_7755; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7757 = 8'h4d == io_state_in_6 ? 8'h13 : _GEN_7756; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7758 = 8'h4e == io_state_in_6 ? 8'h8 : _GEN_7757; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7759 = 8'h4f == io_state_in_6 ? 8'h1 : _GEN_7758; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7760 = 8'h50 == io_state_in_6 ? 8'he6 : _GEN_7759; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7761 = 8'h51 == io_state_in_6 ? 8'hef : _GEN_7760; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7762 = 8'h52 == io_state_in_6 ? 8'hf4 : _GEN_7761; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7763 = 8'h53 == io_state_in_6 ? 8'hfd : _GEN_7762; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7764 = 8'h54 == io_state_in_6 ? 8'hc2 : _GEN_7763; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7765 = 8'h55 == io_state_in_6 ? 8'hcb : _GEN_7764; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7766 = 8'h56 == io_state_in_6 ? 8'hd0 : _GEN_7765; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7767 = 8'h57 == io_state_in_6 ? 8'hd9 : _GEN_7766; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7768 = 8'h58 == io_state_in_6 ? 8'hae : _GEN_7767; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7769 = 8'h59 == io_state_in_6 ? 8'ha7 : _GEN_7768; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7770 = 8'h5a == io_state_in_6 ? 8'hbc : _GEN_7769; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7771 = 8'h5b == io_state_in_6 ? 8'hb5 : _GEN_7770; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7772 = 8'h5c == io_state_in_6 ? 8'h8a : _GEN_7771; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7773 = 8'h5d == io_state_in_6 ? 8'h83 : _GEN_7772; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7774 = 8'h5e == io_state_in_6 ? 8'h98 : _GEN_7773; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7775 = 8'h5f == io_state_in_6 ? 8'h91 : _GEN_7774; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7776 = 8'h60 == io_state_in_6 ? 8'h4d : _GEN_7775; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7777 = 8'h61 == io_state_in_6 ? 8'h44 : _GEN_7776; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7778 = 8'h62 == io_state_in_6 ? 8'h5f : _GEN_7777; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7779 = 8'h63 == io_state_in_6 ? 8'h56 : _GEN_7778; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7780 = 8'h64 == io_state_in_6 ? 8'h69 : _GEN_7779; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7781 = 8'h65 == io_state_in_6 ? 8'h60 : _GEN_7780; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7782 = 8'h66 == io_state_in_6 ? 8'h7b : _GEN_7781; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7783 = 8'h67 == io_state_in_6 ? 8'h72 : _GEN_7782; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7784 = 8'h68 == io_state_in_6 ? 8'h5 : _GEN_7783; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7785 = 8'h69 == io_state_in_6 ? 8'hc : _GEN_7784; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7786 = 8'h6a == io_state_in_6 ? 8'h17 : _GEN_7785; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7787 = 8'h6b == io_state_in_6 ? 8'h1e : _GEN_7786; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7788 = 8'h6c == io_state_in_6 ? 8'h21 : _GEN_7787; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7789 = 8'h6d == io_state_in_6 ? 8'h28 : _GEN_7788; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7790 = 8'h6e == io_state_in_6 ? 8'h33 : _GEN_7789; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7791 = 8'h6f == io_state_in_6 ? 8'h3a : _GEN_7790; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7792 = 8'h70 == io_state_in_6 ? 8'hdd : _GEN_7791; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7793 = 8'h71 == io_state_in_6 ? 8'hd4 : _GEN_7792; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7794 = 8'h72 == io_state_in_6 ? 8'hcf : _GEN_7793; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7795 = 8'h73 == io_state_in_6 ? 8'hc6 : _GEN_7794; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7796 = 8'h74 == io_state_in_6 ? 8'hf9 : _GEN_7795; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7797 = 8'h75 == io_state_in_6 ? 8'hf0 : _GEN_7796; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7798 = 8'h76 == io_state_in_6 ? 8'heb : _GEN_7797; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7799 = 8'h77 == io_state_in_6 ? 8'he2 : _GEN_7798; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7800 = 8'h78 == io_state_in_6 ? 8'h95 : _GEN_7799; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7801 = 8'h79 == io_state_in_6 ? 8'h9c : _GEN_7800; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7802 = 8'h7a == io_state_in_6 ? 8'h87 : _GEN_7801; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7803 = 8'h7b == io_state_in_6 ? 8'h8e : _GEN_7802; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7804 = 8'h7c == io_state_in_6 ? 8'hb1 : _GEN_7803; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7805 = 8'h7d == io_state_in_6 ? 8'hb8 : _GEN_7804; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7806 = 8'h7e == io_state_in_6 ? 8'ha3 : _GEN_7805; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7807 = 8'h7f == io_state_in_6 ? 8'haa : _GEN_7806; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7808 = 8'h80 == io_state_in_6 ? 8'hec : _GEN_7807; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7809 = 8'h81 == io_state_in_6 ? 8'he5 : _GEN_7808; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7810 = 8'h82 == io_state_in_6 ? 8'hfe : _GEN_7809; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7811 = 8'h83 == io_state_in_6 ? 8'hf7 : _GEN_7810; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7812 = 8'h84 == io_state_in_6 ? 8'hc8 : _GEN_7811; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7813 = 8'h85 == io_state_in_6 ? 8'hc1 : _GEN_7812; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7814 = 8'h86 == io_state_in_6 ? 8'hda : _GEN_7813; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7815 = 8'h87 == io_state_in_6 ? 8'hd3 : _GEN_7814; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7816 = 8'h88 == io_state_in_6 ? 8'ha4 : _GEN_7815; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7817 = 8'h89 == io_state_in_6 ? 8'had : _GEN_7816; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7818 = 8'h8a == io_state_in_6 ? 8'hb6 : _GEN_7817; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7819 = 8'h8b == io_state_in_6 ? 8'hbf : _GEN_7818; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7820 = 8'h8c == io_state_in_6 ? 8'h80 : _GEN_7819; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7821 = 8'h8d == io_state_in_6 ? 8'h89 : _GEN_7820; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7822 = 8'h8e == io_state_in_6 ? 8'h92 : _GEN_7821; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7823 = 8'h8f == io_state_in_6 ? 8'h9b : _GEN_7822; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7824 = 8'h90 == io_state_in_6 ? 8'h7c : _GEN_7823; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7825 = 8'h91 == io_state_in_6 ? 8'h75 : _GEN_7824; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7826 = 8'h92 == io_state_in_6 ? 8'h6e : _GEN_7825; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7827 = 8'h93 == io_state_in_6 ? 8'h67 : _GEN_7826; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7828 = 8'h94 == io_state_in_6 ? 8'h58 : _GEN_7827; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7829 = 8'h95 == io_state_in_6 ? 8'h51 : _GEN_7828; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7830 = 8'h96 == io_state_in_6 ? 8'h4a : _GEN_7829; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7831 = 8'h97 == io_state_in_6 ? 8'h43 : _GEN_7830; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7832 = 8'h98 == io_state_in_6 ? 8'h34 : _GEN_7831; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7833 = 8'h99 == io_state_in_6 ? 8'h3d : _GEN_7832; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7834 = 8'h9a == io_state_in_6 ? 8'h26 : _GEN_7833; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7835 = 8'h9b == io_state_in_6 ? 8'h2f : _GEN_7834; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7836 = 8'h9c == io_state_in_6 ? 8'h10 : _GEN_7835; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7837 = 8'h9d == io_state_in_6 ? 8'h19 : _GEN_7836; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7838 = 8'h9e == io_state_in_6 ? 8'h2 : _GEN_7837; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7839 = 8'h9f == io_state_in_6 ? 8'hb : _GEN_7838; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7840 = 8'ha0 == io_state_in_6 ? 8'hd7 : _GEN_7839; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7841 = 8'ha1 == io_state_in_6 ? 8'hde : _GEN_7840; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7842 = 8'ha2 == io_state_in_6 ? 8'hc5 : _GEN_7841; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7843 = 8'ha3 == io_state_in_6 ? 8'hcc : _GEN_7842; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7844 = 8'ha4 == io_state_in_6 ? 8'hf3 : _GEN_7843; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7845 = 8'ha5 == io_state_in_6 ? 8'hfa : _GEN_7844; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7846 = 8'ha6 == io_state_in_6 ? 8'he1 : _GEN_7845; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7847 = 8'ha7 == io_state_in_6 ? 8'he8 : _GEN_7846; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7848 = 8'ha8 == io_state_in_6 ? 8'h9f : _GEN_7847; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7849 = 8'ha9 == io_state_in_6 ? 8'h96 : _GEN_7848; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7850 = 8'haa == io_state_in_6 ? 8'h8d : _GEN_7849; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7851 = 8'hab == io_state_in_6 ? 8'h84 : _GEN_7850; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7852 = 8'hac == io_state_in_6 ? 8'hbb : _GEN_7851; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7853 = 8'had == io_state_in_6 ? 8'hb2 : _GEN_7852; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7854 = 8'hae == io_state_in_6 ? 8'ha9 : _GEN_7853; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7855 = 8'haf == io_state_in_6 ? 8'ha0 : _GEN_7854; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7856 = 8'hb0 == io_state_in_6 ? 8'h47 : _GEN_7855; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7857 = 8'hb1 == io_state_in_6 ? 8'h4e : _GEN_7856; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7858 = 8'hb2 == io_state_in_6 ? 8'h55 : _GEN_7857; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7859 = 8'hb3 == io_state_in_6 ? 8'h5c : _GEN_7858; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7860 = 8'hb4 == io_state_in_6 ? 8'h63 : _GEN_7859; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7861 = 8'hb5 == io_state_in_6 ? 8'h6a : _GEN_7860; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7862 = 8'hb6 == io_state_in_6 ? 8'h71 : _GEN_7861; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7863 = 8'hb7 == io_state_in_6 ? 8'h78 : _GEN_7862; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7864 = 8'hb8 == io_state_in_6 ? 8'hf : _GEN_7863; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7865 = 8'hb9 == io_state_in_6 ? 8'h6 : _GEN_7864; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7866 = 8'hba == io_state_in_6 ? 8'h1d : _GEN_7865; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7867 = 8'hbb == io_state_in_6 ? 8'h14 : _GEN_7866; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7868 = 8'hbc == io_state_in_6 ? 8'h2b : _GEN_7867; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7869 = 8'hbd == io_state_in_6 ? 8'h22 : _GEN_7868; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7870 = 8'hbe == io_state_in_6 ? 8'h39 : _GEN_7869; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7871 = 8'hbf == io_state_in_6 ? 8'h30 : _GEN_7870; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7872 = 8'hc0 == io_state_in_6 ? 8'h9a : _GEN_7871; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7873 = 8'hc1 == io_state_in_6 ? 8'h93 : _GEN_7872; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7874 = 8'hc2 == io_state_in_6 ? 8'h88 : _GEN_7873; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7875 = 8'hc3 == io_state_in_6 ? 8'h81 : _GEN_7874; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7876 = 8'hc4 == io_state_in_6 ? 8'hbe : _GEN_7875; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7877 = 8'hc5 == io_state_in_6 ? 8'hb7 : _GEN_7876; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7878 = 8'hc6 == io_state_in_6 ? 8'hac : _GEN_7877; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7879 = 8'hc7 == io_state_in_6 ? 8'ha5 : _GEN_7878; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7880 = 8'hc8 == io_state_in_6 ? 8'hd2 : _GEN_7879; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7881 = 8'hc9 == io_state_in_6 ? 8'hdb : _GEN_7880; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7882 = 8'hca == io_state_in_6 ? 8'hc0 : _GEN_7881; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7883 = 8'hcb == io_state_in_6 ? 8'hc9 : _GEN_7882; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7884 = 8'hcc == io_state_in_6 ? 8'hf6 : _GEN_7883; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7885 = 8'hcd == io_state_in_6 ? 8'hff : _GEN_7884; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7886 = 8'hce == io_state_in_6 ? 8'he4 : _GEN_7885; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7887 = 8'hcf == io_state_in_6 ? 8'hed : _GEN_7886; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7888 = 8'hd0 == io_state_in_6 ? 8'ha : _GEN_7887; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7889 = 8'hd1 == io_state_in_6 ? 8'h3 : _GEN_7888; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7890 = 8'hd2 == io_state_in_6 ? 8'h18 : _GEN_7889; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7891 = 8'hd3 == io_state_in_6 ? 8'h11 : _GEN_7890; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7892 = 8'hd4 == io_state_in_6 ? 8'h2e : _GEN_7891; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7893 = 8'hd5 == io_state_in_6 ? 8'h27 : _GEN_7892; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7894 = 8'hd6 == io_state_in_6 ? 8'h3c : _GEN_7893; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7895 = 8'hd7 == io_state_in_6 ? 8'h35 : _GEN_7894; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7896 = 8'hd8 == io_state_in_6 ? 8'h42 : _GEN_7895; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7897 = 8'hd9 == io_state_in_6 ? 8'h4b : _GEN_7896; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7898 = 8'hda == io_state_in_6 ? 8'h50 : _GEN_7897; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7899 = 8'hdb == io_state_in_6 ? 8'h59 : _GEN_7898; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7900 = 8'hdc == io_state_in_6 ? 8'h66 : _GEN_7899; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7901 = 8'hdd == io_state_in_6 ? 8'h6f : _GEN_7900; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7902 = 8'hde == io_state_in_6 ? 8'h74 : _GEN_7901; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7903 = 8'hdf == io_state_in_6 ? 8'h7d : _GEN_7902; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7904 = 8'he0 == io_state_in_6 ? 8'ha1 : _GEN_7903; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7905 = 8'he1 == io_state_in_6 ? 8'ha8 : _GEN_7904; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7906 = 8'he2 == io_state_in_6 ? 8'hb3 : _GEN_7905; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7907 = 8'he3 == io_state_in_6 ? 8'hba : _GEN_7906; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7908 = 8'he4 == io_state_in_6 ? 8'h85 : _GEN_7907; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7909 = 8'he5 == io_state_in_6 ? 8'h8c : _GEN_7908; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7910 = 8'he6 == io_state_in_6 ? 8'h97 : _GEN_7909; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7911 = 8'he7 == io_state_in_6 ? 8'h9e : _GEN_7910; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7912 = 8'he8 == io_state_in_6 ? 8'he9 : _GEN_7911; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7913 = 8'he9 == io_state_in_6 ? 8'he0 : _GEN_7912; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7914 = 8'hea == io_state_in_6 ? 8'hfb : _GEN_7913; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7915 = 8'heb == io_state_in_6 ? 8'hf2 : _GEN_7914; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7916 = 8'hec == io_state_in_6 ? 8'hcd : _GEN_7915; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7917 = 8'hed == io_state_in_6 ? 8'hc4 : _GEN_7916; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7918 = 8'hee == io_state_in_6 ? 8'hdf : _GEN_7917; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7919 = 8'hef == io_state_in_6 ? 8'hd6 : _GEN_7918; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7920 = 8'hf0 == io_state_in_6 ? 8'h31 : _GEN_7919; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7921 = 8'hf1 == io_state_in_6 ? 8'h38 : _GEN_7920; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7922 = 8'hf2 == io_state_in_6 ? 8'h23 : _GEN_7921; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7923 = 8'hf3 == io_state_in_6 ? 8'h2a : _GEN_7922; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7924 = 8'hf4 == io_state_in_6 ? 8'h15 : _GEN_7923; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7925 = 8'hf5 == io_state_in_6 ? 8'h1c : _GEN_7924; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7926 = 8'hf6 == io_state_in_6 ? 8'h7 : _GEN_7925; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7927 = 8'hf7 == io_state_in_6 ? 8'he : _GEN_7926; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7928 = 8'hf8 == io_state_in_6 ? 8'h79 : _GEN_7927; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7929 = 8'hf9 == io_state_in_6 ? 8'h70 : _GEN_7928; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7930 = 8'hfa == io_state_in_6 ? 8'h6b : _GEN_7929; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7931 = 8'hfb == io_state_in_6 ? 8'h62 : _GEN_7930; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7932 = 8'hfc == io_state_in_6 ? 8'h5d : _GEN_7931; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7933 = 8'hfd == io_state_in_6 ? 8'h54 : _GEN_7932; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7934 = 8'hfe == io_state_in_6 ? 8'h4f : _GEN_7933; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _GEN_7935 = 8'hff == io_state_in_6 ? 8'h46 : _GEN_7934; // @[InvMixColumns.scala 134:{65,65}]
  wire [7:0] _tmp_state_7_T_1 = _tmp_state_7_T ^ _GEN_7935; // @[InvMixColumns.scala 134:65]
  wire [7:0] _GEN_7937 = 8'h1 == io_state_in_7 ? 8'he : 8'h0; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7938 = 8'h2 == io_state_in_7 ? 8'h1c : _GEN_7937; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7939 = 8'h3 == io_state_in_7 ? 8'h12 : _GEN_7938; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7940 = 8'h4 == io_state_in_7 ? 8'h38 : _GEN_7939; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7941 = 8'h5 == io_state_in_7 ? 8'h36 : _GEN_7940; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7942 = 8'h6 == io_state_in_7 ? 8'h24 : _GEN_7941; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7943 = 8'h7 == io_state_in_7 ? 8'h2a : _GEN_7942; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7944 = 8'h8 == io_state_in_7 ? 8'h70 : _GEN_7943; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7945 = 8'h9 == io_state_in_7 ? 8'h7e : _GEN_7944; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7946 = 8'ha == io_state_in_7 ? 8'h6c : _GEN_7945; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7947 = 8'hb == io_state_in_7 ? 8'h62 : _GEN_7946; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7948 = 8'hc == io_state_in_7 ? 8'h48 : _GEN_7947; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7949 = 8'hd == io_state_in_7 ? 8'h46 : _GEN_7948; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7950 = 8'he == io_state_in_7 ? 8'h54 : _GEN_7949; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7951 = 8'hf == io_state_in_7 ? 8'h5a : _GEN_7950; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7952 = 8'h10 == io_state_in_7 ? 8'he0 : _GEN_7951; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7953 = 8'h11 == io_state_in_7 ? 8'hee : _GEN_7952; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7954 = 8'h12 == io_state_in_7 ? 8'hfc : _GEN_7953; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7955 = 8'h13 == io_state_in_7 ? 8'hf2 : _GEN_7954; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7956 = 8'h14 == io_state_in_7 ? 8'hd8 : _GEN_7955; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7957 = 8'h15 == io_state_in_7 ? 8'hd6 : _GEN_7956; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7958 = 8'h16 == io_state_in_7 ? 8'hc4 : _GEN_7957; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7959 = 8'h17 == io_state_in_7 ? 8'hca : _GEN_7958; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7960 = 8'h18 == io_state_in_7 ? 8'h90 : _GEN_7959; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7961 = 8'h19 == io_state_in_7 ? 8'h9e : _GEN_7960; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7962 = 8'h1a == io_state_in_7 ? 8'h8c : _GEN_7961; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7963 = 8'h1b == io_state_in_7 ? 8'h82 : _GEN_7962; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7964 = 8'h1c == io_state_in_7 ? 8'ha8 : _GEN_7963; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7965 = 8'h1d == io_state_in_7 ? 8'ha6 : _GEN_7964; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7966 = 8'h1e == io_state_in_7 ? 8'hb4 : _GEN_7965; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7967 = 8'h1f == io_state_in_7 ? 8'hba : _GEN_7966; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7968 = 8'h20 == io_state_in_7 ? 8'hdb : _GEN_7967; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7969 = 8'h21 == io_state_in_7 ? 8'hd5 : _GEN_7968; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7970 = 8'h22 == io_state_in_7 ? 8'hc7 : _GEN_7969; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7971 = 8'h23 == io_state_in_7 ? 8'hc9 : _GEN_7970; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7972 = 8'h24 == io_state_in_7 ? 8'he3 : _GEN_7971; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7973 = 8'h25 == io_state_in_7 ? 8'hed : _GEN_7972; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7974 = 8'h26 == io_state_in_7 ? 8'hff : _GEN_7973; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7975 = 8'h27 == io_state_in_7 ? 8'hf1 : _GEN_7974; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7976 = 8'h28 == io_state_in_7 ? 8'hab : _GEN_7975; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7977 = 8'h29 == io_state_in_7 ? 8'ha5 : _GEN_7976; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7978 = 8'h2a == io_state_in_7 ? 8'hb7 : _GEN_7977; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7979 = 8'h2b == io_state_in_7 ? 8'hb9 : _GEN_7978; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7980 = 8'h2c == io_state_in_7 ? 8'h93 : _GEN_7979; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7981 = 8'h2d == io_state_in_7 ? 8'h9d : _GEN_7980; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7982 = 8'h2e == io_state_in_7 ? 8'h8f : _GEN_7981; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7983 = 8'h2f == io_state_in_7 ? 8'h81 : _GEN_7982; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7984 = 8'h30 == io_state_in_7 ? 8'h3b : _GEN_7983; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7985 = 8'h31 == io_state_in_7 ? 8'h35 : _GEN_7984; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7986 = 8'h32 == io_state_in_7 ? 8'h27 : _GEN_7985; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7987 = 8'h33 == io_state_in_7 ? 8'h29 : _GEN_7986; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7988 = 8'h34 == io_state_in_7 ? 8'h3 : _GEN_7987; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7989 = 8'h35 == io_state_in_7 ? 8'hd : _GEN_7988; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7990 = 8'h36 == io_state_in_7 ? 8'h1f : _GEN_7989; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7991 = 8'h37 == io_state_in_7 ? 8'h11 : _GEN_7990; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7992 = 8'h38 == io_state_in_7 ? 8'h4b : _GEN_7991; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7993 = 8'h39 == io_state_in_7 ? 8'h45 : _GEN_7992; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7994 = 8'h3a == io_state_in_7 ? 8'h57 : _GEN_7993; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7995 = 8'h3b == io_state_in_7 ? 8'h59 : _GEN_7994; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7996 = 8'h3c == io_state_in_7 ? 8'h73 : _GEN_7995; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7997 = 8'h3d == io_state_in_7 ? 8'h7d : _GEN_7996; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7998 = 8'h3e == io_state_in_7 ? 8'h6f : _GEN_7997; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_7999 = 8'h3f == io_state_in_7 ? 8'h61 : _GEN_7998; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8000 = 8'h40 == io_state_in_7 ? 8'had : _GEN_7999; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8001 = 8'h41 == io_state_in_7 ? 8'ha3 : _GEN_8000; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8002 = 8'h42 == io_state_in_7 ? 8'hb1 : _GEN_8001; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8003 = 8'h43 == io_state_in_7 ? 8'hbf : _GEN_8002; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8004 = 8'h44 == io_state_in_7 ? 8'h95 : _GEN_8003; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8005 = 8'h45 == io_state_in_7 ? 8'h9b : _GEN_8004; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8006 = 8'h46 == io_state_in_7 ? 8'h89 : _GEN_8005; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8007 = 8'h47 == io_state_in_7 ? 8'h87 : _GEN_8006; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8008 = 8'h48 == io_state_in_7 ? 8'hdd : _GEN_8007; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8009 = 8'h49 == io_state_in_7 ? 8'hd3 : _GEN_8008; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8010 = 8'h4a == io_state_in_7 ? 8'hc1 : _GEN_8009; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8011 = 8'h4b == io_state_in_7 ? 8'hcf : _GEN_8010; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8012 = 8'h4c == io_state_in_7 ? 8'he5 : _GEN_8011; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8013 = 8'h4d == io_state_in_7 ? 8'heb : _GEN_8012; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8014 = 8'h4e == io_state_in_7 ? 8'hf9 : _GEN_8013; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8015 = 8'h4f == io_state_in_7 ? 8'hf7 : _GEN_8014; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8016 = 8'h50 == io_state_in_7 ? 8'h4d : _GEN_8015; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8017 = 8'h51 == io_state_in_7 ? 8'h43 : _GEN_8016; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8018 = 8'h52 == io_state_in_7 ? 8'h51 : _GEN_8017; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8019 = 8'h53 == io_state_in_7 ? 8'h5f : _GEN_8018; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8020 = 8'h54 == io_state_in_7 ? 8'h75 : _GEN_8019; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8021 = 8'h55 == io_state_in_7 ? 8'h7b : _GEN_8020; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8022 = 8'h56 == io_state_in_7 ? 8'h69 : _GEN_8021; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8023 = 8'h57 == io_state_in_7 ? 8'h67 : _GEN_8022; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8024 = 8'h58 == io_state_in_7 ? 8'h3d : _GEN_8023; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8025 = 8'h59 == io_state_in_7 ? 8'h33 : _GEN_8024; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8026 = 8'h5a == io_state_in_7 ? 8'h21 : _GEN_8025; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8027 = 8'h5b == io_state_in_7 ? 8'h2f : _GEN_8026; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8028 = 8'h5c == io_state_in_7 ? 8'h5 : _GEN_8027; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8029 = 8'h5d == io_state_in_7 ? 8'hb : _GEN_8028; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8030 = 8'h5e == io_state_in_7 ? 8'h19 : _GEN_8029; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8031 = 8'h5f == io_state_in_7 ? 8'h17 : _GEN_8030; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8032 = 8'h60 == io_state_in_7 ? 8'h76 : _GEN_8031; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8033 = 8'h61 == io_state_in_7 ? 8'h78 : _GEN_8032; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8034 = 8'h62 == io_state_in_7 ? 8'h6a : _GEN_8033; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8035 = 8'h63 == io_state_in_7 ? 8'h64 : _GEN_8034; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8036 = 8'h64 == io_state_in_7 ? 8'h4e : _GEN_8035; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8037 = 8'h65 == io_state_in_7 ? 8'h40 : _GEN_8036; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8038 = 8'h66 == io_state_in_7 ? 8'h52 : _GEN_8037; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8039 = 8'h67 == io_state_in_7 ? 8'h5c : _GEN_8038; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8040 = 8'h68 == io_state_in_7 ? 8'h6 : _GEN_8039; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8041 = 8'h69 == io_state_in_7 ? 8'h8 : _GEN_8040; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8042 = 8'h6a == io_state_in_7 ? 8'h1a : _GEN_8041; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8043 = 8'h6b == io_state_in_7 ? 8'h14 : _GEN_8042; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8044 = 8'h6c == io_state_in_7 ? 8'h3e : _GEN_8043; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8045 = 8'h6d == io_state_in_7 ? 8'h30 : _GEN_8044; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8046 = 8'h6e == io_state_in_7 ? 8'h22 : _GEN_8045; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8047 = 8'h6f == io_state_in_7 ? 8'h2c : _GEN_8046; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8048 = 8'h70 == io_state_in_7 ? 8'h96 : _GEN_8047; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8049 = 8'h71 == io_state_in_7 ? 8'h98 : _GEN_8048; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8050 = 8'h72 == io_state_in_7 ? 8'h8a : _GEN_8049; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8051 = 8'h73 == io_state_in_7 ? 8'h84 : _GEN_8050; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8052 = 8'h74 == io_state_in_7 ? 8'hae : _GEN_8051; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8053 = 8'h75 == io_state_in_7 ? 8'ha0 : _GEN_8052; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8054 = 8'h76 == io_state_in_7 ? 8'hb2 : _GEN_8053; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8055 = 8'h77 == io_state_in_7 ? 8'hbc : _GEN_8054; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8056 = 8'h78 == io_state_in_7 ? 8'he6 : _GEN_8055; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8057 = 8'h79 == io_state_in_7 ? 8'he8 : _GEN_8056; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8058 = 8'h7a == io_state_in_7 ? 8'hfa : _GEN_8057; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8059 = 8'h7b == io_state_in_7 ? 8'hf4 : _GEN_8058; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8060 = 8'h7c == io_state_in_7 ? 8'hde : _GEN_8059; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8061 = 8'h7d == io_state_in_7 ? 8'hd0 : _GEN_8060; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8062 = 8'h7e == io_state_in_7 ? 8'hc2 : _GEN_8061; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8063 = 8'h7f == io_state_in_7 ? 8'hcc : _GEN_8062; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8064 = 8'h80 == io_state_in_7 ? 8'h41 : _GEN_8063; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8065 = 8'h81 == io_state_in_7 ? 8'h4f : _GEN_8064; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8066 = 8'h82 == io_state_in_7 ? 8'h5d : _GEN_8065; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8067 = 8'h83 == io_state_in_7 ? 8'h53 : _GEN_8066; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8068 = 8'h84 == io_state_in_7 ? 8'h79 : _GEN_8067; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8069 = 8'h85 == io_state_in_7 ? 8'h77 : _GEN_8068; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8070 = 8'h86 == io_state_in_7 ? 8'h65 : _GEN_8069; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8071 = 8'h87 == io_state_in_7 ? 8'h6b : _GEN_8070; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8072 = 8'h88 == io_state_in_7 ? 8'h31 : _GEN_8071; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8073 = 8'h89 == io_state_in_7 ? 8'h3f : _GEN_8072; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8074 = 8'h8a == io_state_in_7 ? 8'h2d : _GEN_8073; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8075 = 8'h8b == io_state_in_7 ? 8'h23 : _GEN_8074; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8076 = 8'h8c == io_state_in_7 ? 8'h9 : _GEN_8075; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8077 = 8'h8d == io_state_in_7 ? 8'h7 : _GEN_8076; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8078 = 8'h8e == io_state_in_7 ? 8'h15 : _GEN_8077; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8079 = 8'h8f == io_state_in_7 ? 8'h1b : _GEN_8078; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8080 = 8'h90 == io_state_in_7 ? 8'ha1 : _GEN_8079; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8081 = 8'h91 == io_state_in_7 ? 8'haf : _GEN_8080; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8082 = 8'h92 == io_state_in_7 ? 8'hbd : _GEN_8081; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8083 = 8'h93 == io_state_in_7 ? 8'hb3 : _GEN_8082; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8084 = 8'h94 == io_state_in_7 ? 8'h99 : _GEN_8083; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8085 = 8'h95 == io_state_in_7 ? 8'h97 : _GEN_8084; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8086 = 8'h96 == io_state_in_7 ? 8'h85 : _GEN_8085; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8087 = 8'h97 == io_state_in_7 ? 8'h8b : _GEN_8086; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8088 = 8'h98 == io_state_in_7 ? 8'hd1 : _GEN_8087; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8089 = 8'h99 == io_state_in_7 ? 8'hdf : _GEN_8088; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8090 = 8'h9a == io_state_in_7 ? 8'hcd : _GEN_8089; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8091 = 8'h9b == io_state_in_7 ? 8'hc3 : _GEN_8090; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8092 = 8'h9c == io_state_in_7 ? 8'he9 : _GEN_8091; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8093 = 8'h9d == io_state_in_7 ? 8'he7 : _GEN_8092; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8094 = 8'h9e == io_state_in_7 ? 8'hf5 : _GEN_8093; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8095 = 8'h9f == io_state_in_7 ? 8'hfb : _GEN_8094; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8096 = 8'ha0 == io_state_in_7 ? 8'h9a : _GEN_8095; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8097 = 8'ha1 == io_state_in_7 ? 8'h94 : _GEN_8096; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8098 = 8'ha2 == io_state_in_7 ? 8'h86 : _GEN_8097; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8099 = 8'ha3 == io_state_in_7 ? 8'h88 : _GEN_8098; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8100 = 8'ha4 == io_state_in_7 ? 8'ha2 : _GEN_8099; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8101 = 8'ha5 == io_state_in_7 ? 8'hac : _GEN_8100; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8102 = 8'ha6 == io_state_in_7 ? 8'hbe : _GEN_8101; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8103 = 8'ha7 == io_state_in_7 ? 8'hb0 : _GEN_8102; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8104 = 8'ha8 == io_state_in_7 ? 8'hea : _GEN_8103; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8105 = 8'ha9 == io_state_in_7 ? 8'he4 : _GEN_8104; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8106 = 8'haa == io_state_in_7 ? 8'hf6 : _GEN_8105; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8107 = 8'hab == io_state_in_7 ? 8'hf8 : _GEN_8106; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8108 = 8'hac == io_state_in_7 ? 8'hd2 : _GEN_8107; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8109 = 8'had == io_state_in_7 ? 8'hdc : _GEN_8108; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8110 = 8'hae == io_state_in_7 ? 8'hce : _GEN_8109; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8111 = 8'haf == io_state_in_7 ? 8'hc0 : _GEN_8110; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8112 = 8'hb0 == io_state_in_7 ? 8'h7a : _GEN_8111; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8113 = 8'hb1 == io_state_in_7 ? 8'h74 : _GEN_8112; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8114 = 8'hb2 == io_state_in_7 ? 8'h66 : _GEN_8113; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8115 = 8'hb3 == io_state_in_7 ? 8'h68 : _GEN_8114; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8116 = 8'hb4 == io_state_in_7 ? 8'h42 : _GEN_8115; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8117 = 8'hb5 == io_state_in_7 ? 8'h4c : _GEN_8116; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8118 = 8'hb6 == io_state_in_7 ? 8'h5e : _GEN_8117; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8119 = 8'hb7 == io_state_in_7 ? 8'h50 : _GEN_8118; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8120 = 8'hb8 == io_state_in_7 ? 8'ha : _GEN_8119; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8121 = 8'hb9 == io_state_in_7 ? 8'h4 : _GEN_8120; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8122 = 8'hba == io_state_in_7 ? 8'h16 : _GEN_8121; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8123 = 8'hbb == io_state_in_7 ? 8'h18 : _GEN_8122; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8124 = 8'hbc == io_state_in_7 ? 8'h32 : _GEN_8123; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8125 = 8'hbd == io_state_in_7 ? 8'h3c : _GEN_8124; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8126 = 8'hbe == io_state_in_7 ? 8'h2e : _GEN_8125; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8127 = 8'hbf == io_state_in_7 ? 8'h20 : _GEN_8126; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8128 = 8'hc0 == io_state_in_7 ? 8'hec : _GEN_8127; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8129 = 8'hc1 == io_state_in_7 ? 8'he2 : _GEN_8128; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8130 = 8'hc2 == io_state_in_7 ? 8'hf0 : _GEN_8129; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8131 = 8'hc3 == io_state_in_7 ? 8'hfe : _GEN_8130; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8132 = 8'hc4 == io_state_in_7 ? 8'hd4 : _GEN_8131; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8133 = 8'hc5 == io_state_in_7 ? 8'hda : _GEN_8132; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8134 = 8'hc6 == io_state_in_7 ? 8'hc8 : _GEN_8133; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8135 = 8'hc7 == io_state_in_7 ? 8'hc6 : _GEN_8134; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8136 = 8'hc8 == io_state_in_7 ? 8'h9c : _GEN_8135; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8137 = 8'hc9 == io_state_in_7 ? 8'h92 : _GEN_8136; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8138 = 8'hca == io_state_in_7 ? 8'h80 : _GEN_8137; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8139 = 8'hcb == io_state_in_7 ? 8'h8e : _GEN_8138; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8140 = 8'hcc == io_state_in_7 ? 8'ha4 : _GEN_8139; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8141 = 8'hcd == io_state_in_7 ? 8'haa : _GEN_8140; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8142 = 8'hce == io_state_in_7 ? 8'hb8 : _GEN_8141; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8143 = 8'hcf == io_state_in_7 ? 8'hb6 : _GEN_8142; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8144 = 8'hd0 == io_state_in_7 ? 8'hc : _GEN_8143; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8145 = 8'hd1 == io_state_in_7 ? 8'h2 : _GEN_8144; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8146 = 8'hd2 == io_state_in_7 ? 8'h10 : _GEN_8145; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8147 = 8'hd3 == io_state_in_7 ? 8'h1e : _GEN_8146; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8148 = 8'hd4 == io_state_in_7 ? 8'h34 : _GEN_8147; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8149 = 8'hd5 == io_state_in_7 ? 8'h3a : _GEN_8148; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8150 = 8'hd6 == io_state_in_7 ? 8'h28 : _GEN_8149; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8151 = 8'hd7 == io_state_in_7 ? 8'h26 : _GEN_8150; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8152 = 8'hd8 == io_state_in_7 ? 8'h7c : _GEN_8151; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8153 = 8'hd9 == io_state_in_7 ? 8'h72 : _GEN_8152; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8154 = 8'hda == io_state_in_7 ? 8'h60 : _GEN_8153; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8155 = 8'hdb == io_state_in_7 ? 8'h6e : _GEN_8154; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8156 = 8'hdc == io_state_in_7 ? 8'h44 : _GEN_8155; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8157 = 8'hdd == io_state_in_7 ? 8'h4a : _GEN_8156; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8158 = 8'hde == io_state_in_7 ? 8'h58 : _GEN_8157; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8159 = 8'hdf == io_state_in_7 ? 8'h56 : _GEN_8158; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8160 = 8'he0 == io_state_in_7 ? 8'h37 : _GEN_8159; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8161 = 8'he1 == io_state_in_7 ? 8'h39 : _GEN_8160; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8162 = 8'he2 == io_state_in_7 ? 8'h2b : _GEN_8161; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8163 = 8'he3 == io_state_in_7 ? 8'h25 : _GEN_8162; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8164 = 8'he4 == io_state_in_7 ? 8'hf : _GEN_8163; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8165 = 8'he5 == io_state_in_7 ? 8'h1 : _GEN_8164; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8166 = 8'he6 == io_state_in_7 ? 8'h13 : _GEN_8165; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8167 = 8'he7 == io_state_in_7 ? 8'h1d : _GEN_8166; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8168 = 8'he8 == io_state_in_7 ? 8'h47 : _GEN_8167; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8169 = 8'he9 == io_state_in_7 ? 8'h49 : _GEN_8168; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8170 = 8'hea == io_state_in_7 ? 8'h5b : _GEN_8169; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8171 = 8'heb == io_state_in_7 ? 8'h55 : _GEN_8170; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8172 = 8'hec == io_state_in_7 ? 8'h7f : _GEN_8171; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8173 = 8'hed == io_state_in_7 ? 8'h71 : _GEN_8172; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8174 = 8'hee == io_state_in_7 ? 8'h63 : _GEN_8173; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8175 = 8'hef == io_state_in_7 ? 8'h6d : _GEN_8174; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8176 = 8'hf0 == io_state_in_7 ? 8'hd7 : _GEN_8175; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8177 = 8'hf1 == io_state_in_7 ? 8'hd9 : _GEN_8176; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8178 = 8'hf2 == io_state_in_7 ? 8'hcb : _GEN_8177; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8179 = 8'hf3 == io_state_in_7 ? 8'hc5 : _GEN_8178; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8180 = 8'hf4 == io_state_in_7 ? 8'hef : _GEN_8179; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8181 = 8'hf5 == io_state_in_7 ? 8'he1 : _GEN_8180; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8182 = 8'hf6 == io_state_in_7 ? 8'hf3 : _GEN_8181; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8183 = 8'hf7 == io_state_in_7 ? 8'hfd : _GEN_8182; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8184 = 8'hf8 == io_state_in_7 ? 8'ha7 : _GEN_8183; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8185 = 8'hf9 == io_state_in_7 ? 8'ha9 : _GEN_8184; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8186 = 8'hfa == io_state_in_7 ? 8'hbb : _GEN_8185; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8187 = 8'hfb == io_state_in_7 ? 8'hb5 : _GEN_8186; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8188 = 8'hfc == io_state_in_7 ? 8'h9f : _GEN_8187; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8189 = 8'hfd == io_state_in_7 ? 8'h91 : _GEN_8188; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8190 = 8'hfe == io_state_in_7 ? 8'h83 : _GEN_8189; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8191 = 8'hff == io_state_in_7 ? 8'h8d : _GEN_8190; // @[InvMixColumns.scala 134:{89,89}]
  wire [7:0] _GEN_8193 = 8'h1 == io_state_in_8 ? 8'he : 8'h0; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8194 = 8'h2 == io_state_in_8 ? 8'h1c : _GEN_8193; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8195 = 8'h3 == io_state_in_8 ? 8'h12 : _GEN_8194; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8196 = 8'h4 == io_state_in_8 ? 8'h38 : _GEN_8195; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8197 = 8'h5 == io_state_in_8 ? 8'h36 : _GEN_8196; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8198 = 8'h6 == io_state_in_8 ? 8'h24 : _GEN_8197; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8199 = 8'h7 == io_state_in_8 ? 8'h2a : _GEN_8198; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8200 = 8'h8 == io_state_in_8 ? 8'h70 : _GEN_8199; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8201 = 8'h9 == io_state_in_8 ? 8'h7e : _GEN_8200; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8202 = 8'ha == io_state_in_8 ? 8'h6c : _GEN_8201; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8203 = 8'hb == io_state_in_8 ? 8'h62 : _GEN_8202; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8204 = 8'hc == io_state_in_8 ? 8'h48 : _GEN_8203; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8205 = 8'hd == io_state_in_8 ? 8'h46 : _GEN_8204; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8206 = 8'he == io_state_in_8 ? 8'h54 : _GEN_8205; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8207 = 8'hf == io_state_in_8 ? 8'h5a : _GEN_8206; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8208 = 8'h10 == io_state_in_8 ? 8'he0 : _GEN_8207; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8209 = 8'h11 == io_state_in_8 ? 8'hee : _GEN_8208; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8210 = 8'h12 == io_state_in_8 ? 8'hfc : _GEN_8209; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8211 = 8'h13 == io_state_in_8 ? 8'hf2 : _GEN_8210; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8212 = 8'h14 == io_state_in_8 ? 8'hd8 : _GEN_8211; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8213 = 8'h15 == io_state_in_8 ? 8'hd6 : _GEN_8212; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8214 = 8'h16 == io_state_in_8 ? 8'hc4 : _GEN_8213; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8215 = 8'h17 == io_state_in_8 ? 8'hca : _GEN_8214; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8216 = 8'h18 == io_state_in_8 ? 8'h90 : _GEN_8215; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8217 = 8'h19 == io_state_in_8 ? 8'h9e : _GEN_8216; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8218 = 8'h1a == io_state_in_8 ? 8'h8c : _GEN_8217; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8219 = 8'h1b == io_state_in_8 ? 8'h82 : _GEN_8218; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8220 = 8'h1c == io_state_in_8 ? 8'ha8 : _GEN_8219; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8221 = 8'h1d == io_state_in_8 ? 8'ha6 : _GEN_8220; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8222 = 8'h1e == io_state_in_8 ? 8'hb4 : _GEN_8221; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8223 = 8'h1f == io_state_in_8 ? 8'hba : _GEN_8222; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8224 = 8'h20 == io_state_in_8 ? 8'hdb : _GEN_8223; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8225 = 8'h21 == io_state_in_8 ? 8'hd5 : _GEN_8224; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8226 = 8'h22 == io_state_in_8 ? 8'hc7 : _GEN_8225; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8227 = 8'h23 == io_state_in_8 ? 8'hc9 : _GEN_8226; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8228 = 8'h24 == io_state_in_8 ? 8'he3 : _GEN_8227; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8229 = 8'h25 == io_state_in_8 ? 8'hed : _GEN_8228; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8230 = 8'h26 == io_state_in_8 ? 8'hff : _GEN_8229; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8231 = 8'h27 == io_state_in_8 ? 8'hf1 : _GEN_8230; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8232 = 8'h28 == io_state_in_8 ? 8'hab : _GEN_8231; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8233 = 8'h29 == io_state_in_8 ? 8'ha5 : _GEN_8232; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8234 = 8'h2a == io_state_in_8 ? 8'hb7 : _GEN_8233; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8235 = 8'h2b == io_state_in_8 ? 8'hb9 : _GEN_8234; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8236 = 8'h2c == io_state_in_8 ? 8'h93 : _GEN_8235; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8237 = 8'h2d == io_state_in_8 ? 8'h9d : _GEN_8236; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8238 = 8'h2e == io_state_in_8 ? 8'h8f : _GEN_8237; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8239 = 8'h2f == io_state_in_8 ? 8'h81 : _GEN_8238; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8240 = 8'h30 == io_state_in_8 ? 8'h3b : _GEN_8239; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8241 = 8'h31 == io_state_in_8 ? 8'h35 : _GEN_8240; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8242 = 8'h32 == io_state_in_8 ? 8'h27 : _GEN_8241; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8243 = 8'h33 == io_state_in_8 ? 8'h29 : _GEN_8242; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8244 = 8'h34 == io_state_in_8 ? 8'h3 : _GEN_8243; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8245 = 8'h35 == io_state_in_8 ? 8'hd : _GEN_8244; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8246 = 8'h36 == io_state_in_8 ? 8'h1f : _GEN_8245; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8247 = 8'h37 == io_state_in_8 ? 8'h11 : _GEN_8246; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8248 = 8'h38 == io_state_in_8 ? 8'h4b : _GEN_8247; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8249 = 8'h39 == io_state_in_8 ? 8'h45 : _GEN_8248; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8250 = 8'h3a == io_state_in_8 ? 8'h57 : _GEN_8249; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8251 = 8'h3b == io_state_in_8 ? 8'h59 : _GEN_8250; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8252 = 8'h3c == io_state_in_8 ? 8'h73 : _GEN_8251; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8253 = 8'h3d == io_state_in_8 ? 8'h7d : _GEN_8252; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8254 = 8'h3e == io_state_in_8 ? 8'h6f : _GEN_8253; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8255 = 8'h3f == io_state_in_8 ? 8'h61 : _GEN_8254; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8256 = 8'h40 == io_state_in_8 ? 8'had : _GEN_8255; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8257 = 8'h41 == io_state_in_8 ? 8'ha3 : _GEN_8256; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8258 = 8'h42 == io_state_in_8 ? 8'hb1 : _GEN_8257; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8259 = 8'h43 == io_state_in_8 ? 8'hbf : _GEN_8258; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8260 = 8'h44 == io_state_in_8 ? 8'h95 : _GEN_8259; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8261 = 8'h45 == io_state_in_8 ? 8'h9b : _GEN_8260; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8262 = 8'h46 == io_state_in_8 ? 8'h89 : _GEN_8261; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8263 = 8'h47 == io_state_in_8 ? 8'h87 : _GEN_8262; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8264 = 8'h48 == io_state_in_8 ? 8'hdd : _GEN_8263; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8265 = 8'h49 == io_state_in_8 ? 8'hd3 : _GEN_8264; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8266 = 8'h4a == io_state_in_8 ? 8'hc1 : _GEN_8265; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8267 = 8'h4b == io_state_in_8 ? 8'hcf : _GEN_8266; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8268 = 8'h4c == io_state_in_8 ? 8'he5 : _GEN_8267; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8269 = 8'h4d == io_state_in_8 ? 8'heb : _GEN_8268; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8270 = 8'h4e == io_state_in_8 ? 8'hf9 : _GEN_8269; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8271 = 8'h4f == io_state_in_8 ? 8'hf7 : _GEN_8270; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8272 = 8'h50 == io_state_in_8 ? 8'h4d : _GEN_8271; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8273 = 8'h51 == io_state_in_8 ? 8'h43 : _GEN_8272; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8274 = 8'h52 == io_state_in_8 ? 8'h51 : _GEN_8273; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8275 = 8'h53 == io_state_in_8 ? 8'h5f : _GEN_8274; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8276 = 8'h54 == io_state_in_8 ? 8'h75 : _GEN_8275; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8277 = 8'h55 == io_state_in_8 ? 8'h7b : _GEN_8276; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8278 = 8'h56 == io_state_in_8 ? 8'h69 : _GEN_8277; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8279 = 8'h57 == io_state_in_8 ? 8'h67 : _GEN_8278; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8280 = 8'h58 == io_state_in_8 ? 8'h3d : _GEN_8279; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8281 = 8'h59 == io_state_in_8 ? 8'h33 : _GEN_8280; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8282 = 8'h5a == io_state_in_8 ? 8'h21 : _GEN_8281; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8283 = 8'h5b == io_state_in_8 ? 8'h2f : _GEN_8282; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8284 = 8'h5c == io_state_in_8 ? 8'h5 : _GEN_8283; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8285 = 8'h5d == io_state_in_8 ? 8'hb : _GEN_8284; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8286 = 8'h5e == io_state_in_8 ? 8'h19 : _GEN_8285; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8287 = 8'h5f == io_state_in_8 ? 8'h17 : _GEN_8286; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8288 = 8'h60 == io_state_in_8 ? 8'h76 : _GEN_8287; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8289 = 8'h61 == io_state_in_8 ? 8'h78 : _GEN_8288; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8290 = 8'h62 == io_state_in_8 ? 8'h6a : _GEN_8289; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8291 = 8'h63 == io_state_in_8 ? 8'h64 : _GEN_8290; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8292 = 8'h64 == io_state_in_8 ? 8'h4e : _GEN_8291; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8293 = 8'h65 == io_state_in_8 ? 8'h40 : _GEN_8292; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8294 = 8'h66 == io_state_in_8 ? 8'h52 : _GEN_8293; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8295 = 8'h67 == io_state_in_8 ? 8'h5c : _GEN_8294; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8296 = 8'h68 == io_state_in_8 ? 8'h6 : _GEN_8295; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8297 = 8'h69 == io_state_in_8 ? 8'h8 : _GEN_8296; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8298 = 8'h6a == io_state_in_8 ? 8'h1a : _GEN_8297; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8299 = 8'h6b == io_state_in_8 ? 8'h14 : _GEN_8298; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8300 = 8'h6c == io_state_in_8 ? 8'h3e : _GEN_8299; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8301 = 8'h6d == io_state_in_8 ? 8'h30 : _GEN_8300; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8302 = 8'h6e == io_state_in_8 ? 8'h22 : _GEN_8301; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8303 = 8'h6f == io_state_in_8 ? 8'h2c : _GEN_8302; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8304 = 8'h70 == io_state_in_8 ? 8'h96 : _GEN_8303; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8305 = 8'h71 == io_state_in_8 ? 8'h98 : _GEN_8304; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8306 = 8'h72 == io_state_in_8 ? 8'h8a : _GEN_8305; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8307 = 8'h73 == io_state_in_8 ? 8'h84 : _GEN_8306; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8308 = 8'h74 == io_state_in_8 ? 8'hae : _GEN_8307; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8309 = 8'h75 == io_state_in_8 ? 8'ha0 : _GEN_8308; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8310 = 8'h76 == io_state_in_8 ? 8'hb2 : _GEN_8309; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8311 = 8'h77 == io_state_in_8 ? 8'hbc : _GEN_8310; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8312 = 8'h78 == io_state_in_8 ? 8'he6 : _GEN_8311; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8313 = 8'h79 == io_state_in_8 ? 8'he8 : _GEN_8312; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8314 = 8'h7a == io_state_in_8 ? 8'hfa : _GEN_8313; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8315 = 8'h7b == io_state_in_8 ? 8'hf4 : _GEN_8314; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8316 = 8'h7c == io_state_in_8 ? 8'hde : _GEN_8315; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8317 = 8'h7d == io_state_in_8 ? 8'hd0 : _GEN_8316; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8318 = 8'h7e == io_state_in_8 ? 8'hc2 : _GEN_8317; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8319 = 8'h7f == io_state_in_8 ? 8'hcc : _GEN_8318; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8320 = 8'h80 == io_state_in_8 ? 8'h41 : _GEN_8319; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8321 = 8'h81 == io_state_in_8 ? 8'h4f : _GEN_8320; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8322 = 8'h82 == io_state_in_8 ? 8'h5d : _GEN_8321; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8323 = 8'h83 == io_state_in_8 ? 8'h53 : _GEN_8322; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8324 = 8'h84 == io_state_in_8 ? 8'h79 : _GEN_8323; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8325 = 8'h85 == io_state_in_8 ? 8'h77 : _GEN_8324; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8326 = 8'h86 == io_state_in_8 ? 8'h65 : _GEN_8325; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8327 = 8'h87 == io_state_in_8 ? 8'h6b : _GEN_8326; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8328 = 8'h88 == io_state_in_8 ? 8'h31 : _GEN_8327; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8329 = 8'h89 == io_state_in_8 ? 8'h3f : _GEN_8328; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8330 = 8'h8a == io_state_in_8 ? 8'h2d : _GEN_8329; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8331 = 8'h8b == io_state_in_8 ? 8'h23 : _GEN_8330; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8332 = 8'h8c == io_state_in_8 ? 8'h9 : _GEN_8331; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8333 = 8'h8d == io_state_in_8 ? 8'h7 : _GEN_8332; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8334 = 8'h8e == io_state_in_8 ? 8'h15 : _GEN_8333; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8335 = 8'h8f == io_state_in_8 ? 8'h1b : _GEN_8334; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8336 = 8'h90 == io_state_in_8 ? 8'ha1 : _GEN_8335; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8337 = 8'h91 == io_state_in_8 ? 8'haf : _GEN_8336; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8338 = 8'h92 == io_state_in_8 ? 8'hbd : _GEN_8337; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8339 = 8'h93 == io_state_in_8 ? 8'hb3 : _GEN_8338; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8340 = 8'h94 == io_state_in_8 ? 8'h99 : _GEN_8339; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8341 = 8'h95 == io_state_in_8 ? 8'h97 : _GEN_8340; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8342 = 8'h96 == io_state_in_8 ? 8'h85 : _GEN_8341; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8343 = 8'h97 == io_state_in_8 ? 8'h8b : _GEN_8342; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8344 = 8'h98 == io_state_in_8 ? 8'hd1 : _GEN_8343; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8345 = 8'h99 == io_state_in_8 ? 8'hdf : _GEN_8344; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8346 = 8'h9a == io_state_in_8 ? 8'hcd : _GEN_8345; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8347 = 8'h9b == io_state_in_8 ? 8'hc3 : _GEN_8346; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8348 = 8'h9c == io_state_in_8 ? 8'he9 : _GEN_8347; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8349 = 8'h9d == io_state_in_8 ? 8'he7 : _GEN_8348; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8350 = 8'h9e == io_state_in_8 ? 8'hf5 : _GEN_8349; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8351 = 8'h9f == io_state_in_8 ? 8'hfb : _GEN_8350; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8352 = 8'ha0 == io_state_in_8 ? 8'h9a : _GEN_8351; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8353 = 8'ha1 == io_state_in_8 ? 8'h94 : _GEN_8352; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8354 = 8'ha2 == io_state_in_8 ? 8'h86 : _GEN_8353; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8355 = 8'ha3 == io_state_in_8 ? 8'h88 : _GEN_8354; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8356 = 8'ha4 == io_state_in_8 ? 8'ha2 : _GEN_8355; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8357 = 8'ha5 == io_state_in_8 ? 8'hac : _GEN_8356; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8358 = 8'ha6 == io_state_in_8 ? 8'hbe : _GEN_8357; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8359 = 8'ha7 == io_state_in_8 ? 8'hb0 : _GEN_8358; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8360 = 8'ha8 == io_state_in_8 ? 8'hea : _GEN_8359; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8361 = 8'ha9 == io_state_in_8 ? 8'he4 : _GEN_8360; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8362 = 8'haa == io_state_in_8 ? 8'hf6 : _GEN_8361; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8363 = 8'hab == io_state_in_8 ? 8'hf8 : _GEN_8362; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8364 = 8'hac == io_state_in_8 ? 8'hd2 : _GEN_8363; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8365 = 8'had == io_state_in_8 ? 8'hdc : _GEN_8364; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8366 = 8'hae == io_state_in_8 ? 8'hce : _GEN_8365; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8367 = 8'haf == io_state_in_8 ? 8'hc0 : _GEN_8366; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8368 = 8'hb0 == io_state_in_8 ? 8'h7a : _GEN_8367; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8369 = 8'hb1 == io_state_in_8 ? 8'h74 : _GEN_8368; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8370 = 8'hb2 == io_state_in_8 ? 8'h66 : _GEN_8369; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8371 = 8'hb3 == io_state_in_8 ? 8'h68 : _GEN_8370; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8372 = 8'hb4 == io_state_in_8 ? 8'h42 : _GEN_8371; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8373 = 8'hb5 == io_state_in_8 ? 8'h4c : _GEN_8372; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8374 = 8'hb6 == io_state_in_8 ? 8'h5e : _GEN_8373; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8375 = 8'hb7 == io_state_in_8 ? 8'h50 : _GEN_8374; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8376 = 8'hb8 == io_state_in_8 ? 8'ha : _GEN_8375; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8377 = 8'hb9 == io_state_in_8 ? 8'h4 : _GEN_8376; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8378 = 8'hba == io_state_in_8 ? 8'h16 : _GEN_8377; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8379 = 8'hbb == io_state_in_8 ? 8'h18 : _GEN_8378; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8380 = 8'hbc == io_state_in_8 ? 8'h32 : _GEN_8379; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8381 = 8'hbd == io_state_in_8 ? 8'h3c : _GEN_8380; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8382 = 8'hbe == io_state_in_8 ? 8'h2e : _GEN_8381; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8383 = 8'hbf == io_state_in_8 ? 8'h20 : _GEN_8382; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8384 = 8'hc0 == io_state_in_8 ? 8'hec : _GEN_8383; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8385 = 8'hc1 == io_state_in_8 ? 8'he2 : _GEN_8384; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8386 = 8'hc2 == io_state_in_8 ? 8'hf0 : _GEN_8385; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8387 = 8'hc3 == io_state_in_8 ? 8'hfe : _GEN_8386; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8388 = 8'hc4 == io_state_in_8 ? 8'hd4 : _GEN_8387; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8389 = 8'hc5 == io_state_in_8 ? 8'hda : _GEN_8388; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8390 = 8'hc6 == io_state_in_8 ? 8'hc8 : _GEN_8389; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8391 = 8'hc7 == io_state_in_8 ? 8'hc6 : _GEN_8390; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8392 = 8'hc8 == io_state_in_8 ? 8'h9c : _GEN_8391; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8393 = 8'hc9 == io_state_in_8 ? 8'h92 : _GEN_8392; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8394 = 8'hca == io_state_in_8 ? 8'h80 : _GEN_8393; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8395 = 8'hcb == io_state_in_8 ? 8'h8e : _GEN_8394; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8396 = 8'hcc == io_state_in_8 ? 8'ha4 : _GEN_8395; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8397 = 8'hcd == io_state_in_8 ? 8'haa : _GEN_8396; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8398 = 8'hce == io_state_in_8 ? 8'hb8 : _GEN_8397; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8399 = 8'hcf == io_state_in_8 ? 8'hb6 : _GEN_8398; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8400 = 8'hd0 == io_state_in_8 ? 8'hc : _GEN_8399; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8401 = 8'hd1 == io_state_in_8 ? 8'h2 : _GEN_8400; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8402 = 8'hd2 == io_state_in_8 ? 8'h10 : _GEN_8401; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8403 = 8'hd3 == io_state_in_8 ? 8'h1e : _GEN_8402; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8404 = 8'hd4 == io_state_in_8 ? 8'h34 : _GEN_8403; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8405 = 8'hd5 == io_state_in_8 ? 8'h3a : _GEN_8404; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8406 = 8'hd6 == io_state_in_8 ? 8'h28 : _GEN_8405; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8407 = 8'hd7 == io_state_in_8 ? 8'h26 : _GEN_8406; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8408 = 8'hd8 == io_state_in_8 ? 8'h7c : _GEN_8407; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8409 = 8'hd9 == io_state_in_8 ? 8'h72 : _GEN_8408; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8410 = 8'hda == io_state_in_8 ? 8'h60 : _GEN_8409; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8411 = 8'hdb == io_state_in_8 ? 8'h6e : _GEN_8410; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8412 = 8'hdc == io_state_in_8 ? 8'h44 : _GEN_8411; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8413 = 8'hdd == io_state_in_8 ? 8'h4a : _GEN_8412; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8414 = 8'hde == io_state_in_8 ? 8'h58 : _GEN_8413; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8415 = 8'hdf == io_state_in_8 ? 8'h56 : _GEN_8414; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8416 = 8'he0 == io_state_in_8 ? 8'h37 : _GEN_8415; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8417 = 8'he1 == io_state_in_8 ? 8'h39 : _GEN_8416; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8418 = 8'he2 == io_state_in_8 ? 8'h2b : _GEN_8417; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8419 = 8'he3 == io_state_in_8 ? 8'h25 : _GEN_8418; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8420 = 8'he4 == io_state_in_8 ? 8'hf : _GEN_8419; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8421 = 8'he5 == io_state_in_8 ? 8'h1 : _GEN_8420; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8422 = 8'he6 == io_state_in_8 ? 8'h13 : _GEN_8421; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8423 = 8'he7 == io_state_in_8 ? 8'h1d : _GEN_8422; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8424 = 8'he8 == io_state_in_8 ? 8'h47 : _GEN_8423; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8425 = 8'he9 == io_state_in_8 ? 8'h49 : _GEN_8424; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8426 = 8'hea == io_state_in_8 ? 8'h5b : _GEN_8425; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8427 = 8'heb == io_state_in_8 ? 8'h55 : _GEN_8426; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8428 = 8'hec == io_state_in_8 ? 8'h7f : _GEN_8427; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8429 = 8'hed == io_state_in_8 ? 8'h71 : _GEN_8428; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8430 = 8'hee == io_state_in_8 ? 8'h63 : _GEN_8429; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8431 = 8'hef == io_state_in_8 ? 8'h6d : _GEN_8430; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8432 = 8'hf0 == io_state_in_8 ? 8'hd7 : _GEN_8431; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8433 = 8'hf1 == io_state_in_8 ? 8'hd9 : _GEN_8432; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8434 = 8'hf2 == io_state_in_8 ? 8'hcb : _GEN_8433; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8435 = 8'hf3 == io_state_in_8 ? 8'hc5 : _GEN_8434; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8436 = 8'hf4 == io_state_in_8 ? 8'hef : _GEN_8435; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8437 = 8'hf5 == io_state_in_8 ? 8'he1 : _GEN_8436; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8438 = 8'hf6 == io_state_in_8 ? 8'hf3 : _GEN_8437; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8439 = 8'hf7 == io_state_in_8 ? 8'hfd : _GEN_8438; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8440 = 8'hf8 == io_state_in_8 ? 8'ha7 : _GEN_8439; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8441 = 8'hf9 == io_state_in_8 ? 8'ha9 : _GEN_8440; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8442 = 8'hfa == io_state_in_8 ? 8'hbb : _GEN_8441; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8443 = 8'hfb == io_state_in_8 ? 8'hb5 : _GEN_8442; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8444 = 8'hfc == io_state_in_8 ? 8'h9f : _GEN_8443; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8445 = 8'hfd == io_state_in_8 ? 8'h91 : _GEN_8444; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8446 = 8'hfe == io_state_in_8 ? 8'h83 : _GEN_8445; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8447 = 8'hff == io_state_in_8 ? 8'h8d : _GEN_8446; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8449 = 8'h1 == io_state_in_9 ? 8'hb : 8'h0; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8450 = 8'h2 == io_state_in_9 ? 8'h16 : _GEN_8449; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8451 = 8'h3 == io_state_in_9 ? 8'h1d : _GEN_8450; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8452 = 8'h4 == io_state_in_9 ? 8'h2c : _GEN_8451; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8453 = 8'h5 == io_state_in_9 ? 8'h27 : _GEN_8452; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8454 = 8'h6 == io_state_in_9 ? 8'h3a : _GEN_8453; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8455 = 8'h7 == io_state_in_9 ? 8'h31 : _GEN_8454; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8456 = 8'h8 == io_state_in_9 ? 8'h58 : _GEN_8455; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8457 = 8'h9 == io_state_in_9 ? 8'h53 : _GEN_8456; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8458 = 8'ha == io_state_in_9 ? 8'h4e : _GEN_8457; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8459 = 8'hb == io_state_in_9 ? 8'h45 : _GEN_8458; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8460 = 8'hc == io_state_in_9 ? 8'h74 : _GEN_8459; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8461 = 8'hd == io_state_in_9 ? 8'h7f : _GEN_8460; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8462 = 8'he == io_state_in_9 ? 8'h62 : _GEN_8461; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8463 = 8'hf == io_state_in_9 ? 8'h69 : _GEN_8462; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8464 = 8'h10 == io_state_in_9 ? 8'hb0 : _GEN_8463; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8465 = 8'h11 == io_state_in_9 ? 8'hbb : _GEN_8464; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8466 = 8'h12 == io_state_in_9 ? 8'ha6 : _GEN_8465; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8467 = 8'h13 == io_state_in_9 ? 8'had : _GEN_8466; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8468 = 8'h14 == io_state_in_9 ? 8'h9c : _GEN_8467; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8469 = 8'h15 == io_state_in_9 ? 8'h97 : _GEN_8468; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8470 = 8'h16 == io_state_in_9 ? 8'h8a : _GEN_8469; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8471 = 8'h17 == io_state_in_9 ? 8'h81 : _GEN_8470; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8472 = 8'h18 == io_state_in_9 ? 8'he8 : _GEN_8471; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8473 = 8'h19 == io_state_in_9 ? 8'he3 : _GEN_8472; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8474 = 8'h1a == io_state_in_9 ? 8'hfe : _GEN_8473; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8475 = 8'h1b == io_state_in_9 ? 8'hf5 : _GEN_8474; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8476 = 8'h1c == io_state_in_9 ? 8'hc4 : _GEN_8475; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8477 = 8'h1d == io_state_in_9 ? 8'hcf : _GEN_8476; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8478 = 8'h1e == io_state_in_9 ? 8'hd2 : _GEN_8477; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8479 = 8'h1f == io_state_in_9 ? 8'hd9 : _GEN_8478; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8480 = 8'h20 == io_state_in_9 ? 8'h7b : _GEN_8479; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8481 = 8'h21 == io_state_in_9 ? 8'h70 : _GEN_8480; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8482 = 8'h22 == io_state_in_9 ? 8'h6d : _GEN_8481; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8483 = 8'h23 == io_state_in_9 ? 8'h66 : _GEN_8482; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8484 = 8'h24 == io_state_in_9 ? 8'h57 : _GEN_8483; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8485 = 8'h25 == io_state_in_9 ? 8'h5c : _GEN_8484; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8486 = 8'h26 == io_state_in_9 ? 8'h41 : _GEN_8485; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8487 = 8'h27 == io_state_in_9 ? 8'h4a : _GEN_8486; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8488 = 8'h28 == io_state_in_9 ? 8'h23 : _GEN_8487; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8489 = 8'h29 == io_state_in_9 ? 8'h28 : _GEN_8488; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8490 = 8'h2a == io_state_in_9 ? 8'h35 : _GEN_8489; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8491 = 8'h2b == io_state_in_9 ? 8'h3e : _GEN_8490; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8492 = 8'h2c == io_state_in_9 ? 8'hf : _GEN_8491; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8493 = 8'h2d == io_state_in_9 ? 8'h4 : _GEN_8492; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8494 = 8'h2e == io_state_in_9 ? 8'h19 : _GEN_8493; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8495 = 8'h2f == io_state_in_9 ? 8'h12 : _GEN_8494; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8496 = 8'h30 == io_state_in_9 ? 8'hcb : _GEN_8495; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8497 = 8'h31 == io_state_in_9 ? 8'hc0 : _GEN_8496; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8498 = 8'h32 == io_state_in_9 ? 8'hdd : _GEN_8497; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8499 = 8'h33 == io_state_in_9 ? 8'hd6 : _GEN_8498; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8500 = 8'h34 == io_state_in_9 ? 8'he7 : _GEN_8499; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8501 = 8'h35 == io_state_in_9 ? 8'hec : _GEN_8500; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8502 = 8'h36 == io_state_in_9 ? 8'hf1 : _GEN_8501; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8503 = 8'h37 == io_state_in_9 ? 8'hfa : _GEN_8502; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8504 = 8'h38 == io_state_in_9 ? 8'h93 : _GEN_8503; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8505 = 8'h39 == io_state_in_9 ? 8'h98 : _GEN_8504; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8506 = 8'h3a == io_state_in_9 ? 8'h85 : _GEN_8505; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8507 = 8'h3b == io_state_in_9 ? 8'h8e : _GEN_8506; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8508 = 8'h3c == io_state_in_9 ? 8'hbf : _GEN_8507; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8509 = 8'h3d == io_state_in_9 ? 8'hb4 : _GEN_8508; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8510 = 8'h3e == io_state_in_9 ? 8'ha9 : _GEN_8509; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8511 = 8'h3f == io_state_in_9 ? 8'ha2 : _GEN_8510; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8512 = 8'h40 == io_state_in_9 ? 8'hf6 : _GEN_8511; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8513 = 8'h41 == io_state_in_9 ? 8'hfd : _GEN_8512; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8514 = 8'h42 == io_state_in_9 ? 8'he0 : _GEN_8513; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8515 = 8'h43 == io_state_in_9 ? 8'heb : _GEN_8514; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8516 = 8'h44 == io_state_in_9 ? 8'hda : _GEN_8515; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8517 = 8'h45 == io_state_in_9 ? 8'hd1 : _GEN_8516; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8518 = 8'h46 == io_state_in_9 ? 8'hcc : _GEN_8517; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8519 = 8'h47 == io_state_in_9 ? 8'hc7 : _GEN_8518; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8520 = 8'h48 == io_state_in_9 ? 8'hae : _GEN_8519; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8521 = 8'h49 == io_state_in_9 ? 8'ha5 : _GEN_8520; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8522 = 8'h4a == io_state_in_9 ? 8'hb8 : _GEN_8521; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8523 = 8'h4b == io_state_in_9 ? 8'hb3 : _GEN_8522; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8524 = 8'h4c == io_state_in_9 ? 8'h82 : _GEN_8523; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8525 = 8'h4d == io_state_in_9 ? 8'h89 : _GEN_8524; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8526 = 8'h4e == io_state_in_9 ? 8'h94 : _GEN_8525; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8527 = 8'h4f == io_state_in_9 ? 8'h9f : _GEN_8526; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8528 = 8'h50 == io_state_in_9 ? 8'h46 : _GEN_8527; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8529 = 8'h51 == io_state_in_9 ? 8'h4d : _GEN_8528; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8530 = 8'h52 == io_state_in_9 ? 8'h50 : _GEN_8529; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8531 = 8'h53 == io_state_in_9 ? 8'h5b : _GEN_8530; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8532 = 8'h54 == io_state_in_9 ? 8'h6a : _GEN_8531; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8533 = 8'h55 == io_state_in_9 ? 8'h61 : _GEN_8532; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8534 = 8'h56 == io_state_in_9 ? 8'h7c : _GEN_8533; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8535 = 8'h57 == io_state_in_9 ? 8'h77 : _GEN_8534; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8536 = 8'h58 == io_state_in_9 ? 8'h1e : _GEN_8535; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8537 = 8'h59 == io_state_in_9 ? 8'h15 : _GEN_8536; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8538 = 8'h5a == io_state_in_9 ? 8'h8 : _GEN_8537; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8539 = 8'h5b == io_state_in_9 ? 8'h3 : _GEN_8538; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8540 = 8'h5c == io_state_in_9 ? 8'h32 : _GEN_8539; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8541 = 8'h5d == io_state_in_9 ? 8'h39 : _GEN_8540; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8542 = 8'h5e == io_state_in_9 ? 8'h24 : _GEN_8541; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8543 = 8'h5f == io_state_in_9 ? 8'h2f : _GEN_8542; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8544 = 8'h60 == io_state_in_9 ? 8'h8d : _GEN_8543; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8545 = 8'h61 == io_state_in_9 ? 8'h86 : _GEN_8544; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8546 = 8'h62 == io_state_in_9 ? 8'h9b : _GEN_8545; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8547 = 8'h63 == io_state_in_9 ? 8'h90 : _GEN_8546; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8548 = 8'h64 == io_state_in_9 ? 8'ha1 : _GEN_8547; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8549 = 8'h65 == io_state_in_9 ? 8'haa : _GEN_8548; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8550 = 8'h66 == io_state_in_9 ? 8'hb7 : _GEN_8549; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8551 = 8'h67 == io_state_in_9 ? 8'hbc : _GEN_8550; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8552 = 8'h68 == io_state_in_9 ? 8'hd5 : _GEN_8551; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8553 = 8'h69 == io_state_in_9 ? 8'hde : _GEN_8552; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8554 = 8'h6a == io_state_in_9 ? 8'hc3 : _GEN_8553; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8555 = 8'h6b == io_state_in_9 ? 8'hc8 : _GEN_8554; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8556 = 8'h6c == io_state_in_9 ? 8'hf9 : _GEN_8555; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8557 = 8'h6d == io_state_in_9 ? 8'hf2 : _GEN_8556; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8558 = 8'h6e == io_state_in_9 ? 8'hef : _GEN_8557; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8559 = 8'h6f == io_state_in_9 ? 8'he4 : _GEN_8558; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8560 = 8'h70 == io_state_in_9 ? 8'h3d : _GEN_8559; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8561 = 8'h71 == io_state_in_9 ? 8'h36 : _GEN_8560; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8562 = 8'h72 == io_state_in_9 ? 8'h2b : _GEN_8561; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8563 = 8'h73 == io_state_in_9 ? 8'h20 : _GEN_8562; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8564 = 8'h74 == io_state_in_9 ? 8'h11 : _GEN_8563; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8565 = 8'h75 == io_state_in_9 ? 8'h1a : _GEN_8564; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8566 = 8'h76 == io_state_in_9 ? 8'h7 : _GEN_8565; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8567 = 8'h77 == io_state_in_9 ? 8'hc : _GEN_8566; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8568 = 8'h78 == io_state_in_9 ? 8'h65 : _GEN_8567; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8569 = 8'h79 == io_state_in_9 ? 8'h6e : _GEN_8568; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8570 = 8'h7a == io_state_in_9 ? 8'h73 : _GEN_8569; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8571 = 8'h7b == io_state_in_9 ? 8'h78 : _GEN_8570; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8572 = 8'h7c == io_state_in_9 ? 8'h49 : _GEN_8571; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8573 = 8'h7d == io_state_in_9 ? 8'h42 : _GEN_8572; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8574 = 8'h7e == io_state_in_9 ? 8'h5f : _GEN_8573; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8575 = 8'h7f == io_state_in_9 ? 8'h54 : _GEN_8574; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8576 = 8'h80 == io_state_in_9 ? 8'hf7 : _GEN_8575; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8577 = 8'h81 == io_state_in_9 ? 8'hfc : _GEN_8576; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8578 = 8'h82 == io_state_in_9 ? 8'he1 : _GEN_8577; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8579 = 8'h83 == io_state_in_9 ? 8'hea : _GEN_8578; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8580 = 8'h84 == io_state_in_9 ? 8'hdb : _GEN_8579; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8581 = 8'h85 == io_state_in_9 ? 8'hd0 : _GEN_8580; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8582 = 8'h86 == io_state_in_9 ? 8'hcd : _GEN_8581; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8583 = 8'h87 == io_state_in_9 ? 8'hc6 : _GEN_8582; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8584 = 8'h88 == io_state_in_9 ? 8'haf : _GEN_8583; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8585 = 8'h89 == io_state_in_9 ? 8'ha4 : _GEN_8584; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8586 = 8'h8a == io_state_in_9 ? 8'hb9 : _GEN_8585; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8587 = 8'h8b == io_state_in_9 ? 8'hb2 : _GEN_8586; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8588 = 8'h8c == io_state_in_9 ? 8'h83 : _GEN_8587; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8589 = 8'h8d == io_state_in_9 ? 8'h88 : _GEN_8588; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8590 = 8'h8e == io_state_in_9 ? 8'h95 : _GEN_8589; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8591 = 8'h8f == io_state_in_9 ? 8'h9e : _GEN_8590; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8592 = 8'h90 == io_state_in_9 ? 8'h47 : _GEN_8591; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8593 = 8'h91 == io_state_in_9 ? 8'h4c : _GEN_8592; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8594 = 8'h92 == io_state_in_9 ? 8'h51 : _GEN_8593; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8595 = 8'h93 == io_state_in_9 ? 8'h5a : _GEN_8594; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8596 = 8'h94 == io_state_in_9 ? 8'h6b : _GEN_8595; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8597 = 8'h95 == io_state_in_9 ? 8'h60 : _GEN_8596; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8598 = 8'h96 == io_state_in_9 ? 8'h7d : _GEN_8597; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8599 = 8'h97 == io_state_in_9 ? 8'h76 : _GEN_8598; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8600 = 8'h98 == io_state_in_9 ? 8'h1f : _GEN_8599; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8601 = 8'h99 == io_state_in_9 ? 8'h14 : _GEN_8600; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8602 = 8'h9a == io_state_in_9 ? 8'h9 : _GEN_8601; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8603 = 8'h9b == io_state_in_9 ? 8'h2 : _GEN_8602; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8604 = 8'h9c == io_state_in_9 ? 8'h33 : _GEN_8603; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8605 = 8'h9d == io_state_in_9 ? 8'h38 : _GEN_8604; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8606 = 8'h9e == io_state_in_9 ? 8'h25 : _GEN_8605; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8607 = 8'h9f == io_state_in_9 ? 8'h2e : _GEN_8606; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8608 = 8'ha0 == io_state_in_9 ? 8'h8c : _GEN_8607; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8609 = 8'ha1 == io_state_in_9 ? 8'h87 : _GEN_8608; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8610 = 8'ha2 == io_state_in_9 ? 8'h9a : _GEN_8609; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8611 = 8'ha3 == io_state_in_9 ? 8'h91 : _GEN_8610; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8612 = 8'ha4 == io_state_in_9 ? 8'ha0 : _GEN_8611; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8613 = 8'ha5 == io_state_in_9 ? 8'hab : _GEN_8612; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8614 = 8'ha6 == io_state_in_9 ? 8'hb6 : _GEN_8613; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8615 = 8'ha7 == io_state_in_9 ? 8'hbd : _GEN_8614; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8616 = 8'ha8 == io_state_in_9 ? 8'hd4 : _GEN_8615; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8617 = 8'ha9 == io_state_in_9 ? 8'hdf : _GEN_8616; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8618 = 8'haa == io_state_in_9 ? 8'hc2 : _GEN_8617; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8619 = 8'hab == io_state_in_9 ? 8'hc9 : _GEN_8618; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8620 = 8'hac == io_state_in_9 ? 8'hf8 : _GEN_8619; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8621 = 8'had == io_state_in_9 ? 8'hf3 : _GEN_8620; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8622 = 8'hae == io_state_in_9 ? 8'hee : _GEN_8621; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8623 = 8'haf == io_state_in_9 ? 8'he5 : _GEN_8622; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8624 = 8'hb0 == io_state_in_9 ? 8'h3c : _GEN_8623; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8625 = 8'hb1 == io_state_in_9 ? 8'h37 : _GEN_8624; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8626 = 8'hb2 == io_state_in_9 ? 8'h2a : _GEN_8625; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8627 = 8'hb3 == io_state_in_9 ? 8'h21 : _GEN_8626; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8628 = 8'hb4 == io_state_in_9 ? 8'h10 : _GEN_8627; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8629 = 8'hb5 == io_state_in_9 ? 8'h1b : _GEN_8628; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8630 = 8'hb6 == io_state_in_9 ? 8'h6 : _GEN_8629; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8631 = 8'hb7 == io_state_in_9 ? 8'hd : _GEN_8630; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8632 = 8'hb8 == io_state_in_9 ? 8'h64 : _GEN_8631; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8633 = 8'hb9 == io_state_in_9 ? 8'h6f : _GEN_8632; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8634 = 8'hba == io_state_in_9 ? 8'h72 : _GEN_8633; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8635 = 8'hbb == io_state_in_9 ? 8'h79 : _GEN_8634; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8636 = 8'hbc == io_state_in_9 ? 8'h48 : _GEN_8635; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8637 = 8'hbd == io_state_in_9 ? 8'h43 : _GEN_8636; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8638 = 8'hbe == io_state_in_9 ? 8'h5e : _GEN_8637; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8639 = 8'hbf == io_state_in_9 ? 8'h55 : _GEN_8638; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8640 = 8'hc0 == io_state_in_9 ? 8'h1 : _GEN_8639; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8641 = 8'hc1 == io_state_in_9 ? 8'ha : _GEN_8640; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8642 = 8'hc2 == io_state_in_9 ? 8'h17 : _GEN_8641; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8643 = 8'hc3 == io_state_in_9 ? 8'h1c : _GEN_8642; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8644 = 8'hc4 == io_state_in_9 ? 8'h2d : _GEN_8643; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8645 = 8'hc5 == io_state_in_9 ? 8'h26 : _GEN_8644; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8646 = 8'hc6 == io_state_in_9 ? 8'h3b : _GEN_8645; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8647 = 8'hc7 == io_state_in_9 ? 8'h30 : _GEN_8646; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8648 = 8'hc8 == io_state_in_9 ? 8'h59 : _GEN_8647; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8649 = 8'hc9 == io_state_in_9 ? 8'h52 : _GEN_8648; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8650 = 8'hca == io_state_in_9 ? 8'h4f : _GEN_8649; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8651 = 8'hcb == io_state_in_9 ? 8'h44 : _GEN_8650; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8652 = 8'hcc == io_state_in_9 ? 8'h75 : _GEN_8651; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8653 = 8'hcd == io_state_in_9 ? 8'h7e : _GEN_8652; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8654 = 8'hce == io_state_in_9 ? 8'h63 : _GEN_8653; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8655 = 8'hcf == io_state_in_9 ? 8'h68 : _GEN_8654; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8656 = 8'hd0 == io_state_in_9 ? 8'hb1 : _GEN_8655; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8657 = 8'hd1 == io_state_in_9 ? 8'hba : _GEN_8656; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8658 = 8'hd2 == io_state_in_9 ? 8'ha7 : _GEN_8657; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8659 = 8'hd3 == io_state_in_9 ? 8'hac : _GEN_8658; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8660 = 8'hd4 == io_state_in_9 ? 8'h9d : _GEN_8659; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8661 = 8'hd5 == io_state_in_9 ? 8'h96 : _GEN_8660; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8662 = 8'hd6 == io_state_in_9 ? 8'h8b : _GEN_8661; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8663 = 8'hd7 == io_state_in_9 ? 8'h80 : _GEN_8662; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8664 = 8'hd8 == io_state_in_9 ? 8'he9 : _GEN_8663; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8665 = 8'hd9 == io_state_in_9 ? 8'he2 : _GEN_8664; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8666 = 8'hda == io_state_in_9 ? 8'hff : _GEN_8665; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8667 = 8'hdb == io_state_in_9 ? 8'hf4 : _GEN_8666; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8668 = 8'hdc == io_state_in_9 ? 8'hc5 : _GEN_8667; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8669 = 8'hdd == io_state_in_9 ? 8'hce : _GEN_8668; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8670 = 8'hde == io_state_in_9 ? 8'hd3 : _GEN_8669; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8671 = 8'hdf == io_state_in_9 ? 8'hd8 : _GEN_8670; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8672 = 8'he0 == io_state_in_9 ? 8'h7a : _GEN_8671; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8673 = 8'he1 == io_state_in_9 ? 8'h71 : _GEN_8672; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8674 = 8'he2 == io_state_in_9 ? 8'h6c : _GEN_8673; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8675 = 8'he3 == io_state_in_9 ? 8'h67 : _GEN_8674; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8676 = 8'he4 == io_state_in_9 ? 8'h56 : _GEN_8675; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8677 = 8'he5 == io_state_in_9 ? 8'h5d : _GEN_8676; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8678 = 8'he6 == io_state_in_9 ? 8'h40 : _GEN_8677; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8679 = 8'he7 == io_state_in_9 ? 8'h4b : _GEN_8678; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8680 = 8'he8 == io_state_in_9 ? 8'h22 : _GEN_8679; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8681 = 8'he9 == io_state_in_9 ? 8'h29 : _GEN_8680; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8682 = 8'hea == io_state_in_9 ? 8'h34 : _GEN_8681; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8683 = 8'heb == io_state_in_9 ? 8'h3f : _GEN_8682; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8684 = 8'hec == io_state_in_9 ? 8'he : _GEN_8683; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8685 = 8'hed == io_state_in_9 ? 8'h5 : _GEN_8684; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8686 = 8'hee == io_state_in_9 ? 8'h18 : _GEN_8685; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8687 = 8'hef == io_state_in_9 ? 8'h13 : _GEN_8686; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8688 = 8'hf0 == io_state_in_9 ? 8'hca : _GEN_8687; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8689 = 8'hf1 == io_state_in_9 ? 8'hc1 : _GEN_8688; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8690 = 8'hf2 == io_state_in_9 ? 8'hdc : _GEN_8689; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8691 = 8'hf3 == io_state_in_9 ? 8'hd7 : _GEN_8690; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8692 = 8'hf4 == io_state_in_9 ? 8'he6 : _GEN_8691; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8693 = 8'hf5 == io_state_in_9 ? 8'hed : _GEN_8692; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8694 = 8'hf6 == io_state_in_9 ? 8'hf0 : _GEN_8693; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8695 = 8'hf7 == io_state_in_9 ? 8'hfb : _GEN_8694; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8696 = 8'hf8 == io_state_in_9 ? 8'h92 : _GEN_8695; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8697 = 8'hf9 == io_state_in_9 ? 8'h99 : _GEN_8696; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8698 = 8'hfa == io_state_in_9 ? 8'h84 : _GEN_8697; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8699 = 8'hfb == io_state_in_9 ? 8'h8f : _GEN_8698; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8700 = 8'hfc == io_state_in_9 ? 8'hbe : _GEN_8699; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8701 = 8'hfd == io_state_in_9 ? 8'hb5 : _GEN_8700; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8702 = 8'hfe == io_state_in_9 ? 8'ha8 : _GEN_8701; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _GEN_8703 = 8'hff == io_state_in_9 ? 8'ha3 : _GEN_8702; // @[InvMixColumns.scala 136:{41,41}]
  wire [7:0] _tmp_state_8_T = _GEN_8447 ^ _GEN_8703; // @[InvMixColumns.scala 136:41]
  wire [7:0] _GEN_8705 = 8'h1 == io_state_in_10 ? 8'hd : 8'h0; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8706 = 8'h2 == io_state_in_10 ? 8'h1a : _GEN_8705; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8707 = 8'h3 == io_state_in_10 ? 8'h17 : _GEN_8706; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8708 = 8'h4 == io_state_in_10 ? 8'h34 : _GEN_8707; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8709 = 8'h5 == io_state_in_10 ? 8'h39 : _GEN_8708; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8710 = 8'h6 == io_state_in_10 ? 8'h2e : _GEN_8709; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8711 = 8'h7 == io_state_in_10 ? 8'h23 : _GEN_8710; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8712 = 8'h8 == io_state_in_10 ? 8'h68 : _GEN_8711; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8713 = 8'h9 == io_state_in_10 ? 8'h65 : _GEN_8712; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8714 = 8'ha == io_state_in_10 ? 8'h72 : _GEN_8713; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8715 = 8'hb == io_state_in_10 ? 8'h7f : _GEN_8714; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8716 = 8'hc == io_state_in_10 ? 8'h5c : _GEN_8715; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8717 = 8'hd == io_state_in_10 ? 8'h51 : _GEN_8716; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8718 = 8'he == io_state_in_10 ? 8'h46 : _GEN_8717; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8719 = 8'hf == io_state_in_10 ? 8'h4b : _GEN_8718; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8720 = 8'h10 == io_state_in_10 ? 8'hd0 : _GEN_8719; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8721 = 8'h11 == io_state_in_10 ? 8'hdd : _GEN_8720; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8722 = 8'h12 == io_state_in_10 ? 8'hca : _GEN_8721; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8723 = 8'h13 == io_state_in_10 ? 8'hc7 : _GEN_8722; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8724 = 8'h14 == io_state_in_10 ? 8'he4 : _GEN_8723; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8725 = 8'h15 == io_state_in_10 ? 8'he9 : _GEN_8724; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8726 = 8'h16 == io_state_in_10 ? 8'hfe : _GEN_8725; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8727 = 8'h17 == io_state_in_10 ? 8'hf3 : _GEN_8726; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8728 = 8'h18 == io_state_in_10 ? 8'hb8 : _GEN_8727; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8729 = 8'h19 == io_state_in_10 ? 8'hb5 : _GEN_8728; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8730 = 8'h1a == io_state_in_10 ? 8'ha2 : _GEN_8729; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8731 = 8'h1b == io_state_in_10 ? 8'haf : _GEN_8730; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8732 = 8'h1c == io_state_in_10 ? 8'h8c : _GEN_8731; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8733 = 8'h1d == io_state_in_10 ? 8'h81 : _GEN_8732; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8734 = 8'h1e == io_state_in_10 ? 8'h96 : _GEN_8733; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8735 = 8'h1f == io_state_in_10 ? 8'h9b : _GEN_8734; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8736 = 8'h20 == io_state_in_10 ? 8'hbb : _GEN_8735; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8737 = 8'h21 == io_state_in_10 ? 8'hb6 : _GEN_8736; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8738 = 8'h22 == io_state_in_10 ? 8'ha1 : _GEN_8737; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8739 = 8'h23 == io_state_in_10 ? 8'hac : _GEN_8738; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8740 = 8'h24 == io_state_in_10 ? 8'h8f : _GEN_8739; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8741 = 8'h25 == io_state_in_10 ? 8'h82 : _GEN_8740; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8742 = 8'h26 == io_state_in_10 ? 8'h95 : _GEN_8741; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8743 = 8'h27 == io_state_in_10 ? 8'h98 : _GEN_8742; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8744 = 8'h28 == io_state_in_10 ? 8'hd3 : _GEN_8743; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8745 = 8'h29 == io_state_in_10 ? 8'hde : _GEN_8744; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8746 = 8'h2a == io_state_in_10 ? 8'hc9 : _GEN_8745; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8747 = 8'h2b == io_state_in_10 ? 8'hc4 : _GEN_8746; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8748 = 8'h2c == io_state_in_10 ? 8'he7 : _GEN_8747; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8749 = 8'h2d == io_state_in_10 ? 8'hea : _GEN_8748; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8750 = 8'h2e == io_state_in_10 ? 8'hfd : _GEN_8749; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8751 = 8'h2f == io_state_in_10 ? 8'hf0 : _GEN_8750; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8752 = 8'h30 == io_state_in_10 ? 8'h6b : _GEN_8751; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8753 = 8'h31 == io_state_in_10 ? 8'h66 : _GEN_8752; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8754 = 8'h32 == io_state_in_10 ? 8'h71 : _GEN_8753; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8755 = 8'h33 == io_state_in_10 ? 8'h7c : _GEN_8754; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8756 = 8'h34 == io_state_in_10 ? 8'h5f : _GEN_8755; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8757 = 8'h35 == io_state_in_10 ? 8'h52 : _GEN_8756; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8758 = 8'h36 == io_state_in_10 ? 8'h45 : _GEN_8757; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8759 = 8'h37 == io_state_in_10 ? 8'h48 : _GEN_8758; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8760 = 8'h38 == io_state_in_10 ? 8'h3 : _GEN_8759; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8761 = 8'h39 == io_state_in_10 ? 8'he : _GEN_8760; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8762 = 8'h3a == io_state_in_10 ? 8'h19 : _GEN_8761; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8763 = 8'h3b == io_state_in_10 ? 8'h14 : _GEN_8762; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8764 = 8'h3c == io_state_in_10 ? 8'h37 : _GEN_8763; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8765 = 8'h3d == io_state_in_10 ? 8'h3a : _GEN_8764; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8766 = 8'h3e == io_state_in_10 ? 8'h2d : _GEN_8765; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8767 = 8'h3f == io_state_in_10 ? 8'h20 : _GEN_8766; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8768 = 8'h40 == io_state_in_10 ? 8'h6d : _GEN_8767; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8769 = 8'h41 == io_state_in_10 ? 8'h60 : _GEN_8768; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8770 = 8'h42 == io_state_in_10 ? 8'h77 : _GEN_8769; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8771 = 8'h43 == io_state_in_10 ? 8'h7a : _GEN_8770; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8772 = 8'h44 == io_state_in_10 ? 8'h59 : _GEN_8771; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8773 = 8'h45 == io_state_in_10 ? 8'h54 : _GEN_8772; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8774 = 8'h46 == io_state_in_10 ? 8'h43 : _GEN_8773; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8775 = 8'h47 == io_state_in_10 ? 8'h4e : _GEN_8774; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8776 = 8'h48 == io_state_in_10 ? 8'h5 : _GEN_8775; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8777 = 8'h49 == io_state_in_10 ? 8'h8 : _GEN_8776; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8778 = 8'h4a == io_state_in_10 ? 8'h1f : _GEN_8777; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8779 = 8'h4b == io_state_in_10 ? 8'h12 : _GEN_8778; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8780 = 8'h4c == io_state_in_10 ? 8'h31 : _GEN_8779; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8781 = 8'h4d == io_state_in_10 ? 8'h3c : _GEN_8780; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8782 = 8'h4e == io_state_in_10 ? 8'h2b : _GEN_8781; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8783 = 8'h4f == io_state_in_10 ? 8'h26 : _GEN_8782; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8784 = 8'h50 == io_state_in_10 ? 8'hbd : _GEN_8783; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8785 = 8'h51 == io_state_in_10 ? 8'hb0 : _GEN_8784; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8786 = 8'h52 == io_state_in_10 ? 8'ha7 : _GEN_8785; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8787 = 8'h53 == io_state_in_10 ? 8'haa : _GEN_8786; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8788 = 8'h54 == io_state_in_10 ? 8'h89 : _GEN_8787; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8789 = 8'h55 == io_state_in_10 ? 8'h84 : _GEN_8788; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8790 = 8'h56 == io_state_in_10 ? 8'h93 : _GEN_8789; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8791 = 8'h57 == io_state_in_10 ? 8'h9e : _GEN_8790; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8792 = 8'h58 == io_state_in_10 ? 8'hd5 : _GEN_8791; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8793 = 8'h59 == io_state_in_10 ? 8'hd8 : _GEN_8792; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8794 = 8'h5a == io_state_in_10 ? 8'hcf : _GEN_8793; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8795 = 8'h5b == io_state_in_10 ? 8'hc2 : _GEN_8794; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8796 = 8'h5c == io_state_in_10 ? 8'he1 : _GEN_8795; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8797 = 8'h5d == io_state_in_10 ? 8'hec : _GEN_8796; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8798 = 8'h5e == io_state_in_10 ? 8'hfb : _GEN_8797; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8799 = 8'h5f == io_state_in_10 ? 8'hf6 : _GEN_8798; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8800 = 8'h60 == io_state_in_10 ? 8'hd6 : _GEN_8799; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8801 = 8'h61 == io_state_in_10 ? 8'hdb : _GEN_8800; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8802 = 8'h62 == io_state_in_10 ? 8'hcc : _GEN_8801; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8803 = 8'h63 == io_state_in_10 ? 8'hc1 : _GEN_8802; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8804 = 8'h64 == io_state_in_10 ? 8'he2 : _GEN_8803; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8805 = 8'h65 == io_state_in_10 ? 8'hef : _GEN_8804; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8806 = 8'h66 == io_state_in_10 ? 8'hf8 : _GEN_8805; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8807 = 8'h67 == io_state_in_10 ? 8'hf5 : _GEN_8806; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8808 = 8'h68 == io_state_in_10 ? 8'hbe : _GEN_8807; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8809 = 8'h69 == io_state_in_10 ? 8'hb3 : _GEN_8808; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8810 = 8'h6a == io_state_in_10 ? 8'ha4 : _GEN_8809; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8811 = 8'h6b == io_state_in_10 ? 8'ha9 : _GEN_8810; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8812 = 8'h6c == io_state_in_10 ? 8'h8a : _GEN_8811; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8813 = 8'h6d == io_state_in_10 ? 8'h87 : _GEN_8812; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8814 = 8'h6e == io_state_in_10 ? 8'h90 : _GEN_8813; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8815 = 8'h6f == io_state_in_10 ? 8'h9d : _GEN_8814; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8816 = 8'h70 == io_state_in_10 ? 8'h6 : _GEN_8815; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8817 = 8'h71 == io_state_in_10 ? 8'hb : _GEN_8816; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8818 = 8'h72 == io_state_in_10 ? 8'h1c : _GEN_8817; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8819 = 8'h73 == io_state_in_10 ? 8'h11 : _GEN_8818; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8820 = 8'h74 == io_state_in_10 ? 8'h32 : _GEN_8819; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8821 = 8'h75 == io_state_in_10 ? 8'h3f : _GEN_8820; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8822 = 8'h76 == io_state_in_10 ? 8'h28 : _GEN_8821; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8823 = 8'h77 == io_state_in_10 ? 8'h25 : _GEN_8822; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8824 = 8'h78 == io_state_in_10 ? 8'h6e : _GEN_8823; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8825 = 8'h79 == io_state_in_10 ? 8'h63 : _GEN_8824; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8826 = 8'h7a == io_state_in_10 ? 8'h74 : _GEN_8825; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8827 = 8'h7b == io_state_in_10 ? 8'h79 : _GEN_8826; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8828 = 8'h7c == io_state_in_10 ? 8'h5a : _GEN_8827; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8829 = 8'h7d == io_state_in_10 ? 8'h57 : _GEN_8828; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8830 = 8'h7e == io_state_in_10 ? 8'h40 : _GEN_8829; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8831 = 8'h7f == io_state_in_10 ? 8'h4d : _GEN_8830; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8832 = 8'h80 == io_state_in_10 ? 8'hda : _GEN_8831; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8833 = 8'h81 == io_state_in_10 ? 8'hd7 : _GEN_8832; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8834 = 8'h82 == io_state_in_10 ? 8'hc0 : _GEN_8833; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8835 = 8'h83 == io_state_in_10 ? 8'hcd : _GEN_8834; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8836 = 8'h84 == io_state_in_10 ? 8'hee : _GEN_8835; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8837 = 8'h85 == io_state_in_10 ? 8'he3 : _GEN_8836; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8838 = 8'h86 == io_state_in_10 ? 8'hf4 : _GEN_8837; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8839 = 8'h87 == io_state_in_10 ? 8'hf9 : _GEN_8838; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8840 = 8'h88 == io_state_in_10 ? 8'hb2 : _GEN_8839; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8841 = 8'h89 == io_state_in_10 ? 8'hbf : _GEN_8840; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8842 = 8'h8a == io_state_in_10 ? 8'ha8 : _GEN_8841; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8843 = 8'h8b == io_state_in_10 ? 8'ha5 : _GEN_8842; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8844 = 8'h8c == io_state_in_10 ? 8'h86 : _GEN_8843; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8845 = 8'h8d == io_state_in_10 ? 8'h8b : _GEN_8844; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8846 = 8'h8e == io_state_in_10 ? 8'h9c : _GEN_8845; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8847 = 8'h8f == io_state_in_10 ? 8'h91 : _GEN_8846; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8848 = 8'h90 == io_state_in_10 ? 8'ha : _GEN_8847; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8849 = 8'h91 == io_state_in_10 ? 8'h7 : _GEN_8848; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8850 = 8'h92 == io_state_in_10 ? 8'h10 : _GEN_8849; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8851 = 8'h93 == io_state_in_10 ? 8'h1d : _GEN_8850; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8852 = 8'h94 == io_state_in_10 ? 8'h3e : _GEN_8851; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8853 = 8'h95 == io_state_in_10 ? 8'h33 : _GEN_8852; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8854 = 8'h96 == io_state_in_10 ? 8'h24 : _GEN_8853; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8855 = 8'h97 == io_state_in_10 ? 8'h29 : _GEN_8854; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8856 = 8'h98 == io_state_in_10 ? 8'h62 : _GEN_8855; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8857 = 8'h99 == io_state_in_10 ? 8'h6f : _GEN_8856; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8858 = 8'h9a == io_state_in_10 ? 8'h78 : _GEN_8857; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8859 = 8'h9b == io_state_in_10 ? 8'h75 : _GEN_8858; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8860 = 8'h9c == io_state_in_10 ? 8'h56 : _GEN_8859; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8861 = 8'h9d == io_state_in_10 ? 8'h5b : _GEN_8860; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8862 = 8'h9e == io_state_in_10 ? 8'h4c : _GEN_8861; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8863 = 8'h9f == io_state_in_10 ? 8'h41 : _GEN_8862; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8864 = 8'ha0 == io_state_in_10 ? 8'h61 : _GEN_8863; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8865 = 8'ha1 == io_state_in_10 ? 8'h6c : _GEN_8864; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8866 = 8'ha2 == io_state_in_10 ? 8'h7b : _GEN_8865; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8867 = 8'ha3 == io_state_in_10 ? 8'h76 : _GEN_8866; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8868 = 8'ha4 == io_state_in_10 ? 8'h55 : _GEN_8867; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8869 = 8'ha5 == io_state_in_10 ? 8'h58 : _GEN_8868; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8870 = 8'ha6 == io_state_in_10 ? 8'h4f : _GEN_8869; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8871 = 8'ha7 == io_state_in_10 ? 8'h42 : _GEN_8870; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8872 = 8'ha8 == io_state_in_10 ? 8'h9 : _GEN_8871; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8873 = 8'ha9 == io_state_in_10 ? 8'h4 : _GEN_8872; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8874 = 8'haa == io_state_in_10 ? 8'h13 : _GEN_8873; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8875 = 8'hab == io_state_in_10 ? 8'h1e : _GEN_8874; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8876 = 8'hac == io_state_in_10 ? 8'h3d : _GEN_8875; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8877 = 8'had == io_state_in_10 ? 8'h30 : _GEN_8876; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8878 = 8'hae == io_state_in_10 ? 8'h27 : _GEN_8877; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8879 = 8'haf == io_state_in_10 ? 8'h2a : _GEN_8878; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8880 = 8'hb0 == io_state_in_10 ? 8'hb1 : _GEN_8879; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8881 = 8'hb1 == io_state_in_10 ? 8'hbc : _GEN_8880; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8882 = 8'hb2 == io_state_in_10 ? 8'hab : _GEN_8881; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8883 = 8'hb3 == io_state_in_10 ? 8'ha6 : _GEN_8882; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8884 = 8'hb4 == io_state_in_10 ? 8'h85 : _GEN_8883; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8885 = 8'hb5 == io_state_in_10 ? 8'h88 : _GEN_8884; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8886 = 8'hb6 == io_state_in_10 ? 8'h9f : _GEN_8885; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8887 = 8'hb7 == io_state_in_10 ? 8'h92 : _GEN_8886; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8888 = 8'hb8 == io_state_in_10 ? 8'hd9 : _GEN_8887; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8889 = 8'hb9 == io_state_in_10 ? 8'hd4 : _GEN_8888; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8890 = 8'hba == io_state_in_10 ? 8'hc3 : _GEN_8889; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8891 = 8'hbb == io_state_in_10 ? 8'hce : _GEN_8890; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8892 = 8'hbc == io_state_in_10 ? 8'hed : _GEN_8891; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8893 = 8'hbd == io_state_in_10 ? 8'he0 : _GEN_8892; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8894 = 8'hbe == io_state_in_10 ? 8'hf7 : _GEN_8893; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8895 = 8'hbf == io_state_in_10 ? 8'hfa : _GEN_8894; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8896 = 8'hc0 == io_state_in_10 ? 8'hb7 : _GEN_8895; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8897 = 8'hc1 == io_state_in_10 ? 8'hba : _GEN_8896; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8898 = 8'hc2 == io_state_in_10 ? 8'had : _GEN_8897; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8899 = 8'hc3 == io_state_in_10 ? 8'ha0 : _GEN_8898; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8900 = 8'hc4 == io_state_in_10 ? 8'h83 : _GEN_8899; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8901 = 8'hc5 == io_state_in_10 ? 8'h8e : _GEN_8900; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8902 = 8'hc6 == io_state_in_10 ? 8'h99 : _GEN_8901; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8903 = 8'hc7 == io_state_in_10 ? 8'h94 : _GEN_8902; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8904 = 8'hc8 == io_state_in_10 ? 8'hdf : _GEN_8903; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8905 = 8'hc9 == io_state_in_10 ? 8'hd2 : _GEN_8904; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8906 = 8'hca == io_state_in_10 ? 8'hc5 : _GEN_8905; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8907 = 8'hcb == io_state_in_10 ? 8'hc8 : _GEN_8906; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8908 = 8'hcc == io_state_in_10 ? 8'heb : _GEN_8907; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8909 = 8'hcd == io_state_in_10 ? 8'he6 : _GEN_8908; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8910 = 8'hce == io_state_in_10 ? 8'hf1 : _GEN_8909; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8911 = 8'hcf == io_state_in_10 ? 8'hfc : _GEN_8910; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8912 = 8'hd0 == io_state_in_10 ? 8'h67 : _GEN_8911; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8913 = 8'hd1 == io_state_in_10 ? 8'h6a : _GEN_8912; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8914 = 8'hd2 == io_state_in_10 ? 8'h7d : _GEN_8913; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8915 = 8'hd3 == io_state_in_10 ? 8'h70 : _GEN_8914; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8916 = 8'hd4 == io_state_in_10 ? 8'h53 : _GEN_8915; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8917 = 8'hd5 == io_state_in_10 ? 8'h5e : _GEN_8916; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8918 = 8'hd6 == io_state_in_10 ? 8'h49 : _GEN_8917; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8919 = 8'hd7 == io_state_in_10 ? 8'h44 : _GEN_8918; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8920 = 8'hd8 == io_state_in_10 ? 8'hf : _GEN_8919; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8921 = 8'hd9 == io_state_in_10 ? 8'h2 : _GEN_8920; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8922 = 8'hda == io_state_in_10 ? 8'h15 : _GEN_8921; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8923 = 8'hdb == io_state_in_10 ? 8'h18 : _GEN_8922; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8924 = 8'hdc == io_state_in_10 ? 8'h3b : _GEN_8923; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8925 = 8'hdd == io_state_in_10 ? 8'h36 : _GEN_8924; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8926 = 8'hde == io_state_in_10 ? 8'h21 : _GEN_8925; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8927 = 8'hdf == io_state_in_10 ? 8'h2c : _GEN_8926; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8928 = 8'he0 == io_state_in_10 ? 8'hc : _GEN_8927; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8929 = 8'he1 == io_state_in_10 ? 8'h1 : _GEN_8928; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8930 = 8'he2 == io_state_in_10 ? 8'h16 : _GEN_8929; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8931 = 8'he3 == io_state_in_10 ? 8'h1b : _GEN_8930; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8932 = 8'he4 == io_state_in_10 ? 8'h38 : _GEN_8931; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8933 = 8'he5 == io_state_in_10 ? 8'h35 : _GEN_8932; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8934 = 8'he6 == io_state_in_10 ? 8'h22 : _GEN_8933; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8935 = 8'he7 == io_state_in_10 ? 8'h2f : _GEN_8934; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8936 = 8'he8 == io_state_in_10 ? 8'h64 : _GEN_8935; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8937 = 8'he9 == io_state_in_10 ? 8'h69 : _GEN_8936; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8938 = 8'hea == io_state_in_10 ? 8'h7e : _GEN_8937; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8939 = 8'heb == io_state_in_10 ? 8'h73 : _GEN_8938; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8940 = 8'hec == io_state_in_10 ? 8'h50 : _GEN_8939; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8941 = 8'hed == io_state_in_10 ? 8'h5d : _GEN_8940; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8942 = 8'hee == io_state_in_10 ? 8'h4a : _GEN_8941; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8943 = 8'hef == io_state_in_10 ? 8'h47 : _GEN_8942; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8944 = 8'hf0 == io_state_in_10 ? 8'hdc : _GEN_8943; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8945 = 8'hf1 == io_state_in_10 ? 8'hd1 : _GEN_8944; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8946 = 8'hf2 == io_state_in_10 ? 8'hc6 : _GEN_8945; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8947 = 8'hf3 == io_state_in_10 ? 8'hcb : _GEN_8946; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8948 = 8'hf4 == io_state_in_10 ? 8'he8 : _GEN_8947; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8949 = 8'hf5 == io_state_in_10 ? 8'he5 : _GEN_8948; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8950 = 8'hf6 == io_state_in_10 ? 8'hf2 : _GEN_8949; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8951 = 8'hf7 == io_state_in_10 ? 8'hff : _GEN_8950; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8952 = 8'hf8 == io_state_in_10 ? 8'hb4 : _GEN_8951; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8953 = 8'hf9 == io_state_in_10 ? 8'hb9 : _GEN_8952; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8954 = 8'hfa == io_state_in_10 ? 8'hae : _GEN_8953; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8955 = 8'hfb == io_state_in_10 ? 8'ha3 : _GEN_8954; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8956 = 8'hfc == io_state_in_10 ? 8'h80 : _GEN_8955; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8957 = 8'hfd == io_state_in_10 ? 8'h8d : _GEN_8956; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8958 = 8'hfe == io_state_in_10 ? 8'h9a : _GEN_8957; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _GEN_8959 = 8'hff == io_state_in_10 ? 8'h97 : _GEN_8958; // @[InvMixColumns.scala 136:{65,65}]
  wire [7:0] _tmp_state_8_T_1 = _tmp_state_8_T ^ _GEN_8959; // @[InvMixColumns.scala 136:65]
  wire [7:0] _GEN_8961 = 8'h1 == io_state_in_11 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8962 = 8'h2 == io_state_in_11 ? 8'h12 : _GEN_8961; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8963 = 8'h3 == io_state_in_11 ? 8'h1b : _GEN_8962; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8964 = 8'h4 == io_state_in_11 ? 8'h24 : _GEN_8963; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8965 = 8'h5 == io_state_in_11 ? 8'h2d : _GEN_8964; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8966 = 8'h6 == io_state_in_11 ? 8'h36 : _GEN_8965; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8967 = 8'h7 == io_state_in_11 ? 8'h3f : _GEN_8966; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8968 = 8'h8 == io_state_in_11 ? 8'h48 : _GEN_8967; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8969 = 8'h9 == io_state_in_11 ? 8'h41 : _GEN_8968; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8970 = 8'ha == io_state_in_11 ? 8'h5a : _GEN_8969; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8971 = 8'hb == io_state_in_11 ? 8'h53 : _GEN_8970; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8972 = 8'hc == io_state_in_11 ? 8'h6c : _GEN_8971; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8973 = 8'hd == io_state_in_11 ? 8'h65 : _GEN_8972; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8974 = 8'he == io_state_in_11 ? 8'h7e : _GEN_8973; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8975 = 8'hf == io_state_in_11 ? 8'h77 : _GEN_8974; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8976 = 8'h10 == io_state_in_11 ? 8'h90 : _GEN_8975; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8977 = 8'h11 == io_state_in_11 ? 8'h99 : _GEN_8976; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8978 = 8'h12 == io_state_in_11 ? 8'h82 : _GEN_8977; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8979 = 8'h13 == io_state_in_11 ? 8'h8b : _GEN_8978; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8980 = 8'h14 == io_state_in_11 ? 8'hb4 : _GEN_8979; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8981 = 8'h15 == io_state_in_11 ? 8'hbd : _GEN_8980; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8982 = 8'h16 == io_state_in_11 ? 8'ha6 : _GEN_8981; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8983 = 8'h17 == io_state_in_11 ? 8'haf : _GEN_8982; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8984 = 8'h18 == io_state_in_11 ? 8'hd8 : _GEN_8983; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8985 = 8'h19 == io_state_in_11 ? 8'hd1 : _GEN_8984; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8986 = 8'h1a == io_state_in_11 ? 8'hca : _GEN_8985; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8987 = 8'h1b == io_state_in_11 ? 8'hc3 : _GEN_8986; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8988 = 8'h1c == io_state_in_11 ? 8'hfc : _GEN_8987; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8989 = 8'h1d == io_state_in_11 ? 8'hf5 : _GEN_8988; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8990 = 8'h1e == io_state_in_11 ? 8'hee : _GEN_8989; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8991 = 8'h1f == io_state_in_11 ? 8'he7 : _GEN_8990; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8992 = 8'h20 == io_state_in_11 ? 8'h3b : _GEN_8991; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8993 = 8'h21 == io_state_in_11 ? 8'h32 : _GEN_8992; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8994 = 8'h22 == io_state_in_11 ? 8'h29 : _GEN_8993; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8995 = 8'h23 == io_state_in_11 ? 8'h20 : _GEN_8994; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8996 = 8'h24 == io_state_in_11 ? 8'h1f : _GEN_8995; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8997 = 8'h25 == io_state_in_11 ? 8'h16 : _GEN_8996; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8998 = 8'h26 == io_state_in_11 ? 8'hd : _GEN_8997; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_8999 = 8'h27 == io_state_in_11 ? 8'h4 : _GEN_8998; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9000 = 8'h28 == io_state_in_11 ? 8'h73 : _GEN_8999; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9001 = 8'h29 == io_state_in_11 ? 8'h7a : _GEN_9000; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9002 = 8'h2a == io_state_in_11 ? 8'h61 : _GEN_9001; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9003 = 8'h2b == io_state_in_11 ? 8'h68 : _GEN_9002; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9004 = 8'h2c == io_state_in_11 ? 8'h57 : _GEN_9003; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9005 = 8'h2d == io_state_in_11 ? 8'h5e : _GEN_9004; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9006 = 8'h2e == io_state_in_11 ? 8'h45 : _GEN_9005; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9007 = 8'h2f == io_state_in_11 ? 8'h4c : _GEN_9006; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9008 = 8'h30 == io_state_in_11 ? 8'hab : _GEN_9007; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9009 = 8'h31 == io_state_in_11 ? 8'ha2 : _GEN_9008; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9010 = 8'h32 == io_state_in_11 ? 8'hb9 : _GEN_9009; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9011 = 8'h33 == io_state_in_11 ? 8'hb0 : _GEN_9010; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9012 = 8'h34 == io_state_in_11 ? 8'h8f : _GEN_9011; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9013 = 8'h35 == io_state_in_11 ? 8'h86 : _GEN_9012; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9014 = 8'h36 == io_state_in_11 ? 8'h9d : _GEN_9013; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9015 = 8'h37 == io_state_in_11 ? 8'h94 : _GEN_9014; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9016 = 8'h38 == io_state_in_11 ? 8'he3 : _GEN_9015; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9017 = 8'h39 == io_state_in_11 ? 8'hea : _GEN_9016; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9018 = 8'h3a == io_state_in_11 ? 8'hf1 : _GEN_9017; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9019 = 8'h3b == io_state_in_11 ? 8'hf8 : _GEN_9018; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9020 = 8'h3c == io_state_in_11 ? 8'hc7 : _GEN_9019; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9021 = 8'h3d == io_state_in_11 ? 8'hce : _GEN_9020; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9022 = 8'h3e == io_state_in_11 ? 8'hd5 : _GEN_9021; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9023 = 8'h3f == io_state_in_11 ? 8'hdc : _GEN_9022; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9024 = 8'h40 == io_state_in_11 ? 8'h76 : _GEN_9023; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9025 = 8'h41 == io_state_in_11 ? 8'h7f : _GEN_9024; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9026 = 8'h42 == io_state_in_11 ? 8'h64 : _GEN_9025; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9027 = 8'h43 == io_state_in_11 ? 8'h6d : _GEN_9026; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9028 = 8'h44 == io_state_in_11 ? 8'h52 : _GEN_9027; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9029 = 8'h45 == io_state_in_11 ? 8'h5b : _GEN_9028; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9030 = 8'h46 == io_state_in_11 ? 8'h40 : _GEN_9029; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9031 = 8'h47 == io_state_in_11 ? 8'h49 : _GEN_9030; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9032 = 8'h48 == io_state_in_11 ? 8'h3e : _GEN_9031; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9033 = 8'h49 == io_state_in_11 ? 8'h37 : _GEN_9032; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9034 = 8'h4a == io_state_in_11 ? 8'h2c : _GEN_9033; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9035 = 8'h4b == io_state_in_11 ? 8'h25 : _GEN_9034; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9036 = 8'h4c == io_state_in_11 ? 8'h1a : _GEN_9035; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9037 = 8'h4d == io_state_in_11 ? 8'h13 : _GEN_9036; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9038 = 8'h4e == io_state_in_11 ? 8'h8 : _GEN_9037; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9039 = 8'h4f == io_state_in_11 ? 8'h1 : _GEN_9038; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9040 = 8'h50 == io_state_in_11 ? 8'he6 : _GEN_9039; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9041 = 8'h51 == io_state_in_11 ? 8'hef : _GEN_9040; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9042 = 8'h52 == io_state_in_11 ? 8'hf4 : _GEN_9041; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9043 = 8'h53 == io_state_in_11 ? 8'hfd : _GEN_9042; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9044 = 8'h54 == io_state_in_11 ? 8'hc2 : _GEN_9043; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9045 = 8'h55 == io_state_in_11 ? 8'hcb : _GEN_9044; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9046 = 8'h56 == io_state_in_11 ? 8'hd0 : _GEN_9045; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9047 = 8'h57 == io_state_in_11 ? 8'hd9 : _GEN_9046; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9048 = 8'h58 == io_state_in_11 ? 8'hae : _GEN_9047; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9049 = 8'h59 == io_state_in_11 ? 8'ha7 : _GEN_9048; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9050 = 8'h5a == io_state_in_11 ? 8'hbc : _GEN_9049; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9051 = 8'h5b == io_state_in_11 ? 8'hb5 : _GEN_9050; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9052 = 8'h5c == io_state_in_11 ? 8'h8a : _GEN_9051; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9053 = 8'h5d == io_state_in_11 ? 8'h83 : _GEN_9052; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9054 = 8'h5e == io_state_in_11 ? 8'h98 : _GEN_9053; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9055 = 8'h5f == io_state_in_11 ? 8'h91 : _GEN_9054; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9056 = 8'h60 == io_state_in_11 ? 8'h4d : _GEN_9055; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9057 = 8'h61 == io_state_in_11 ? 8'h44 : _GEN_9056; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9058 = 8'h62 == io_state_in_11 ? 8'h5f : _GEN_9057; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9059 = 8'h63 == io_state_in_11 ? 8'h56 : _GEN_9058; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9060 = 8'h64 == io_state_in_11 ? 8'h69 : _GEN_9059; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9061 = 8'h65 == io_state_in_11 ? 8'h60 : _GEN_9060; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9062 = 8'h66 == io_state_in_11 ? 8'h7b : _GEN_9061; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9063 = 8'h67 == io_state_in_11 ? 8'h72 : _GEN_9062; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9064 = 8'h68 == io_state_in_11 ? 8'h5 : _GEN_9063; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9065 = 8'h69 == io_state_in_11 ? 8'hc : _GEN_9064; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9066 = 8'h6a == io_state_in_11 ? 8'h17 : _GEN_9065; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9067 = 8'h6b == io_state_in_11 ? 8'h1e : _GEN_9066; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9068 = 8'h6c == io_state_in_11 ? 8'h21 : _GEN_9067; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9069 = 8'h6d == io_state_in_11 ? 8'h28 : _GEN_9068; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9070 = 8'h6e == io_state_in_11 ? 8'h33 : _GEN_9069; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9071 = 8'h6f == io_state_in_11 ? 8'h3a : _GEN_9070; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9072 = 8'h70 == io_state_in_11 ? 8'hdd : _GEN_9071; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9073 = 8'h71 == io_state_in_11 ? 8'hd4 : _GEN_9072; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9074 = 8'h72 == io_state_in_11 ? 8'hcf : _GEN_9073; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9075 = 8'h73 == io_state_in_11 ? 8'hc6 : _GEN_9074; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9076 = 8'h74 == io_state_in_11 ? 8'hf9 : _GEN_9075; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9077 = 8'h75 == io_state_in_11 ? 8'hf0 : _GEN_9076; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9078 = 8'h76 == io_state_in_11 ? 8'heb : _GEN_9077; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9079 = 8'h77 == io_state_in_11 ? 8'he2 : _GEN_9078; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9080 = 8'h78 == io_state_in_11 ? 8'h95 : _GEN_9079; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9081 = 8'h79 == io_state_in_11 ? 8'h9c : _GEN_9080; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9082 = 8'h7a == io_state_in_11 ? 8'h87 : _GEN_9081; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9083 = 8'h7b == io_state_in_11 ? 8'h8e : _GEN_9082; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9084 = 8'h7c == io_state_in_11 ? 8'hb1 : _GEN_9083; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9085 = 8'h7d == io_state_in_11 ? 8'hb8 : _GEN_9084; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9086 = 8'h7e == io_state_in_11 ? 8'ha3 : _GEN_9085; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9087 = 8'h7f == io_state_in_11 ? 8'haa : _GEN_9086; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9088 = 8'h80 == io_state_in_11 ? 8'hec : _GEN_9087; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9089 = 8'h81 == io_state_in_11 ? 8'he5 : _GEN_9088; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9090 = 8'h82 == io_state_in_11 ? 8'hfe : _GEN_9089; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9091 = 8'h83 == io_state_in_11 ? 8'hf7 : _GEN_9090; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9092 = 8'h84 == io_state_in_11 ? 8'hc8 : _GEN_9091; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9093 = 8'h85 == io_state_in_11 ? 8'hc1 : _GEN_9092; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9094 = 8'h86 == io_state_in_11 ? 8'hda : _GEN_9093; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9095 = 8'h87 == io_state_in_11 ? 8'hd3 : _GEN_9094; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9096 = 8'h88 == io_state_in_11 ? 8'ha4 : _GEN_9095; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9097 = 8'h89 == io_state_in_11 ? 8'had : _GEN_9096; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9098 = 8'h8a == io_state_in_11 ? 8'hb6 : _GEN_9097; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9099 = 8'h8b == io_state_in_11 ? 8'hbf : _GEN_9098; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9100 = 8'h8c == io_state_in_11 ? 8'h80 : _GEN_9099; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9101 = 8'h8d == io_state_in_11 ? 8'h89 : _GEN_9100; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9102 = 8'h8e == io_state_in_11 ? 8'h92 : _GEN_9101; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9103 = 8'h8f == io_state_in_11 ? 8'h9b : _GEN_9102; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9104 = 8'h90 == io_state_in_11 ? 8'h7c : _GEN_9103; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9105 = 8'h91 == io_state_in_11 ? 8'h75 : _GEN_9104; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9106 = 8'h92 == io_state_in_11 ? 8'h6e : _GEN_9105; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9107 = 8'h93 == io_state_in_11 ? 8'h67 : _GEN_9106; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9108 = 8'h94 == io_state_in_11 ? 8'h58 : _GEN_9107; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9109 = 8'h95 == io_state_in_11 ? 8'h51 : _GEN_9108; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9110 = 8'h96 == io_state_in_11 ? 8'h4a : _GEN_9109; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9111 = 8'h97 == io_state_in_11 ? 8'h43 : _GEN_9110; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9112 = 8'h98 == io_state_in_11 ? 8'h34 : _GEN_9111; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9113 = 8'h99 == io_state_in_11 ? 8'h3d : _GEN_9112; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9114 = 8'h9a == io_state_in_11 ? 8'h26 : _GEN_9113; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9115 = 8'h9b == io_state_in_11 ? 8'h2f : _GEN_9114; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9116 = 8'h9c == io_state_in_11 ? 8'h10 : _GEN_9115; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9117 = 8'h9d == io_state_in_11 ? 8'h19 : _GEN_9116; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9118 = 8'h9e == io_state_in_11 ? 8'h2 : _GEN_9117; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9119 = 8'h9f == io_state_in_11 ? 8'hb : _GEN_9118; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9120 = 8'ha0 == io_state_in_11 ? 8'hd7 : _GEN_9119; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9121 = 8'ha1 == io_state_in_11 ? 8'hde : _GEN_9120; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9122 = 8'ha2 == io_state_in_11 ? 8'hc5 : _GEN_9121; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9123 = 8'ha3 == io_state_in_11 ? 8'hcc : _GEN_9122; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9124 = 8'ha4 == io_state_in_11 ? 8'hf3 : _GEN_9123; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9125 = 8'ha5 == io_state_in_11 ? 8'hfa : _GEN_9124; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9126 = 8'ha6 == io_state_in_11 ? 8'he1 : _GEN_9125; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9127 = 8'ha7 == io_state_in_11 ? 8'he8 : _GEN_9126; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9128 = 8'ha8 == io_state_in_11 ? 8'h9f : _GEN_9127; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9129 = 8'ha9 == io_state_in_11 ? 8'h96 : _GEN_9128; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9130 = 8'haa == io_state_in_11 ? 8'h8d : _GEN_9129; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9131 = 8'hab == io_state_in_11 ? 8'h84 : _GEN_9130; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9132 = 8'hac == io_state_in_11 ? 8'hbb : _GEN_9131; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9133 = 8'had == io_state_in_11 ? 8'hb2 : _GEN_9132; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9134 = 8'hae == io_state_in_11 ? 8'ha9 : _GEN_9133; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9135 = 8'haf == io_state_in_11 ? 8'ha0 : _GEN_9134; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9136 = 8'hb0 == io_state_in_11 ? 8'h47 : _GEN_9135; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9137 = 8'hb1 == io_state_in_11 ? 8'h4e : _GEN_9136; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9138 = 8'hb2 == io_state_in_11 ? 8'h55 : _GEN_9137; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9139 = 8'hb3 == io_state_in_11 ? 8'h5c : _GEN_9138; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9140 = 8'hb4 == io_state_in_11 ? 8'h63 : _GEN_9139; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9141 = 8'hb5 == io_state_in_11 ? 8'h6a : _GEN_9140; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9142 = 8'hb6 == io_state_in_11 ? 8'h71 : _GEN_9141; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9143 = 8'hb7 == io_state_in_11 ? 8'h78 : _GEN_9142; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9144 = 8'hb8 == io_state_in_11 ? 8'hf : _GEN_9143; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9145 = 8'hb9 == io_state_in_11 ? 8'h6 : _GEN_9144; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9146 = 8'hba == io_state_in_11 ? 8'h1d : _GEN_9145; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9147 = 8'hbb == io_state_in_11 ? 8'h14 : _GEN_9146; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9148 = 8'hbc == io_state_in_11 ? 8'h2b : _GEN_9147; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9149 = 8'hbd == io_state_in_11 ? 8'h22 : _GEN_9148; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9150 = 8'hbe == io_state_in_11 ? 8'h39 : _GEN_9149; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9151 = 8'hbf == io_state_in_11 ? 8'h30 : _GEN_9150; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9152 = 8'hc0 == io_state_in_11 ? 8'h9a : _GEN_9151; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9153 = 8'hc1 == io_state_in_11 ? 8'h93 : _GEN_9152; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9154 = 8'hc2 == io_state_in_11 ? 8'h88 : _GEN_9153; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9155 = 8'hc3 == io_state_in_11 ? 8'h81 : _GEN_9154; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9156 = 8'hc4 == io_state_in_11 ? 8'hbe : _GEN_9155; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9157 = 8'hc5 == io_state_in_11 ? 8'hb7 : _GEN_9156; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9158 = 8'hc6 == io_state_in_11 ? 8'hac : _GEN_9157; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9159 = 8'hc7 == io_state_in_11 ? 8'ha5 : _GEN_9158; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9160 = 8'hc8 == io_state_in_11 ? 8'hd2 : _GEN_9159; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9161 = 8'hc9 == io_state_in_11 ? 8'hdb : _GEN_9160; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9162 = 8'hca == io_state_in_11 ? 8'hc0 : _GEN_9161; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9163 = 8'hcb == io_state_in_11 ? 8'hc9 : _GEN_9162; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9164 = 8'hcc == io_state_in_11 ? 8'hf6 : _GEN_9163; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9165 = 8'hcd == io_state_in_11 ? 8'hff : _GEN_9164; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9166 = 8'hce == io_state_in_11 ? 8'he4 : _GEN_9165; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9167 = 8'hcf == io_state_in_11 ? 8'hed : _GEN_9166; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9168 = 8'hd0 == io_state_in_11 ? 8'ha : _GEN_9167; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9169 = 8'hd1 == io_state_in_11 ? 8'h3 : _GEN_9168; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9170 = 8'hd2 == io_state_in_11 ? 8'h18 : _GEN_9169; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9171 = 8'hd3 == io_state_in_11 ? 8'h11 : _GEN_9170; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9172 = 8'hd4 == io_state_in_11 ? 8'h2e : _GEN_9171; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9173 = 8'hd5 == io_state_in_11 ? 8'h27 : _GEN_9172; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9174 = 8'hd6 == io_state_in_11 ? 8'h3c : _GEN_9173; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9175 = 8'hd7 == io_state_in_11 ? 8'h35 : _GEN_9174; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9176 = 8'hd8 == io_state_in_11 ? 8'h42 : _GEN_9175; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9177 = 8'hd9 == io_state_in_11 ? 8'h4b : _GEN_9176; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9178 = 8'hda == io_state_in_11 ? 8'h50 : _GEN_9177; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9179 = 8'hdb == io_state_in_11 ? 8'h59 : _GEN_9178; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9180 = 8'hdc == io_state_in_11 ? 8'h66 : _GEN_9179; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9181 = 8'hdd == io_state_in_11 ? 8'h6f : _GEN_9180; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9182 = 8'hde == io_state_in_11 ? 8'h74 : _GEN_9181; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9183 = 8'hdf == io_state_in_11 ? 8'h7d : _GEN_9182; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9184 = 8'he0 == io_state_in_11 ? 8'ha1 : _GEN_9183; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9185 = 8'he1 == io_state_in_11 ? 8'ha8 : _GEN_9184; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9186 = 8'he2 == io_state_in_11 ? 8'hb3 : _GEN_9185; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9187 = 8'he3 == io_state_in_11 ? 8'hba : _GEN_9186; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9188 = 8'he4 == io_state_in_11 ? 8'h85 : _GEN_9187; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9189 = 8'he5 == io_state_in_11 ? 8'h8c : _GEN_9188; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9190 = 8'he6 == io_state_in_11 ? 8'h97 : _GEN_9189; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9191 = 8'he7 == io_state_in_11 ? 8'h9e : _GEN_9190; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9192 = 8'he8 == io_state_in_11 ? 8'he9 : _GEN_9191; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9193 = 8'he9 == io_state_in_11 ? 8'he0 : _GEN_9192; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9194 = 8'hea == io_state_in_11 ? 8'hfb : _GEN_9193; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9195 = 8'heb == io_state_in_11 ? 8'hf2 : _GEN_9194; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9196 = 8'hec == io_state_in_11 ? 8'hcd : _GEN_9195; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9197 = 8'hed == io_state_in_11 ? 8'hc4 : _GEN_9196; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9198 = 8'hee == io_state_in_11 ? 8'hdf : _GEN_9197; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9199 = 8'hef == io_state_in_11 ? 8'hd6 : _GEN_9198; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9200 = 8'hf0 == io_state_in_11 ? 8'h31 : _GEN_9199; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9201 = 8'hf1 == io_state_in_11 ? 8'h38 : _GEN_9200; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9202 = 8'hf2 == io_state_in_11 ? 8'h23 : _GEN_9201; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9203 = 8'hf3 == io_state_in_11 ? 8'h2a : _GEN_9202; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9204 = 8'hf4 == io_state_in_11 ? 8'h15 : _GEN_9203; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9205 = 8'hf5 == io_state_in_11 ? 8'h1c : _GEN_9204; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9206 = 8'hf6 == io_state_in_11 ? 8'h7 : _GEN_9205; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9207 = 8'hf7 == io_state_in_11 ? 8'he : _GEN_9206; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9208 = 8'hf8 == io_state_in_11 ? 8'h79 : _GEN_9207; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9209 = 8'hf9 == io_state_in_11 ? 8'h70 : _GEN_9208; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9210 = 8'hfa == io_state_in_11 ? 8'h6b : _GEN_9209; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9211 = 8'hfb == io_state_in_11 ? 8'h62 : _GEN_9210; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9212 = 8'hfc == io_state_in_11 ? 8'h5d : _GEN_9211; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9213 = 8'hfd == io_state_in_11 ? 8'h54 : _GEN_9212; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9214 = 8'hfe == io_state_in_11 ? 8'h4f : _GEN_9213; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9215 = 8'hff == io_state_in_11 ? 8'h46 : _GEN_9214; // @[InvMixColumns.scala 136:{90,90}]
  wire [7:0] _GEN_9217 = 8'h1 == io_state_in_8 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9218 = 8'h2 == io_state_in_8 ? 8'h12 : _GEN_9217; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9219 = 8'h3 == io_state_in_8 ? 8'h1b : _GEN_9218; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9220 = 8'h4 == io_state_in_8 ? 8'h24 : _GEN_9219; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9221 = 8'h5 == io_state_in_8 ? 8'h2d : _GEN_9220; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9222 = 8'h6 == io_state_in_8 ? 8'h36 : _GEN_9221; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9223 = 8'h7 == io_state_in_8 ? 8'h3f : _GEN_9222; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9224 = 8'h8 == io_state_in_8 ? 8'h48 : _GEN_9223; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9225 = 8'h9 == io_state_in_8 ? 8'h41 : _GEN_9224; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9226 = 8'ha == io_state_in_8 ? 8'h5a : _GEN_9225; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9227 = 8'hb == io_state_in_8 ? 8'h53 : _GEN_9226; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9228 = 8'hc == io_state_in_8 ? 8'h6c : _GEN_9227; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9229 = 8'hd == io_state_in_8 ? 8'h65 : _GEN_9228; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9230 = 8'he == io_state_in_8 ? 8'h7e : _GEN_9229; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9231 = 8'hf == io_state_in_8 ? 8'h77 : _GEN_9230; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9232 = 8'h10 == io_state_in_8 ? 8'h90 : _GEN_9231; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9233 = 8'h11 == io_state_in_8 ? 8'h99 : _GEN_9232; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9234 = 8'h12 == io_state_in_8 ? 8'h82 : _GEN_9233; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9235 = 8'h13 == io_state_in_8 ? 8'h8b : _GEN_9234; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9236 = 8'h14 == io_state_in_8 ? 8'hb4 : _GEN_9235; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9237 = 8'h15 == io_state_in_8 ? 8'hbd : _GEN_9236; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9238 = 8'h16 == io_state_in_8 ? 8'ha6 : _GEN_9237; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9239 = 8'h17 == io_state_in_8 ? 8'haf : _GEN_9238; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9240 = 8'h18 == io_state_in_8 ? 8'hd8 : _GEN_9239; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9241 = 8'h19 == io_state_in_8 ? 8'hd1 : _GEN_9240; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9242 = 8'h1a == io_state_in_8 ? 8'hca : _GEN_9241; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9243 = 8'h1b == io_state_in_8 ? 8'hc3 : _GEN_9242; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9244 = 8'h1c == io_state_in_8 ? 8'hfc : _GEN_9243; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9245 = 8'h1d == io_state_in_8 ? 8'hf5 : _GEN_9244; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9246 = 8'h1e == io_state_in_8 ? 8'hee : _GEN_9245; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9247 = 8'h1f == io_state_in_8 ? 8'he7 : _GEN_9246; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9248 = 8'h20 == io_state_in_8 ? 8'h3b : _GEN_9247; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9249 = 8'h21 == io_state_in_8 ? 8'h32 : _GEN_9248; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9250 = 8'h22 == io_state_in_8 ? 8'h29 : _GEN_9249; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9251 = 8'h23 == io_state_in_8 ? 8'h20 : _GEN_9250; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9252 = 8'h24 == io_state_in_8 ? 8'h1f : _GEN_9251; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9253 = 8'h25 == io_state_in_8 ? 8'h16 : _GEN_9252; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9254 = 8'h26 == io_state_in_8 ? 8'hd : _GEN_9253; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9255 = 8'h27 == io_state_in_8 ? 8'h4 : _GEN_9254; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9256 = 8'h28 == io_state_in_8 ? 8'h73 : _GEN_9255; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9257 = 8'h29 == io_state_in_8 ? 8'h7a : _GEN_9256; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9258 = 8'h2a == io_state_in_8 ? 8'h61 : _GEN_9257; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9259 = 8'h2b == io_state_in_8 ? 8'h68 : _GEN_9258; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9260 = 8'h2c == io_state_in_8 ? 8'h57 : _GEN_9259; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9261 = 8'h2d == io_state_in_8 ? 8'h5e : _GEN_9260; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9262 = 8'h2e == io_state_in_8 ? 8'h45 : _GEN_9261; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9263 = 8'h2f == io_state_in_8 ? 8'h4c : _GEN_9262; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9264 = 8'h30 == io_state_in_8 ? 8'hab : _GEN_9263; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9265 = 8'h31 == io_state_in_8 ? 8'ha2 : _GEN_9264; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9266 = 8'h32 == io_state_in_8 ? 8'hb9 : _GEN_9265; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9267 = 8'h33 == io_state_in_8 ? 8'hb0 : _GEN_9266; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9268 = 8'h34 == io_state_in_8 ? 8'h8f : _GEN_9267; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9269 = 8'h35 == io_state_in_8 ? 8'h86 : _GEN_9268; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9270 = 8'h36 == io_state_in_8 ? 8'h9d : _GEN_9269; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9271 = 8'h37 == io_state_in_8 ? 8'h94 : _GEN_9270; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9272 = 8'h38 == io_state_in_8 ? 8'he3 : _GEN_9271; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9273 = 8'h39 == io_state_in_8 ? 8'hea : _GEN_9272; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9274 = 8'h3a == io_state_in_8 ? 8'hf1 : _GEN_9273; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9275 = 8'h3b == io_state_in_8 ? 8'hf8 : _GEN_9274; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9276 = 8'h3c == io_state_in_8 ? 8'hc7 : _GEN_9275; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9277 = 8'h3d == io_state_in_8 ? 8'hce : _GEN_9276; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9278 = 8'h3e == io_state_in_8 ? 8'hd5 : _GEN_9277; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9279 = 8'h3f == io_state_in_8 ? 8'hdc : _GEN_9278; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9280 = 8'h40 == io_state_in_8 ? 8'h76 : _GEN_9279; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9281 = 8'h41 == io_state_in_8 ? 8'h7f : _GEN_9280; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9282 = 8'h42 == io_state_in_8 ? 8'h64 : _GEN_9281; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9283 = 8'h43 == io_state_in_8 ? 8'h6d : _GEN_9282; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9284 = 8'h44 == io_state_in_8 ? 8'h52 : _GEN_9283; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9285 = 8'h45 == io_state_in_8 ? 8'h5b : _GEN_9284; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9286 = 8'h46 == io_state_in_8 ? 8'h40 : _GEN_9285; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9287 = 8'h47 == io_state_in_8 ? 8'h49 : _GEN_9286; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9288 = 8'h48 == io_state_in_8 ? 8'h3e : _GEN_9287; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9289 = 8'h49 == io_state_in_8 ? 8'h37 : _GEN_9288; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9290 = 8'h4a == io_state_in_8 ? 8'h2c : _GEN_9289; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9291 = 8'h4b == io_state_in_8 ? 8'h25 : _GEN_9290; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9292 = 8'h4c == io_state_in_8 ? 8'h1a : _GEN_9291; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9293 = 8'h4d == io_state_in_8 ? 8'h13 : _GEN_9292; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9294 = 8'h4e == io_state_in_8 ? 8'h8 : _GEN_9293; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9295 = 8'h4f == io_state_in_8 ? 8'h1 : _GEN_9294; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9296 = 8'h50 == io_state_in_8 ? 8'he6 : _GEN_9295; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9297 = 8'h51 == io_state_in_8 ? 8'hef : _GEN_9296; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9298 = 8'h52 == io_state_in_8 ? 8'hf4 : _GEN_9297; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9299 = 8'h53 == io_state_in_8 ? 8'hfd : _GEN_9298; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9300 = 8'h54 == io_state_in_8 ? 8'hc2 : _GEN_9299; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9301 = 8'h55 == io_state_in_8 ? 8'hcb : _GEN_9300; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9302 = 8'h56 == io_state_in_8 ? 8'hd0 : _GEN_9301; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9303 = 8'h57 == io_state_in_8 ? 8'hd9 : _GEN_9302; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9304 = 8'h58 == io_state_in_8 ? 8'hae : _GEN_9303; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9305 = 8'h59 == io_state_in_8 ? 8'ha7 : _GEN_9304; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9306 = 8'h5a == io_state_in_8 ? 8'hbc : _GEN_9305; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9307 = 8'h5b == io_state_in_8 ? 8'hb5 : _GEN_9306; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9308 = 8'h5c == io_state_in_8 ? 8'h8a : _GEN_9307; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9309 = 8'h5d == io_state_in_8 ? 8'h83 : _GEN_9308; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9310 = 8'h5e == io_state_in_8 ? 8'h98 : _GEN_9309; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9311 = 8'h5f == io_state_in_8 ? 8'h91 : _GEN_9310; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9312 = 8'h60 == io_state_in_8 ? 8'h4d : _GEN_9311; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9313 = 8'h61 == io_state_in_8 ? 8'h44 : _GEN_9312; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9314 = 8'h62 == io_state_in_8 ? 8'h5f : _GEN_9313; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9315 = 8'h63 == io_state_in_8 ? 8'h56 : _GEN_9314; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9316 = 8'h64 == io_state_in_8 ? 8'h69 : _GEN_9315; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9317 = 8'h65 == io_state_in_8 ? 8'h60 : _GEN_9316; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9318 = 8'h66 == io_state_in_8 ? 8'h7b : _GEN_9317; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9319 = 8'h67 == io_state_in_8 ? 8'h72 : _GEN_9318; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9320 = 8'h68 == io_state_in_8 ? 8'h5 : _GEN_9319; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9321 = 8'h69 == io_state_in_8 ? 8'hc : _GEN_9320; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9322 = 8'h6a == io_state_in_8 ? 8'h17 : _GEN_9321; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9323 = 8'h6b == io_state_in_8 ? 8'h1e : _GEN_9322; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9324 = 8'h6c == io_state_in_8 ? 8'h21 : _GEN_9323; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9325 = 8'h6d == io_state_in_8 ? 8'h28 : _GEN_9324; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9326 = 8'h6e == io_state_in_8 ? 8'h33 : _GEN_9325; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9327 = 8'h6f == io_state_in_8 ? 8'h3a : _GEN_9326; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9328 = 8'h70 == io_state_in_8 ? 8'hdd : _GEN_9327; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9329 = 8'h71 == io_state_in_8 ? 8'hd4 : _GEN_9328; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9330 = 8'h72 == io_state_in_8 ? 8'hcf : _GEN_9329; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9331 = 8'h73 == io_state_in_8 ? 8'hc6 : _GEN_9330; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9332 = 8'h74 == io_state_in_8 ? 8'hf9 : _GEN_9331; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9333 = 8'h75 == io_state_in_8 ? 8'hf0 : _GEN_9332; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9334 = 8'h76 == io_state_in_8 ? 8'heb : _GEN_9333; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9335 = 8'h77 == io_state_in_8 ? 8'he2 : _GEN_9334; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9336 = 8'h78 == io_state_in_8 ? 8'h95 : _GEN_9335; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9337 = 8'h79 == io_state_in_8 ? 8'h9c : _GEN_9336; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9338 = 8'h7a == io_state_in_8 ? 8'h87 : _GEN_9337; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9339 = 8'h7b == io_state_in_8 ? 8'h8e : _GEN_9338; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9340 = 8'h7c == io_state_in_8 ? 8'hb1 : _GEN_9339; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9341 = 8'h7d == io_state_in_8 ? 8'hb8 : _GEN_9340; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9342 = 8'h7e == io_state_in_8 ? 8'ha3 : _GEN_9341; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9343 = 8'h7f == io_state_in_8 ? 8'haa : _GEN_9342; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9344 = 8'h80 == io_state_in_8 ? 8'hec : _GEN_9343; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9345 = 8'h81 == io_state_in_8 ? 8'he5 : _GEN_9344; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9346 = 8'h82 == io_state_in_8 ? 8'hfe : _GEN_9345; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9347 = 8'h83 == io_state_in_8 ? 8'hf7 : _GEN_9346; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9348 = 8'h84 == io_state_in_8 ? 8'hc8 : _GEN_9347; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9349 = 8'h85 == io_state_in_8 ? 8'hc1 : _GEN_9348; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9350 = 8'h86 == io_state_in_8 ? 8'hda : _GEN_9349; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9351 = 8'h87 == io_state_in_8 ? 8'hd3 : _GEN_9350; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9352 = 8'h88 == io_state_in_8 ? 8'ha4 : _GEN_9351; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9353 = 8'h89 == io_state_in_8 ? 8'had : _GEN_9352; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9354 = 8'h8a == io_state_in_8 ? 8'hb6 : _GEN_9353; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9355 = 8'h8b == io_state_in_8 ? 8'hbf : _GEN_9354; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9356 = 8'h8c == io_state_in_8 ? 8'h80 : _GEN_9355; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9357 = 8'h8d == io_state_in_8 ? 8'h89 : _GEN_9356; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9358 = 8'h8e == io_state_in_8 ? 8'h92 : _GEN_9357; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9359 = 8'h8f == io_state_in_8 ? 8'h9b : _GEN_9358; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9360 = 8'h90 == io_state_in_8 ? 8'h7c : _GEN_9359; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9361 = 8'h91 == io_state_in_8 ? 8'h75 : _GEN_9360; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9362 = 8'h92 == io_state_in_8 ? 8'h6e : _GEN_9361; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9363 = 8'h93 == io_state_in_8 ? 8'h67 : _GEN_9362; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9364 = 8'h94 == io_state_in_8 ? 8'h58 : _GEN_9363; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9365 = 8'h95 == io_state_in_8 ? 8'h51 : _GEN_9364; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9366 = 8'h96 == io_state_in_8 ? 8'h4a : _GEN_9365; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9367 = 8'h97 == io_state_in_8 ? 8'h43 : _GEN_9366; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9368 = 8'h98 == io_state_in_8 ? 8'h34 : _GEN_9367; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9369 = 8'h99 == io_state_in_8 ? 8'h3d : _GEN_9368; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9370 = 8'h9a == io_state_in_8 ? 8'h26 : _GEN_9369; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9371 = 8'h9b == io_state_in_8 ? 8'h2f : _GEN_9370; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9372 = 8'h9c == io_state_in_8 ? 8'h10 : _GEN_9371; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9373 = 8'h9d == io_state_in_8 ? 8'h19 : _GEN_9372; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9374 = 8'h9e == io_state_in_8 ? 8'h2 : _GEN_9373; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9375 = 8'h9f == io_state_in_8 ? 8'hb : _GEN_9374; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9376 = 8'ha0 == io_state_in_8 ? 8'hd7 : _GEN_9375; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9377 = 8'ha1 == io_state_in_8 ? 8'hde : _GEN_9376; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9378 = 8'ha2 == io_state_in_8 ? 8'hc5 : _GEN_9377; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9379 = 8'ha3 == io_state_in_8 ? 8'hcc : _GEN_9378; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9380 = 8'ha4 == io_state_in_8 ? 8'hf3 : _GEN_9379; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9381 = 8'ha5 == io_state_in_8 ? 8'hfa : _GEN_9380; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9382 = 8'ha6 == io_state_in_8 ? 8'he1 : _GEN_9381; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9383 = 8'ha7 == io_state_in_8 ? 8'he8 : _GEN_9382; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9384 = 8'ha8 == io_state_in_8 ? 8'h9f : _GEN_9383; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9385 = 8'ha9 == io_state_in_8 ? 8'h96 : _GEN_9384; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9386 = 8'haa == io_state_in_8 ? 8'h8d : _GEN_9385; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9387 = 8'hab == io_state_in_8 ? 8'h84 : _GEN_9386; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9388 = 8'hac == io_state_in_8 ? 8'hbb : _GEN_9387; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9389 = 8'had == io_state_in_8 ? 8'hb2 : _GEN_9388; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9390 = 8'hae == io_state_in_8 ? 8'ha9 : _GEN_9389; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9391 = 8'haf == io_state_in_8 ? 8'ha0 : _GEN_9390; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9392 = 8'hb0 == io_state_in_8 ? 8'h47 : _GEN_9391; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9393 = 8'hb1 == io_state_in_8 ? 8'h4e : _GEN_9392; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9394 = 8'hb2 == io_state_in_8 ? 8'h55 : _GEN_9393; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9395 = 8'hb3 == io_state_in_8 ? 8'h5c : _GEN_9394; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9396 = 8'hb4 == io_state_in_8 ? 8'h63 : _GEN_9395; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9397 = 8'hb5 == io_state_in_8 ? 8'h6a : _GEN_9396; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9398 = 8'hb6 == io_state_in_8 ? 8'h71 : _GEN_9397; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9399 = 8'hb7 == io_state_in_8 ? 8'h78 : _GEN_9398; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9400 = 8'hb8 == io_state_in_8 ? 8'hf : _GEN_9399; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9401 = 8'hb9 == io_state_in_8 ? 8'h6 : _GEN_9400; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9402 = 8'hba == io_state_in_8 ? 8'h1d : _GEN_9401; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9403 = 8'hbb == io_state_in_8 ? 8'h14 : _GEN_9402; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9404 = 8'hbc == io_state_in_8 ? 8'h2b : _GEN_9403; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9405 = 8'hbd == io_state_in_8 ? 8'h22 : _GEN_9404; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9406 = 8'hbe == io_state_in_8 ? 8'h39 : _GEN_9405; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9407 = 8'hbf == io_state_in_8 ? 8'h30 : _GEN_9406; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9408 = 8'hc0 == io_state_in_8 ? 8'h9a : _GEN_9407; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9409 = 8'hc1 == io_state_in_8 ? 8'h93 : _GEN_9408; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9410 = 8'hc2 == io_state_in_8 ? 8'h88 : _GEN_9409; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9411 = 8'hc3 == io_state_in_8 ? 8'h81 : _GEN_9410; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9412 = 8'hc4 == io_state_in_8 ? 8'hbe : _GEN_9411; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9413 = 8'hc5 == io_state_in_8 ? 8'hb7 : _GEN_9412; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9414 = 8'hc6 == io_state_in_8 ? 8'hac : _GEN_9413; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9415 = 8'hc7 == io_state_in_8 ? 8'ha5 : _GEN_9414; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9416 = 8'hc8 == io_state_in_8 ? 8'hd2 : _GEN_9415; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9417 = 8'hc9 == io_state_in_8 ? 8'hdb : _GEN_9416; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9418 = 8'hca == io_state_in_8 ? 8'hc0 : _GEN_9417; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9419 = 8'hcb == io_state_in_8 ? 8'hc9 : _GEN_9418; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9420 = 8'hcc == io_state_in_8 ? 8'hf6 : _GEN_9419; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9421 = 8'hcd == io_state_in_8 ? 8'hff : _GEN_9420; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9422 = 8'hce == io_state_in_8 ? 8'he4 : _GEN_9421; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9423 = 8'hcf == io_state_in_8 ? 8'hed : _GEN_9422; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9424 = 8'hd0 == io_state_in_8 ? 8'ha : _GEN_9423; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9425 = 8'hd1 == io_state_in_8 ? 8'h3 : _GEN_9424; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9426 = 8'hd2 == io_state_in_8 ? 8'h18 : _GEN_9425; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9427 = 8'hd3 == io_state_in_8 ? 8'h11 : _GEN_9426; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9428 = 8'hd4 == io_state_in_8 ? 8'h2e : _GEN_9427; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9429 = 8'hd5 == io_state_in_8 ? 8'h27 : _GEN_9428; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9430 = 8'hd6 == io_state_in_8 ? 8'h3c : _GEN_9429; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9431 = 8'hd7 == io_state_in_8 ? 8'h35 : _GEN_9430; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9432 = 8'hd8 == io_state_in_8 ? 8'h42 : _GEN_9431; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9433 = 8'hd9 == io_state_in_8 ? 8'h4b : _GEN_9432; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9434 = 8'hda == io_state_in_8 ? 8'h50 : _GEN_9433; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9435 = 8'hdb == io_state_in_8 ? 8'h59 : _GEN_9434; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9436 = 8'hdc == io_state_in_8 ? 8'h66 : _GEN_9435; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9437 = 8'hdd == io_state_in_8 ? 8'h6f : _GEN_9436; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9438 = 8'hde == io_state_in_8 ? 8'h74 : _GEN_9437; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9439 = 8'hdf == io_state_in_8 ? 8'h7d : _GEN_9438; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9440 = 8'he0 == io_state_in_8 ? 8'ha1 : _GEN_9439; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9441 = 8'he1 == io_state_in_8 ? 8'ha8 : _GEN_9440; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9442 = 8'he2 == io_state_in_8 ? 8'hb3 : _GEN_9441; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9443 = 8'he3 == io_state_in_8 ? 8'hba : _GEN_9442; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9444 = 8'he4 == io_state_in_8 ? 8'h85 : _GEN_9443; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9445 = 8'he5 == io_state_in_8 ? 8'h8c : _GEN_9444; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9446 = 8'he6 == io_state_in_8 ? 8'h97 : _GEN_9445; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9447 = 8'he7 == io_state_in_8 ? 8'h9e : _GEN_9446; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9448 = 8'he8 == io_state_in_8 ? 8'he9 : _GEN_9447; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9449 = 8'he9 == io_state_in_8 ? 8'he0 : _GEN_9448; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9450 = 8'hea == io_state_in_8 ? 8'hfb : _GEN_9449; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9451 = 8'heb == io_state_in_8 ? 8'hf2 : _GEN_9450; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9452 = 8'hec == io_state_in_8 ? 8'hcd : _GEN_9451; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9453 = 8'hed == io_state_in_8 ? 8'hc4 : _GEN_9452; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9454 = 8'hee == io_state_in_8 ? 8'hdf : _GEN_9453; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9455 = 8'hef == io_state_in_8 ? 8'hd6 : _GEN_9454; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9456 = 8'hf0 == io_state_in_8 ? 8'h31 : _GEN_9455; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9457 = 8'hf1 == io_state_in_8 ? 8'h38 : _GEN_9456; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9458 = 8'hf2 == io_state_in_8 ? 8'h23 : _GEN_9457; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9459 = 8'hf3 == io_state_in_8 ? 8'h2a : _GEN_9458; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9460 = 8'hf4 == io_state_in_8 ? 8'h15 : _GEN_9459; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9461 = 8'hf5 == io_state_in_8 ? 8'h1c : _GEN_9460; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9462 = 8'hf6 == io_state_in_8 ? 8'h7 : _GEN_9461; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9463 = 8'hf7 == io_state_in_8 ? 8'he : _GEN_9462; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9464 = 8'hf8 == io_state_in_8 ? 8'h79 : _GEN_9463; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9465 = 8'hf9 == io_state_in_8 ? 8'h70 : _GEN_9464; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9466 = 8'hfa == io_state_in_8 ? 8'h6b : _GEN_9465; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9467 = 8'hfb == io_state_in_8 ? 8'h62 : _GEN_9466; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9468 = 8'hfc == io_state_in_8 ? 8'h5d : _GEN_9467; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9469 = 8'hfd == io_state_in_8 ? 8'h54 : _GEN_9468; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9470 = 8'hfe == io_state_in_8 ? 8'h4f : _GEN_9469; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9471 = 8'hff == io_state_in_8 ? 8'h46 : _GEN_9470; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9473 = 8'h1 == io_state_in_9 ? 8'he : 8'h0; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9474 = 8'h2 == io_state_in_9 ? 8'h1c : _GEN_9473; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9475 = 8'h3 == io_state_in_9 ? 8'h12 : _GEN_9474; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9476 = 8'h4 == io_state_in_9 ? 8'h38 : _GEN_9475; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9477 = 8'h5 == io_state_in_9 ? 8'h36 : _GEN_9476; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9478 = 8'h6 == io_state_in_9 ? 8'h24 : _GEN_9477; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9479 = 8'h7 == io_state_in_9 ? 8'h2a : _GEN_9478; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9480 = 8'h8 == io_state_in_9 ? 8'h70 : _GEN_9479; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9481 = 8'h9 == io_state_in_9 ? 8'h7e : _GEN_9480; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9482 = 8'ha == io_state_in_9 ? 8'h6c : _GEN_9481; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9483 = 8'hb == io_state_in_9 ? 8'h62 : _GEN_9482; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9484 = 8'hc == io_state_in_9 ? 8'h48 : _GEN_9483; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9485 = 8'hd == io_state_in_9 ? 8'h46 : _GEN_9484; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9486 = 8'he == io_state_in_9 ? 8'h54 : _GEN_9485; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9487 = 8'hf == io_state_in_9 ? 8'h5a : _GEN_9486; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9488 = 8'h10 == io_state_in_9 ? 8'he0 : _GEN_9487; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9489 = 8'h11 == io_state_in_9 ? 8'hee : _GEN_9488; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9490 = 8'h12 == io_state_in_9 ? 8'hfc : _GEN_9489; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9491 = 8'h13 == io_state_in_9 ? 8'hf2 : _GEN_9490; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9492 = 8'h14 == io_state_in_9 ? 8'hd8 : _GEN_9491; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9493 = 8'h15 == io_state_in_9 ? 8'hd6 : _GEN_9492; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9494 = 8'h16 == io_state_in_9 ? 8'hc4 : _GEN_9493; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9495 = 8'h17 == io_state_in_9 ? 8'hca : _GEN_9494; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9496 = 8'h18 == io_state_in_9 ? 8'h90 : _GEN_9495; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9497 = 8'h19 == io_state_in_9 ? 8'h9e : _GEN_9496; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9498 = 8'h1a == io_state_in_9 ? 8'h8c : _GEN_9497; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9499 = 8'h1b == io_state_in_9 ? 8'h82 : _GEN_9498; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9500 = 8'h1c == io_state_in_9 ? 8'ha8 : _GEN_9499; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9501 = 8'h1d == io_state_in_9 ? 8'ha6 : _GEN_9500; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9502 = 8'h1e == io_state_in_9 ? 8'hb4 : _GEN_9501; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9503 = 8'h1f == io_state_in_9 ? 8'hba : _GEN_9502; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9504 = 8'h20 == io_state_in_9 ? 8'hdb : _GEN_9503; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9505 = 8'h21 == io_state_in_9 ? 8'hd5 : _GEN_9504; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9506 = 8'h22 == io_state_in_9 ? 8'hc7 : _GEN_9505; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9507 = 8'h23 == io_state_in_9 ? 8'hc9 : _GEN_9506; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9508 = 8'h24 == io_state_in_9 ? 8'he3 : _GEN_9507; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9509 = 8'h25 == io_state_in_9 ? 8'hed : _GEN_9508; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9510 = 8'h26 == io_state_in_9 ? 8'hff : _GEN_9509; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9511 = 8'h27 == io_state_in_9 ? 8'hf1 : _GEN_9510; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9512 = 8'h28 == io_state_in_9 ? 8'hab : _GEN_9511; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9513 = 8'h29 == io_state_in_9 ? 8'ha5 : _GEN_9512; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9514 = 8'h2a == io_state_in_9 ? 8'hb7 : _GEN_9513; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9515 = 8'h2b == io_state_in_9 ? 8'hb9 : _GEN_9514; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9516 = 8'h2c == io_state_in_9 ? 8'h93 : _GEN_9515; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9517 = 8'h2d == io_state_in_9 ? 8'h9d : _GEN_9516; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9518 = 8'h2e == io_state_in_9 ? 8'h8f : _GEN_9517; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9519 = 8'h2f == io_state_in_9 ? 8'h81 : _GEN_9518; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9520 = 8'h30 == io_state_in_9 ? 8'h3b : _GEN_9519; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9521 = 8'h31 == io_state_in_9 ? 8'h35 : _GEN_9520; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9522 = 8'h32 == io_state_in_9 ? 8'h27 : _GEN_9521; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9523 = 8'h33 == io_state_in_9 ? 8'h29 : _GEN_9522; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9524 = 8'h34 == io_state_in_9 ? 8'h3 : _GEN_9523; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9525 = 8'h35 == io_state_in_9 ? 8'hd : _GEN_9524; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9526 = 8'h36 == io_state_in_9 ? 8'h1f : _GEN_9525; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9527 = 8'h37 == io_state_in_9 ? 8'h11 : _GEN_9526; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9528 = 8'h38 == io_state_in_9 ? 8'h4b : _GEN_9527; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9529 = 8'h39 == io_state_in_9 ? 8'h45 : _GEN_9528; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9530 = 8'h3a == io_state_in_9 ? 8'h57 : _GEN_9529; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9531 = 8'h3b == io_state_in_9 ? 8'h59 : _GEN_9530; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9532 = 8'h3c == io_state_in_9 ? 8'h73 : _GEN_9531; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9533 = 8'h3d == io_state_in_9 ? 8'h7d : _GEN_9532; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9534 = 8'h3e == io_state_in_9 ? 8'h6f : _GEN_9533; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9535 = 8'h3f == io_state_in_9 ? 8'h61 : _GEN_9534; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9536 = 8'h40 == io_state_in_9 ? 8'had : _GEN_9535; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9537 = 8'h41 == io_state_in_9 ? 8'ha3 : _GEN_9536; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9538 = 8'h42 == io_state_in_9 ? 8'hb1 : _GEN_9537; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9539 = 8'h43 == io_state_in_9 ? 8'hbf : _GEN_9538; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9540 = 8'h44 == io_state_in_9 ? 8'h95 : _GEN_9539; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9541 = 8'h45 == io_state_in_9 ? 8'h9b : _GEN_9540; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9542 = 8'h46 == io_state_in_9 ? 8'h89 : _GEN_9541; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9543 = 8'h47 == io_state_in_9 ? 8'h87 : _GEN_9542; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9544 = 8'h48 == io_state_in_9 ? 8'hdd : _GEN_9543; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9545 = 8'h49 == io_state_in_9 ? 8'hd3 : _GEN_9544; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9546 = 8'h4a == io_state_in_9 ? 8'hc1 : _GEN_9545; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9547 = 8'h4b == io_state_in_9 ? 8'hcf : _GEN_9546; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9548 = 8'h4c == io_state_in_9 ? 8'he5 : _GEN_9547; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9549 = 8'h4d == io_state_in_9 ? 8'heb : _GEN_9548; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9550 = 8'h4e == io_state_in_9 ? 8'hf9 : _GEN_9549; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9551 = 8'h4f == io_state_in_9 ? 8'hf7 : _GEN_9550; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9552 = 8'h50 == io_state_in_9 ? 8'h4d : _GEN_9551; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9553 = 8'h51 == io_state_in_9 ? 8'h43 : _GEN_9552; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9554 = 8'h52 == io_state_in_9 ? 8'h51 : _GEN_9553; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9555 = 8'h53 == io_state_in_9 ? 8'h5f : _GEN_9554; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9556 = 8'h54 == io_state_in_9 ? 8'h75 : _GEN_9555; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9557 = 8'h55 == io_state_in_9 ? 8'h7b : _GEN_9556; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9558 = 8'h56 == io_state_in_9 ? 8'h69 : _GEN_9557; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9559 = 8'h57 == io_state_in_9 ? 8'h67 : _GEN_9558; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9560 = 8'h58 == io_state_in_9 ? 8'h3d : _GEN_9559; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9561 = 8'h59 == io_state_in_9 ? 8'h33 : _GEN_9560; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9562 = 8'h5a == io_state_in_9 ? 8'h21 : _GEN_9561; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9563 = 8'h5b == io_state_in_9 ? 8'h2f : _GEN_9562; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9564 = 8'h5c == io_state_in_9 ? 8'h5 : _GEN_9563; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9565 = 8'h5d == io_state_in_9 ? 8'hb : _GEN_9564; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9566 = 8'h5e == io_state_in_9 ? 8'h19 : _GEN_9565; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9567 = 8'h5f == io_state_in_9 ? 8'h17 : _GEN_9566; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9568 = 8'h60 == io_state_in_9 ? 8'h76 : _GEN_9567; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9569 = 8'h61 == io_state_in_9 ? 8'h78 : _GEN_9568; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9570 = 8'h62 == io_state_in_9 ? 8'h6a : _GEN_9569; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9571 = 8'h63 == io_state_in_9 ? 8'h64 : _GEN_9570; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9572 = 8'h64 == io_state_in_9 ? 8'h4e : _GEN_9571; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9573 = 8'h65 == io_state_in_9 ? 8'h40 : _GEN_9572; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9574 = 8'h66 == io_state_in_9 ? 8'h52 : _GEN_9573; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9575 = 8'h67 == io_state_in_9 ? 8'h5c : _GEN_9574; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9576 = 8'h68 == io_state_in_9 ? 8'h6 : _GEN_9575; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9577 = 8'h69 == io_state_in_9 ? 8'h8 : _GEN_9576; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9578 = 8'h6a == io_state_in_9 ? 8'h1a : _GEN_9577; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9579 = 8'h6b == io_state_in_9 ? 8'h14 : _GEN_9578; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9580 = 8'h6c == io_state_in_9 ? 8'h3e : _GEN_9579; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9581 = 8'h6d == io_state_in_9 ? 8'h30 : _GEN_9580; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9582 = 8'h6e == io_state_in_9 ? 8'h22 : _GEN_9581; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9583 = 8'h6f == io_state_in_9 ? 8'h2c : _GEN_9582; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9584 = 8'h70 == io_state_in_9 ? 8'h96 : _GEN_9583; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9585 = 8'h71 == io_state_in_9 ? 8'h98 : _GEN_9584; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9586 = 8'h72 == io_state_in_9 ? 8'h8a : _GEN_9585; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9587 = 8'h73 == io_state_in_9 ? 8'h84 : _GEN_9586; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9588 = 8'h74 == io_state_in_9 ? 8'hae : _GEN_9587; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9589 = 8'h75 == io_state_in_9 ? 8'ha0 : _GEN_9588; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9590 = 8'h76 == io_state_in_9 ? 8'hb2 : _GEN_9589; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9591 = 8'h77 == io_state_in_9 ? 8'hbc : _GEN_9590; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9592 = 8'h78 == io_state_in_9 ? 8'he6 : _GEN_9591; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9593 = 8'h79 == io_state_in_9 ? 8'he8 : _GEN_9592; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9594 = 8'h7a == io_state_in_9 ? 8'hfa : _GEN_9593; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9595 = 8'h7b == io_state_in_9 ? 8'hf4 : _GEN_9594; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9596 = 8'h7c == io_state_in_9 ? 8'hde : _GEN_9595; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9597 = 8'h7d == io_state_in_9 ? 8'hd0 : _GEN_9596; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9598 = 8'h7e == io_state_in_9 ? 8'hc2 : _GEN_9597; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9599 = 8'h7f == io_state_in_9 ? 8'hcc : _GEN_9598; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9600 = 8'h80 == io_state_in_9 ? 8'h41 : _GEN_9599; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9601 = 8'h81 == io_state_in_9 ? 8'h4f : _GEN_9600; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9602 = 8'h82 == io_state_in_9 ? 8'h5d : _GEN_9601; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9603 = 8'h83 == io_state_in_9 ? 8'h53 : _GEN_9602; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9604 = 8'h84 == io_state_in_9 ? 8'h79 : _GEN_9603; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9605 = 8'h85 == io_state_in_9 ? 8'h77 : _GEN_9604; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9606 = 8'h86 == io_state_in_9 ? 8'h65 : _GEN_9605; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9607 = 8'h87 == io_state_in_9 ? 8'h6b : _GEN_9606; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9608 = 8'h88 == io_state_in_9 ? 8'h31 : _GEN_9607; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9609 = 8'h89 == io_state_in_9 ? 8'h3f : _GEN_9608; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9610 = 8'h8a == io_state_in_9 ? 8'h2d : _GEN_9609; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9611 = 8'h8b == io_state_in_9 ? 8'h23 : _GEN_9610; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9612 = 8'h8c == io_state_in_9 ? 8'h9 : _GEN_9611; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9613 = 8'h8d == io_state_in_9 ? 8'h7 : _GEN_9612; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9614 = 8'h8e == io_state_in_9 ? 8'h15 : _GEN_9613; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9615 = 8'h8f == io_state_in_9 ? 8'h1b : _GEN_9614; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9616 = 8'h90 == io_state_in_9 ? 8'ha1 : _GEN_9615; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9617 = 8'h91 == io_state_in_9 ? 8'haf : _GEN_9616; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9618 = 8'h92 == io_state_in_9 ? 8'hbd : _GEN_9617; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9619 = 8'h93 == io_state_in_9 ? 8'hb3 : _GEN_9618; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9620 = 8'h94 == io_state_in_9 ? 8'h99 : _GEN_9619; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9621 = 8'h95 == io_state_in_9 ? 8'h97 : _GEN_9620; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9622 = 8'h96 == io_state_in_9 ? 8'h85 : _GEN_9621; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9623 = 8'h97 == io_state_in_9 ? 8'h8b : _GEN_9622; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9624 = 8'h98 == io_state_in_9 ? 8'hd1 : _GEN_9623; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9625 = 8'h99 == io_state_in_9 ? 8'hdf : _GEN_9624; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9626 = 8'h9a == io_state_in_9 ? 8'hcd : _GEN_9625; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9627 = 8'h9b == io_state_in_9 ? 8'hc3 : _GEN_9626; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9628 = 8'h9c == io_state_in_9 ? 8'he9 : _GEN_9627; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9629 = 8'h9d == io_state_in_9 ? 8'he7 : _GEN_9628; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9630 = 8'h9e == io_state_in_9 ? 8'hf5 : _GEN_9629; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9631 = 8'h9f == io_state_in_9 ? 8'hfb : _GEN_9630; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9632 = 8'ha0 == io_state_in_9 ? 8'h9a : _GEN_9631; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9633 = 8'ha1 == io_state_in_9 ? 8'h94 : _GEN_9632; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9634 = 8'ha2 == io_state_in_9 ? 8'h86 : _GEN_9633; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9635 = 8'ha3 == io_state_in_9 ? 8'h88 : _GEN_9634; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9636 = 8'ha4 == io_state_in_9 ? 8'ha2 : _GEN_9635; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9637 = 8'ha5 == io_state_in_9 ? 8'hac : _GEN_9636; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9638 = 8'ha6 == io_state_in_9 ? 8'hbe : _GEN_9637; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9639 = 8'ha7 == io_state_in_9 ? 8'hb0 : _GEN_9638; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9640 = 8'ha8 == io_state_in_9 ? 8'hea : _GEN_9639; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9641 = 8'ha9 == io_state_in_9 ? 8'he4 : _GEN_9640; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9642 = 8'haa == io_state_in_9 ? 8'hf6 : _GEN_9641; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9643 = 8'hab == io_state_in_9 ? 8'hf8 : _GEN_9642; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9644 = 8'hac == io_state_in_9 ? 8'hd2 : _GEN_9643; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9645 = 8'had == io_state_in_9 ? 8'hdc : _GEN_9644; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9646 = 8'hae == io_state_in_9 ? 8'hce : _GEN_9645; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9647 = 8'haf == io_state_in_9 ? 8'hc0 : _GEN_9646; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9648 = 8'hb0 == io_state_in_9 ? 8'h7a : _GEN_9647; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9649 = 8'hb1 == io_state_in_9 ? 8'h74 : _GEN_9648; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9650 = 8'hb2 == io_state_in_9 ? 8'h66 : _GEN_9649; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9651 = 8'hb3 == io_state_in_9 ? 8'h68 : _GEN_9650; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9652 = 8'hb4 == io_state_in_9 ? 8'h42 : _GEN_9651; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9653 = 8'hb5 == io_state_in_9 ? 8'h4c : _GEN_9652; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9654 = 8'hb6 == io_state_in_9 ? 8'h5e : _GEN_9653; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9655 = 8'hb7 == io_state_in_9 ? 8'h50 : _GEN_9654; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9656 = 8'hb8 == io_state_in_9 ? 8'ha : _GEN_9655; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9657 = 8'hb9 == io_state_in_9 ? 8'h4 : _GEN_9656; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9658 = 8'hba == io_state_in_9 ? 8'h16 : _GEN_9657; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9659 = 8'hbb == io_state_in_9 ? 8'h18 : _GEN_9658; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9660 = 8'hbc == io_state_in_9 ? 8'h32 : _GEN_9659; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9661 = 8'hbd == io_state_in_9 ? 8'h3c : _GEN_9660; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9662 = 8'hbe == io_state_in_9 ? 8'h2e : _GEN_9661; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9663 = 8'hbf == io_state_in_9 ? 8'h20 : _GEN_9662; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9664 = 8'hc0 == io_state_in_9 ? 8'hec : _GEN_9663; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9665 = 8'hc1 == io_state_in_9 ? 8'he2 : _GEN_9664; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9666 = 8'hc2 == io_state_in_9 ? 8'hf0 : _GEN_9665; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9667 = 8'hc3 == io_state_in_9 ? 8'hfe : _GEN_9666; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9668 = 8'hc4 == io_state_in_9 ? 8'hd4 : _GEN_9667; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9669 = 8'hc5 == io_state_in_9 ? 8'hda : _GEN_9668; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9670 = 8'hc6 == io_state_in_9 ? 8'hc8 : _GEN_9669; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9671 = 8'hc7 == io_state_in_9 ? 8'hc6 : _GEN_9670; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9672 = 8'hc8 == io_state_in_9 ? 8'h9c : _GEN_9671; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9673 = 8'hc9 == io_state_in_9 ? 8'h92 : _GEN_9672; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9674 = 8'hca == io_state_in_9 ? 8'h80 : _GEN_9673; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9675 = 8'hcb == io_state_in_9 ? 8'h8e : _GEN_9674; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9676 = 8'hcc == io_state_in_9 ? 8'ha4 : _GEN_9675; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9677 = 8'hcd == io_state_in_9 ? 8'haa : _GEN_9676; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9678 = 8'hce == io_state_in_9 ? 8'hb8 : _GEN_9677; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9679 = 8'hcf == io_state_in_9 ? 8'hb6 : _GEN_9678; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9680 = 8'hd0 == io_state_in_9 ? 8'hc : _GEN_9679; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9681 = 8'hd1 == io_state_in_9 ? 8'h2 : _GEN_9680; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9682 = 8'hd2 == io_state_in_9 ? 8'h10 : _GEN_9681; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9683 = 8'hd3 == io_state_in_9 ? 8'h1e : _GEN_9682; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9684 = 8'hd4 == io_state_in_9 ? 8'h34 : _GEN_9683; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9685 = 8'hd5 == io_state_in_9 ? 8'h3a : _GEN_9684; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9686 = 8'hd6 == io_state_in_9 ? 8'h28 : _GEN_9685; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9687 = 8'hd7 == io_state_in_9 ? 8'h26 : _GEN_9686; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9688 = 8'hd8 == io_state_in_9 ? 8'h7c : _GEN_9687; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9689 = 8'hd9 == io_state_in_9 ? 8'h72 : _GEN_9688; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9690 = 8'hda == io_state_in_9 ? 8'h60 : _GEN_9689; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9691 = 8'hdb == io_state_in_9 ? 8'h6e : _GEN_9690; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9692 = 8'hdc == io_state_in_9 ? 8'h44 : _GEN_9691; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9693 = 8'hdd == io_state_in_9 ? 8'h4a : _GEN_9692; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9694 = 8'hde == io_state_in_9 ? 8'h58 : _GEN_9693; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9695 = 8'hdf == io_state_in_9 ? 8'h56 : _GEN_9694; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9696 = 8'he0 == io_state_in_9 ? 8'h37 : _GEN_9695; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9697 = 8'he1 == io_state_in_9 ? 8'h39 : _GEN_9696; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9698 = 8'he2 == io_state_in_9 ? 8'h2b : _GEN_9697; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9699 = 8'he3 == io_state_in_9 ? 8'h25 : _GEN_9698; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9700 = 8'he4 == io_state_in_9 ? 8'hf : _GEN_9699; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9701 = 8'he5 == io_state_in_9 ? 8'h1 : _GEN_9700; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9702 = 8'he6 == io_state_in_9 ? 8'h13 : _GEN_9701; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9703 = 8'he7 == io_state_in_9 ? 8'h1d : _GEN_9702; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9704 = 8'he8 == io_state_in_9 ? 8'h47 : _GEN_9703; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9705 = 8'he9 == io_state_in_9 ? 8'h49 : _GEN_9704; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9706 = 8'hea == io_state_in_9 ? 8'h5b : _GEN_9705; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9707 = 8'heb == io_state_in_9 ? 8'h55 : _GEN_9706; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9708 = 8'hec == io_state_in_9 ? 8'h7f : _GEN_9707; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9709 = 8'hed == io_state_in_9 ? 8'h71 : _GEN_9708; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9710 = 8'hee == io_state_in_9 ? 8'h63 : _GEN_9709; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9711 = 8'hef == io_state_in_9 ? 8'h6d : _GEN_9710; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9712 = 8'hf0 == io_state_in_9 ? 8'hd7 : _GEN_9711; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9713 = 8'hf1 == io_state_in_9 ? 8'hd9 : _GEN_9712; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9714 = 8'hf2 == io_state_in_9 ? 8'hcb : _GEN_9713; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9715 = 8'hf3 == io_state_in_9 ? 8'hc5 : _GEN_9714; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9716 = 8'hf4 == io_state_in_9 ? 8'hef : _GEN_9715; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9717 = 8'hf5 == io_state_in_9 ? 8'he1 : _GEN_9716; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9718 = 8'hf6 == io_state_in_9 ? 8'hf3 : _GEN_9717; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9719 = 8'hf7 == io_state_in_9 ? 8'hfd : _GEN_9718; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9720 = 8'hf8 == io_state_in_9 ? 8'ha7 : _GEN_9719; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9721 = 8'hf9 == io_state_in_9 ? 8'ha9 : _GEN_9720; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9722 = 8'hfa == io_state_in_9 ? 8'hbb : _GEN_9721; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9723 = 8'hfb == io_state_in_9 ? 8'hb5 : _GEN_9722; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9724 = 8'hfc == io_state_in_9 ? 8'h9f : _GEN_9723; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9725 = 8'hfd == io_state_in_9 ? 8'h91 : _GEN_9724; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9726 = 8'hfe == io_state_in_9 ? 8'h83 : _GEN_9725; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _GEN_9727 = 8'hff == io_state_in_9 ? 8'h8d : _GEN_9726; // @[InvMixColumns.scala 137:{41,41}]
  wire [7:0] _tmp_state_9_T = _GEN_9471 ^ _GEN_9727; // @[InvMixColumns.scala 137:41]
  wire [7:0] _GEN_9729 = 8'h1 == io_state_in_10 ? 8'hb : 8'h0; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9730 = 8'h2 == io_state_in_10 ? 8'h16 : _GEN_9729; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9731 = 8'h3 == io_state_in_10 ? 8'h1d : _GEN_9730; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9732 = 8'h4 == io_state_in_10 ? 8'h2c : _GEN_9731; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9733 = 8'h5 == io_state_in_10 ? 8'h27 : _GEN_9732; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9734 = 8'h6 == io_state_in_10 ? 8'h3a : _GEN_9733; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9735 = 8'h7 == io_state_in_10 ? 8'h31 : _GEN_9734; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9736 = 8'h8 == io_state_in_10 ? 8'h58 : _GEN_9735; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9737 = 8'h9 == io_state_in_10 ? 8'h53 : _GEN_9736; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9738 = 8'ha == io_state_in_10 ? 8'h4e : _GEN_9737; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9739 = 8'hb == io_state_in_10 ? 8'h45 : _GEN_9738; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9740 = 8'hc == io_state_in_10 ? 8'h74 : _GEN_9739; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9741 = 8'hd == io_state_in_10 ? 8'h7f : _GEN_9740; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9742 = 8'he == io_state_in_10 ? 8'h62 : _GEN_9741; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9743 = 8'hf == io_state_in_10 ? 8'h69 : _GEN_9742; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9744 = 8'h10 == io_state_in_10 ? 8'hb0 : _GEN_9743; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9745 = 8'h11 == io_state_in_10 ? 8'hbb : _GEN_9744; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9746 = 8'h12 == io_state_in_10 ? 8'ha6 : _GEN_9745; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9747 = 8'h13 == io_state_in_10 ? 8'had : _GEN_9746; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9748 = 8'h14 == io_state_in_10 ? 8'h9c : _GEN_9747; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9749 = 8'h15 == io_state_in_10 ? 8'h97 : _GEN_9748; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9750 = 8'h16 == io_state_in_10 ? 8'h8a : _GEN_9749; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9751 = 8'h17 == io_state_in_10 ? 8'h81 : _GEN_9750; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9752 = 8'h18 == io_state_in_10 ? 8'he8 : _GEN_9751; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9753 = 8'h19 == io_state_in_10 ? 8'he3 : _GEN_9752; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9754 = 8'h1a == io_state_in_10 ? 8'hfe : _GEN_9753; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9755 = 8'h1b == io_state_in_10 ? 8'hf5 : _GEN_9754; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9756 = 8'h1c == io_state_in_10 ? 8'hc4 : _GEN_9755; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9757 = 8'h1d == io_state_in_10 ? 8'hcf : _GEN_9756; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9758 = 8'h1e == io_state_in_10 ? 8'hd2 : _GEN_9757; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9759 = 8'h1f == io_state_in_10 ? 8'hd9 : _GEN_9758; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9760 = 8'h20 == io_state_in_10 ? 8'h7b : _GEN_9759; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9761 = 8'h21 == io_state_in_10 ? 8'h70 : _GEN_9760; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9762 = 8'h22 == io_state_in_10 ? 8'h6d : _GEN_9761; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9763 = 8'h23 == io_state_in_10 ? 8'h66 : _GEN_9762; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9764 = 8'h24 == io_state_in_10 ? 8'h57 : _GEN_9763; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9765 = 8'h25 == io_state_in_10 ? 8'h5c : _GEN_9764; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9766 = 8'h26 == io_state_in_10 ? 8'h41 : _GEN_9765; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9767 = 8'h27 == io_state_in_10 ? 8'h4a : _GEN_9766; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9768 = 8'h28 == io_state_in_10 ? 8'h23 : _GEN_9767; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9769 = 8'h29 == io_state_in_10 ? 8'h28 : _GEN_9768; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9770 = 8'h2a == io_state_in_10 ? 8'h35 : _GEN_9769; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9771 = 8'h2b == io_state_in_10 ? 8'h3e : _GEN_9770; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9772 = 8'h2c == io_state_in_10 ? 8'hf : _GEN_9771; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9773 = 8'h2d == io_state_in_10 ? 8'h4 : _GEN_9772; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9774 = 8'h2e == io_state_in_10 ? 8'h19 : _GEN_9773; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9775 = 8'h2f == io_state_in_10 ? 8'h12 : _GEN_9774; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9776 = 8'h30 == io_state_in_10 ? 8'hcb : _GEN_9775; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9777 = 8'h31 == io_state_in_10 ? 8'hc0 : _GEN_9776; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9778 = 8'h32 == io_state_in_10 ? 8'hdd : _GEN_9777; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9779 = 8'h33 == io_state_in_10 ? 8'hd6 : _GEN_9778; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9780 = 8'h34 == io_state_in_10 ? 8'he7 : _GEN_9779; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9781 = 8'h35 == io_state_in_10 ? 8'hec : _GEN_9780; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9782 = 8'h36 == io_state_in_10 ? 8'hf1 : _GEN_9781; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9783 = 8'h37 == io_state_in_10 ? 8'hfa : _GEN_9782; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9784 = 8'h38 == io_state_in_10 ? 8'h93 : _GEN_9783; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9785 = 8'h39 == io_state_in_10 ? 8'h98 : _GEN_9784; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9786 = 8'h3a == io_state_in_10 ? 8'h85 : _GEN_9785; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9787 = 8'h3b == io_state_in_10 ? 8'h8e : _GEN_9786; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9788 = 8'h3c == io_state_in_10 ? 8'hbf : _GEN_9787; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9789 = 8'h3d == io_state_in_10 ? 8'hb4 : _GEN_9788; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9790 = 8'h3e == io_state_in_10 ? 8'ha9 : _GEN_9789; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9791 = 8'h3f == io_state_in_10 ? 8'ha2 : _GEN_9790; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9792 = 8'h40 == io_state_in_10 ? 8'hf6 : _GEN_9791; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9793 = 8'h41 == io_state_in_10 ? 8'hfd : _GEN_9792; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9794 = 8'h42 == io_state_in_10 ? 8'he0 : _GEN_9793; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9795 = 8'h43 == io_state_in_10 ? 8'heb : _GEN_9794; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9796 = 8'h44 == io_state_in_10 ? 8'hda : _GEN_9795; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9797 = 8'h45 == io_state_in_10 ? 8'hd1 : _GEN_9796; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9798 = 8'h46 == io_state_in_10 ? 8'hcc : _GEN_9797; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9799 = 8'h47 == io_state_in_10 ? 8'hc7 : _GEN_9798; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9800 = 8'h48 == io_state_in_10 ? 8'hae : _GEN_9799; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9801 = 8'h49 == io_state_in_10 ? 8'ha5 : _GEN_9800; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9802 = 8'h4a == io_state_in_10 ? 8'hb8 : _GEN_9801; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9803 = 8'h4b == io_state_in_10 ? 8'hb3 : _GEN_9802; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9804 = 8'h4c == io_state_in_10 ? 8'h82 : _GEN_9803; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9805 = 8'h4d == io_state_in_10 ? 8'h89 : _GEN_9804; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9806 = 8'h4e == io_state_in_10 ? 8'h94 : _GEN_9805; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9807 = 8'h4f == io_state_in_10 ? 8'h9f : _GEN_9806; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9808 = 8'h50 == io_state_in_10 ? 8'h46 : _GEN_9807; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9809 = 8'h51 == io_state_in_10 ? 8'h4d : _GEN_9808; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9810 = 8'h52 == io_state_in_10 ? 8'h50 : _GEN_9809; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9811 = 8'h53 == io_state_in_10 ? 8'h5b : _GEN_9810; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9812 = 8'h54 == io_state_in_10 ? 8'h6a : _GEN_9811; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9813 = 8'h55 == io_state_in_10 ? 8'h61 : _GEN_9812; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9814 = 8'h56 == io_state_in_10 ? 8'h7c : _GEN_9813; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9815 = 8'h57 == io_state_in_10 ? 8'h77 : _GEN_9814; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9816 = 8'h58 == io_state_in_10 ? 8'h1e : _GEN_9815; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9817 = 8'h59 == io_state_in_10 ? 8'h15 : _GEN_9816; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9818 = 8'h5a == io_state_in_10 ? 8'h8 : _GEN_9817; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9819 = 8'h5b == io_state_in_10 ? 8'h3 : _GEN_9818; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9820 = 8'h5c == io_state_in_10 ? 8'h32 : _GEN_9819; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9821 = 8'h5d == io_state_in_10 ? 8'h39 : _GEN_9820; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9822 = 8'h5e == io_state_in_10 ? 8'h24 : _GEN_9821; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9823 = 8'h5f == io_state_in_10 ? 8'h2f : _GEN_9822; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9824 = 8'h60 == io_state_in_10 ? 8'h8d : _GEN_9823; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9825 = 8'h61 == io_state_in_10 ? 8'h86 : _GEN_9824; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9826 = 8'h62 == io_state_in_10 ? 8'h9b : _GEN_9825; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9827 = 8'h63 == io_state_in_10 ? 8'h90 : _GEN_9826; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9828 = 8'h64 == io_state_in_10 ? 8'ha1 : _GEN_9827; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9829 = 8'h65 == io_state_in_10 ? 8'haa : _GEN_9828; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9830 = 8'h66 == io_state_in_10 ? 8'hb7 : _GEN_9829; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9831 = 8'h67 == io_state_in_10 ? 8'hbc : _GEN_9830; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9832 = 8'h68 == io_state_in_10 ? 8'hd5 : _GEN_9831; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9833 = 8'h69 == io_state_in_10 ? 8'hde : _GEN_9832; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9834 = 8'h6a == io_state_in_10 ? 8'hc3 : _GEN_9833; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9835 = 8'h6b == io_state_in_10 ? 8'hc8 : _GEN_9834; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9836 = 8'h6c == io_state_in_10 ? 8'hf9 : _GEN_9835; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9837 = 8'h6d == io_state_in_10 ? 8'hf2 : _GEN_9836; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9838 = 8'h6e == io_state_in_10 ? 8'hef : _GEN_9837; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9839 = 8'h6f == io_state_in_10 ? 8'he4 : _GEN_9838; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9840 = 8'h70 == io_state_in_10 ? 8'h3d : _GEN_9839; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9841 = 8'h71 == io_state_in_10 ? 8'h36 : _GEN_9840; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9842 = 8'h72 == io_state_in_10 ? 8'h2b : _GEN_9841; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9843 = 8'h73 == io_state_in_10 ? 8'h20 : _GEN_9842; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9844 = 8'h74 == io_state_in_10 ? 8'h11 : _GEN_9843; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9845 = 8'h75 == io_state_in_10 ? 8'h1a : _GEN_9844; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9846 = 8'h76 == io_state_in_10 ? 8'h7 : _GEN_9845; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9847 = 8'h77 == io_state_in_10 ? 8'hc : _GEN_9846; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9848 = 8'h78 == io_state_in_10 ? 8'h65 : _GEN_9847; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9849 = 8'h79 == io_state_in_10 ? 8'h6e : _GEN_9848; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9850 = 8'h7a == io_state_in_10 ? 8'h73 : _GEN_9849; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9851 = 8'h7b == io_state_in_10 ? 8'h78 : _GEN_9850; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9852 = 8'h7c == io_state_in_10 ? 8'h49 : _GEN_9851; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9853 = 8'h7d == io_state_in_10 ? 8'h42 : _GEN_9852; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9854 = 8'h7e == io_state_in_10 ? 8'h5f : _GEN_9853; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9855 = 8'h7f == io_state_in_10 ? 8'h54 : _GEN_9854; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9856 = 8'h80 == io_state_in_10 ? 8'hf7 : _GEN_9855; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9857 = 8'h81 == io_state_in_10 ? 8'hfc : _GEN_9856; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9858 = 8'h82 == io_state_in_10 ? 8'he1 : _GEN_9857; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9859 = 8'h83 == io_state_in_10 ? 8'hea : _GEN_9858; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9860 = 8'h84 == io_state_in_10 ? 8'hdb : _GEN_9859; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9861 = 8'h85 == io_state_in_10 ? 8'hd0 : _GEN_9860; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9862 = 8'h86 == io_state_in_10 ? 8'hcd : _GEN_9861; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9863 = 8'h87 == io_state_in_10 ? 8'hc6 : _GEN_9862; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9864 = 8'h88 == io_state_in_10 ? 8'haf : _GEN_9863; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9865 = 8'h89 == io_state_in_10 ? 8'ha4 : _GEN_9864; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9866 = 8'h8a == io_state_in_10 ? 8'hb9 : _GEN_9865; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9867 = 8'h8b == io_state_in_10 ? 8'hb2 : _GEN_9866; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9868 = 8'h8c == io_state_in_10 ? 8'h83 : _GEN_9867; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9869 = 8'h8d == io_state_in_10 ? 8'h88 : _GEN_9868; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9870 = 8'h8e == io_state_in_10 ? 8'h95 : _GEN_9869; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9871 = 8'h8f == io_state_in_10 ? 8'h9e : _GEN_9870; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9872 = 8'h90 == io_state_in_10 ? 8'h47 : _GEN_9871; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9873 = 8'h91 == io_state_in_10 ? 8'h4c : _GEN_9872; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9874 = 8'h92 == io_state_in_10 ? 8'h51 : _GEN_9873; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9875 = 8'h93 == io_state_in_10 ? 8'h5a : _GEN_9874; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9876 = 8'h94 == io_state_in_10 ? 8'h6b : _GEN_9875; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9877 = 8'h95 == io_state_in_10 ? 8'h60 : _GEN_9876; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9878 = 8'h96 == io_state_in_10 ? 8'h7d : _GEN_9877; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9879 = 8'h97 == io_state_in_10 ? 8'h76 : _GEN_9878; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9880 = 8'h98 == io_state_in_10 ? 8'h1f : _GEN_9879; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9881 = 8'h99 == io_state_in_10 ? 8'h14 : _GEN_9880; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9882 = 8'h9a == io_state_in_10 ? 8'h9 : _GEN_9881; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9883 = 8'h9b == io_state_in_10 ? 8'h2 : _GEN_9882; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9884 = 8'h9c == io_state_in_10 ? 8'h33 : _GEN_9883; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9885 = 8'h9d == io_state_in_10 ? 8'h38 : _GEN_9884; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9886 = 8'h9e == io_state_in_10 ? 8'h25 : _GEN_9885; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9887 = 8'h9f == io_state_in_10 ? 8'h2e : _GEN_9886; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9888 = 8'ha0 == io_state_in_10 ? 8'h8c : _GEN_9887; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9889 = 8'ha1 == io_state_in_10 ? 8'h87 : _GEN_9888; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9890 = 8'ha2 == io_state_in_10 ? 8'h9a : _GEN_9889; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9891 = 8'ha3 == io_state_in_10 ? 8'h91 : _GEN_9890; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9892 = 8'ha4 == io_state_in_10 ? 8'ha0 : _GEN_9891; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9893 = 8'ha5 == io_state_in_10 ? 8'hab : _GEN_9892; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9894 = 8'ha6 == io_state_in_10 ? 8'hb6 : _GEN_9893; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9895 = 8'ha7 == io_state_in_10 ? 8'hbd : _GEN_9894; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9896 = 8'ha8 == io_state_in_10 ? 8'hd4 : _GEN_9895; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9897 = 8'ha9 == io_state_in_10 ? 8'hdf : _GEN_9896; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9898 = 8'haa == io_state_in_10 ? 8'hc2 : _GEN_9897; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9899 = 8'hab == io_state_in_10 ? 8'hc9 : _GEN_9898; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9900 = 8'hac == io_state_in_10 ? 8'hf8 : _GEN_9899; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9901 = 8'had == io_state_in_10 ? 8'hf3 : _GEN_9900; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9902 = 8'hae == io_state_in_10 ? 8'hee : _GEN_9901; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9903 = 8'haf == io_state_in_10 ? 8'he5 : _GEN_9902; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9904 = 8'hb0 == io_state_in_10 ? 8'h3c : _GEN_9903; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9905 = 8'hb1 == io_state_in_10 ? 8'h37 : _GEN_9904; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9906 = 8'hb2 == io_state_in_10 ? 8'h2a : _GEN_9905; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9907 = 8'hb3 == io_state_in_10 ? 8'h21 : _GEN_9906; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9908 = 8'hb4 == io_state_in_10 ? 8'h10 : _GEN_9907; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9909 = 8'hb5 == io_state_in_10 ? 8'h1b : _GEN_9908; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9910 = 8'hb6 == io_state_in_10 ? 8'h6 : _GEN_9909; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9911 = 8'hb7 == io_state_in_10 ? 8'hd : _GEN_9910; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9912 = 8'hb8 == io_state_in_10 ? 8'h64 : _GEN_9911; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9913 = 8'hb9 == io_state_in_10 ? 8'h6f : _GEN_9912; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9914 = 8'hba == io_state_in_10 ? 8'h72 : _GEN_9913; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9915 = 8'hbb == io_state_in_10 ? 8'h79 : _GEN_9914; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9916 = 8'hbc == io_state_in_10 ? 8'h48 : _GEN_9915; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9917 = 8'hbd == io_state_in_10 ? 8'h43 : _GEN_9916; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9918 = 8'hbe == io_state_in_10 ? 8'h5e : _GEN_9917; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9919 = 8'hbf == io_state_in_10 ? 8'h55 : _GEN_9918; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9920 = 8'hc0 == io_state_in_10 ? 8'h1 : _GEN_9919; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9921 = 8'hc1 == io_state_in_10 ? 8'ha : _GEN_9920; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9922 = 8'hc2 == io_state_in_10 ? 8'h17 : _GEN_9921; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9923 = 8'hc3 == io_state_in_10 ? 8'h1c : _GEN_9922; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9924 = 8'hc4 == io_state_in_10 ? 8'h2d : _GEN_9923; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9925 = 8'hc5 == io_state_in_10 ? 8'h26 : _GEN_9924; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9926 = 8'hc6 == io_state_in_10 ? 8'h3b : _GEN_9925; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9927 = 8'hc7 == io_state_in_10 ? 8'h30 : _GEN_9926; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9928 = 8'hc8 == io_state_in_10 ? 8'h59 : _GEN_9927; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9929 = 8'hc9 == io_state_in_10 ? 8'h52 : _GEN_9928; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9930 = 8'hca == io_state_in_10 ? 8'h4f : _GEN_9929; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9931 = 8'hcb == io_state_in_10 ? 8'h44 : _GEN_9930; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9932 = 8'hcc == io_state_in_10 ? 8'h75 : _GEN_9931; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9933 = 8'hcd == io_state_in_10 ? 8'h7e : _GEN_9932; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9934 = 8'hce == io_state_in_10 ? 8'h63 : _GEN_9933; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9935 = 8'hcf == io_state_in_10 ? 8'h68 : _GEN_9934; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9936 = 8'hd0 == io_state_in_10 ? 8'hb1 : _GEN_9935; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9937 = 8'hd1 == io_state_in_10 ? 8'hba : _GEN_9936; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9938 = 8'hd2 == io_state_in_10 ? 8'ha7 : _GEN_9937; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9939 = 8'hd3 == io_state_in_10 ? 8'hac : _GEN_9938; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9940 = 8'hd4 == io_state_in_10 ? 8'h9d : _GEN_9939; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9941 = 8'hd5 == io_state_in_10 ? 8'h96 : _GEN_9940; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9942 = 8'hd6 == io_state_in_10 ? 8'h8b : _GEN_9941; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9943 = 8'hd7 == io_state_in_10 ? 8'h80 : _GEN_9942; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9944 = 8'hd8 == io_state_in_10 ? 8'he9 : _GEN_9943; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9945 = 8'hd9 == io_state_in_10 ? 8'he2 : _GEN_9944; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9946 = 8'hda == io_state_in_10 ? 8'hff : _GEN_9945; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9947 = 8'hdb == io_state_in_10 ? 8'hf4 : _GEN_9946; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9948 = 8'hdc == io_state_in_10 ? 8'hc5 : _GEN_9947; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9949 = 8'hdd == io_state_in_10 ? 8'hce : _GEN_9948; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9950 = 8'hde == io_state_in_10 ? 8'hd3 : _GEN_9949; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9951 = 8'hdf == io_state_in_10 ? 8'hd8 : _GEN_9950; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9952 = 8'he0 == io_state_in_10 ? 8'h7a : _GEN_9951; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9953 = 8'he1 == io_state_in_10 ? 8'h71 : _GEN_9952; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9954 = 8'he2 == io_state_in_10 ? 8'h6c : _GEN_9953; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9955 = 8'he3 == io_state_in_10 ? 8'h67 : _GEN_9954; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9956 = 8'he4 == io_state_in_10 ? 8'h56 : _GEN_9955; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9957 = 8'he5 == io_state_in_10 ? 8'h5d : _GEN_9956; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9958 = 8'he6 == io_state_in_10 ? 8'h40 : _GEN_9957; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9959 = 8'he7 == io_state_in_10 ? 8'h4b : _GEN_9958; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9960 = 8'he8 == io_state_in_10 ? 8'h22 : _GEN_9959; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9961 = 8'he9 == io_state_in_10 ? 8'h29 : _GEN_9960; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9962 = 8'hea == io_state_in_10 ? 8'h34 : _GEN_9961; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9963 = 8'heb == io_state_in_10 ? 8'h3f : _GEN_9962; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9964 = 8'hec == io_state_in_10 ? 8'he : _GEN_9963; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9965 = 8'hed == io_state_in_10 ? 8'h5 : _GEN_9964; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9966 = 8'hee == io_state_in_10 ? 8'h18 : _GEN_9965; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9967 = 8'hef == io_state_in_10 ? 8'h13 : _GEN_9966; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9968 = 8'hf0 == io_state_in_10 ? 8'hca : _GEN_9967; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9969 = 8'hf1 == io_state_in_10 ? 8'hc1 : _GEN_9968; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9970 = 8'hf2 == io_state_in_10 ? 8'hdc : _GEN_9969; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9971 = 8'hf3 == io_state_in_10 ? 8'hd7 : _GEN_9970; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9972 = 8'hf4 == io_state_in_10 ? 8'he6 : _GEN_9971; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9973 = 8'hf5 == io_state_in_10 ? 8'hed : _GEN_9972; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9974 = 8'hf6 == io_state_in_10 ? 8'hf0 : _GEN_9973; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9975 = 8'hf7 == io_state_in_10 ? 8'hfb : _GEN_9974; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9976 = 8'hf8 == io_state_in_10 ? 8'h92 : _GEN_9975; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9977 = 8'hf9 == io_state_in_10 ? 8'h99 : _GEN_9976; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9978 = 8'hfa == io_state_in_10 ? 8'h84 : _GEN_9977; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9979 = 8'hfb == io_state_in_10 ? 8'h8f : _GEN_9978; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9980 = 8'hfc == io_state_in_10 ? 8'hbe : _GEN_9979; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9981 = 8'hfd == io_state_in_10 ? 8'hb5 : _GEN_9980; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9982 = 8'hfe == io_state_in_10 ? 8'ha8 : _GEN_9981; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _GEN_9983 = 8'hff == io_state_in_10 ? 8'ha3 : _GEN_9982; // @[InvMixColumns.scala 137:{65,65}]
  wire [7:0] _tmp_state_9_T_1 = _tmp_state_9_T ^ _GEN_9983; // @[InvMixColumns.scala 137:65]
  wire [7:0] _GEN_9985 = 8'h1 == io_state_in_11 ? 8'hd : 8'h0; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9986 = 8'h2 == io_state_in_11 ? 8'h1a : _GEN_9985; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9987 = 8'h3 == io_state_in_11 ? 8'h17 : _GEN_9986; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9988 = 8'h4 == io_state_in_11 ? 8'h34 : _GEN_9987; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9989 = 8'h5 == io_state_in_11 ? 8'h39 : _GEN_9988; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9990 = 8'h6 == io_state_in_11 ? 8'h2e : _GEN_9989; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9991 = 8'h7 == io_state_in_11 ? 8'h23 : _GEN_9990; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9992 = 8'h8 == io_state_in_11 ? 8'h68 : _GEN_9991; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9993 = 8'h9 == io_state_in_11 ? 8'h65 : _GEN_9992; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9994 = 8'ha == io_state_in_11 ? 8'h72 : _GEN_9993; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9995 = 8'hb == io_state_in_11 ? 8'h7f : _GEN_9994; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9996 = 8'hc == io_state_in_11 ? 8'h5c : _GEN_9995; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9997 = 8'hd == io_state_in_11 ? 8'h51 : _GEN_9996; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9998 = 8'he == io_state_in_11 ? 8'h46 : _GEN_9997; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_9999 = 8'hf == io_state_in_11 ? 8'h4b : _GEN_9998; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10000 = 8'h10 == io_state_in_11 ? 8'hd0 : _GEN_9999; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10001 = 8'h11 == io_state_in_11 ? 8'hdd : _GEN_10000; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10002 = 8'h12 == io_state_in_11 ? 8'hca : _GEN_10001; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10003 = 8'h13 == io_state_in_11 ? 8'hc7 : _GEN_10002; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10004 = 8'h14 == io_state_in_11 ? 8'he4 : _GEN_10003; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10005 = 8'h15 == io_state_in_11 ? 8'he9 : _GEN_10004; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10006 = 8'h16 == io_state_in_11 ? 8'hfe : _GEN_10005; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10007 = 8'h17 == io_state_in_11 ? 8'hf3 : _GEN_10006; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10008 = 8'h18 == io_state_in_11 ? 8'hb8 : _GEN_10007; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10009 = 8'h19 == io_state_in_11 ? 8'hb5 : _GEN_10008; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10010 = 8'h1a == io_state_in_11 ? 8'ha2 : _GEN_10009; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10011 = 8'h1b == io_state_in_11 ? 8'haf : _GEN_10010; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10012 = 8'h1c == io_state_in_11 ? 8'h8c : _GEN_10011; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10013 = 8'h1d == io_state_in_11 ? 8'h81 : _GEN_10012; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10014 = 8'h1e == io_state_in_11 ? 8'h96 : _GEN_10013; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10015 = 8'h1f == io_state_in_11 ? 8'h9b : _GEN_10014; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10016 = 8'h20 == io_state_in_11 ? 8'hbb : _GEN_10015; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10017 = 8'h21 == io_state_in_11 ? 8'hb6 : _GEN_10016; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10018 = 8'h22 == io_state_in_11 ? 8'ha1 : _GEN_10017; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10019 = 8'h23 == io_state_in_11 ? 8'hac : _GEN_10018; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10020 = 8'h24 == io_state_in_11 ? 8'h8f : _GEN_10019; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10021 = 8'h25 == io_state_in_11 ? 8'h82 : _GEN_10020; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10022 = 8'h26 == io_state_in_11 ? 8'h95 : _GEN_10021; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10023 = 8'h27 == io_state_in_11 ? 8'h98 : _GEN_10022; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10024 = 8'h28 == io_state_in_11 ? 8'hd3 : _GEN_10023; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10025 = 8'h29 == io_state_in_11 ? 8'hde : _GEN_10024; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10026 = 8'h2a == io_state_in_11 ? 8'hc9 : _GEN_10025; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10027 = 8'h2b == io_state_in_11 ? 8'hc4 : _GEN_10026; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10028 = 8'h2c == io_state_in_11 ? 8'he7 : _GEN_10027; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10029 = 8'h2d == io_state_in_11 ? 8'hea : _GEN_10028; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10030 = 8'h2e == io_state_in_11 ? 8'hfd : _GEN_10029; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10031 = 8'h2f == io_state_in_11 ? 8'hf0 : _GEN_10030; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10032 = 8'h30 == io_state_in_11 ? 8'h6b : _GEN_10031; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10033 = 8'h31 == io_state_in_11 ? 8'h66 : _GEN_10032; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10034 = 8'h32 == io_state_in_11 ? 8'h71 : _GEN_10033; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10035 = 8'h33 == io_state_in_11 ? 8'h7c : _GEN_10034; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10036 = 8'h34 == io_state_in_11 ? 8'h5f : _GEN_10035; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10037 = 8'h35 == io_state_in_11 ? 8'h52 : _GEN_10036; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10038 = 8'h36 == io_state_in_11 ? 8'h45 : _GEN_10037; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10039 = 8'h37 == io_state_in_11 ? 8'h48 : _GEN_10038; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10040 = 8'h38 == io_state_in_11 ? 8'h3 : _GEN_10039; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10041 = 8'h39 == io_state_in_11 ? 8'he : _GEN_10040; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10042 = 8'h3a == io_state_in_11 ? 8'h19 : _GEN_10041; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10043 = 8'h3b == io_state_in_11 ? 8'h14 : _GEN_10042; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10044 = 8'h3c == io_state_in_11 ? 8'h37 : _GEN_10043; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10045 = 8'h3d == io_state_in_11 ? 8'h3a : _GEN_10044; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10046 = 8'h3e == io_state_in_11 ? 8'h2d : _GEN_10045; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10047 = 8'h3f == io_state_in_11 ? 8'h20 : _GEN_10046; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10048 = 8'h40 == io_state_in_11 ? 8'h6d : _GEN_10047; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10049 = 8'h41 == io_state_in_11 ? 8'h60 : _GEN_10048; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10050 = 8'h42 == io_state_in_11 ? 8'h77 : _GEN_10049; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10051 = 8'h43 == io_state_in_11 ? 8'h7a : _GEN_10050; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10052 = 8'h44 == io_state_in_11 ? 8'h59 : _GEN_10051; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10053 = 8'h45 == io_state_in_11 ? 8'h54 : _GEN_10052; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10054 = 8'h46 == io_state_in_11 ? 8'h43 : _GEN_10053; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10055 = 8'h47 == io_state_in_11 ? 8'h4e : _GEN_10054; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10056 = 8'h48 == io_state_in_11 ? 8'h5 : _GEN_10055; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10057 = 8'h49 == io_state_in_11 ? 8'h8 : _GEN_10056; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10058 = 8'h4a == io_state_in_11 ? 8'h1f : _GEN_10057; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10059 = 8'h4b == io_state_in_11 ? 8'h12 : _GEN_10058; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10060 = 8'h4c == io_state_in_11 ? 8'h31 : _GEN_10059; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10061 = 8'h4d == io_state_in_11 ? 8'h3c : _GEN_10060; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10062 = 8'h4e == io_state_in_11 ? 8'h2b : _GEN_10061; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10063 = 8'h4f == io_state_in_11 ? 8'h26 : _GEN_10062; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10064 = 8'h50 == io_state_in_11 ? 8'hbd : _GEN_10063; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10065 = 8'h51 == io_state_in_11 ? 8'hb0 : _GEN_10064; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10066 = 8'h52 == io_state_in_11 ? 8'ha7 : _GEN_10065; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10067 = 8'h53 == io_state_in_11 ? 8'haa : _GEN_10066; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10068 = 8'h54 == io_state_in_11 ? 8'h89 : _GEN_10067; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10069 = 8'h55 == io_state_in_11 ? 8'h84 : _GEN_10068; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10070 = 8'h56 == io_state_in_11 ? 8'h93 : _GEN_10069; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10071 = 8'h57 == io_state_in_11 ? 8'h9e : _GEN_10070; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10072 = 8'h58 == io_state_in_11 ? 8'hd5 : _GEN_10071; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10073 = 8'h59 == io_state_in_11 ? 8'hd8 : _GEN_10072; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10074 = 8'h5a == io_state_in_11 ? 8'hcf : _GEN_10073; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10075 = 8'h5b == io_state_in_11 ? 8'hc2 : _GEN_10074; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10076 = 8'h5c == io_state_in_11 ? 8'he1 : _GEN_10075; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10077 = 8'h5d == io_state_in_11 ? 8'hec : _GEN_10076; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10078 = 8'h5e == io_state_in_11 ? 8'hfb : _GEN_10077; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10079 = 8'h5f == io_state_in_11 ? 8'hf6 : _GEN_10078; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10080 = 8'h60 == io_state_in_11 ? 8'hd6 : _GEN_10079; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10081 = 8'h61 == io_state_in_11 ? 8'hdb : _GEN_10080; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10082 = 8'h62 == io_state_in_11 ? 8'hcc : _GEN_10081; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10083 = 8'h63 == io_state_in_11 ? 8'hc1 : _GEN_10082; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10084 = 8'h64 == io_state_in_11 ? 8'he2 : _GEN_10083; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10085 = 8'h65 == io_state_in_11 ? 8'hef : _GEN_10084; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10086 = 8'h66 == io_state_in_11 ? 8'hf8 : _GEN_10085; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10087 = 8'h67 == io_state_in_11 ? 8'hf5 : _GEN_10086; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10088 = 8'h68 == io_state_in_11 ? 8'hbe : _GEN_10087; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10089 = 8'h69 == io_state_in_11 ? 8'hb3 : _GEN_10088; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10090 = 8'h6a == io_state_in_11 ? 8'ha4 : _GEN_10089; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10091 = 8'h6b == io_state_in_11 ? 8'ha9 : _GEN_10090; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10092 = 8'h6c == io_state_in_11 ? 8'h8a : _GEN_10091; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10093 = 8'h6d == io_state_in_11 ? 8'h87 : _GEN_10092; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10094 = 8'h6e == io_state_in_11 ? 8'h90 : _GEN_10093; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10095 = 8'h6f == io_state_in_11 ? 8'h9d : _GEN_10094; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10096 = 8'h70 == io_state_in_11 ? 8'h6 : _GEN_10095; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10097 = 8'h71 == io_state_in_11 ? 8'hb : _GEN_10096; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10098 = 8'h72 == io_state_in_11 ? 8'h1c : _GEN_10097; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10099 = 8'h73 == io_state_in_11 ? 8'h11 : _GEN_10098; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10100 = 8'h74 == io_state_in_11 ? 8'h32 : _GEN_10099; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10101 = 8'h75 == io_state_in_11 ? 8'h3f : _GEN_10100; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10102 = 8'h76 == io_state_in_11 ? 8'h28 : _GEN_10101; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10103 = 8'h77 == io_state_in_11 ? 8'h25 : _GEN_10102; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10104 = 8'h78 == io_state_in_11 ? 8'h6e : _GEN_10103; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10105 = 8'h79 == io_state_in_11 ? 8'h63 : _GEN_10104; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10106 = 8'h7a == io_state_in_11 ? 8'h74 : _GEN_10105; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10107 = 8'h7b == io_state_in_11 ? 8'h79 : _GEN_10106; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10108 = 8'h7c == io_state_in_11 ? 8'h5a : _GEN_10107; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10109 = 8'h7d == io_state_in_11 ? 8'h57 : _GEN_10108; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10110 = 8'h7e == io_state_in_11 ? 8'h40 : _GEN_10109; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10111 = 8'h7f == io_state_in_11 ? 8'h4d : _GEN_10110; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10112 = 8'h80 == io_state_in_11 ? 8'hda : _GEN_10111; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10113 = 8'h81 == io_state_in_11 ? 8'hd7 : _GEN_10112; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10114 = 8'h82 == io_state_in_11 ? 8'hc0 : _GEN_10113; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10115 = 8'h83 == io_state_in_11 ? 8'hcd : _GEN_10114; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10116 = 8'h84 == io_state_in_11 ? 8'hee : _GEN_10115; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10117 = 8'h85 == io_state_in_11 ? 8'he3 : _GEN_10116; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10118 = 8'h86 == io_state_in_11 ? 8'hf4 : _GEN_10117; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10119 = 8'h87 == io_state_in_11 ? 8'hf9 : _GEN_10118; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10120 = 8'h88 == io_state_in_11 ? 8'hb2 : _GEN_10119; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10121 = 8'h89 == io_state_in_11 ? 8'hbf : _GEN_10120; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10122 = 8'h8a == io_state_in_11 ? 8'ha8 : _GEN_10121; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10123 = 8'h8b == io_state_in_11 ? 8'ha5 : _GEN_10122; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10124 = 8'h8c == io_state_in_11 ? 8'h86 : _GEN_10123; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10125 = 8'h8d == io_state_in_11 ? 8'h8b : _GEN_10124; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10126 = 8'h8e == io_state_in_11 ? 8'h9c : _GEN_10125; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10127 = 8'h8f == io_state_in_11 ? 8'h91 : _GEN_10126; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10128 = 8'h90 == io_state_in_11 ? 8'ha : _GEN_10127; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10129 = 8'h91 == io_state_in_11 ? 8'h7 : _GEN_10128; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10130 = 8'h92 == io_state_in_11 ? 8'h10 : _GEN_10129; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10131 = 8'h93 == io_state_in_11 ? 8'h1d : _GEN_10130; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10132 = 8'h94 == io_state_in_11 ? 8'h3e : _GEN_10131; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10133 = 8'h95 == io_state_in_11 ? 8'h33 : _GEN_10132; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10134 = 8'h96 == io_state_in_11 ? 8'h24 : _GEN_10133; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10135 = 8'h97 == io_state_in_11 ? 8'h29 : _GEN_10134; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10136 = 8'h98 == io_state_in_11 ? 8'h62 : _GEN_10135; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10137 = 8'h99 == io_state_in_11 ? 8'h6f : _GEN_10136; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10138 = 8'h9a == io_state_in_11 ? 8'h78 : _GEN_10137; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10139 = 8'h9b == io_state_in_11 ? 8'h75 : _GEN_10138; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10140 = 8'h9c == io_state_in_11 ? 8'h56 : _GEN_10139; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10141 = 8'h9d == io_state_in_11 ? 8'h5b : _GEN_10140; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10142 = 8'h9e == io_state_in_11 ? 8'h4c : _GEN_10141; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10143 = 8'h9f == io_state_in_11 ? 8'h41 : _GEN_10142; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10144 = 8'ha0 == io_state_in_11 ? 8'h61 : _GEN_10143; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10145 = 8'ha1 == io_state_in_11 ? 8'h6c : _GEN_10144; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10146 = 8'ha2 == io_state_in_11 ? 8'h7b : _GEN_10145; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10147 = 8'ha3 == io_state_in_11 ? 8'h76 : _GEN_10146; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10148 = 8'ha4 == io_state_in_11 ? 8'h55 : _GEN_10147; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10149 = 8'ha5 == io_state_in_11 ? 8'h58 : _GEN_10148; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10150 = 8'ha6 == io_state_in_11 ? 8'h4f : _GEN_10149; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10151 = 8'ha7 == io_state_in_11 ? 8'h42 : _GEN_10150; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10152 = 8'ha8 == io_state_in_11 ? 8'h9 : _GEN_10151; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10153 = 8'ha9 == io_state_in_11 ? 8'h4 : _GEN_10152; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10154 = 8'haa == io_state_in_11 ? 8'h13 : _GEN_10153; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10155 = 8'hab == io_state_in_11 ? 8'h1e : _GEN_10154; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10156 = 8'hac == io_state_in_11 ? 8'h3d : _GEN_10155; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10157 = 8'had == io_state_in_11 ? 8'h30 : _GEN_10156; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10158 = 8'hae == io_state_in_11 ? 8'h27 : _GEN_10157; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10159 = 8'haf == io_state_in_11 ? 8'h2a : _GEN_10158; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10160 = 8'hb0 == io_state_in_11 ? 8'hb1 : _GEN_10159; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10161 = 8'hb1 == io_state_in_11 ? 8'hbc : _GEN_10160; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10162 = 8'hb2 == io_state_in_11 ? 8'hab : _GEN_10161; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10163 = 8'hb3 == io_state_in_11 ? 8'ha6 : _GEN_10162; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10164 = 8'hb4 == io_state_in_11 ? 8'h85 : _GEN_10163; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10165 = 8'hb5 == io_state_in_11 ? 8'h88 : _GEN_10164; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10166 = 8'hb6 == io_state_in_11 ? 8'h9f : _GEN_10165; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10167 = 8'hb7 == io_state_in_11 ? 8'h92 : _GEN_10166; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10168 = 8'hb8 == io_state_in_11 ? 8'hd9 : _GEN_10167; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10169 = 8'hb9 == io_state_in_11 ? 8'hd4 : _GEN_10168; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10170 = 8'hba == io_state_in_11 ? 8'hc3 : _GEN_10169; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10171 = 8'hbb == io_state_in_11 ? 8'hce : _GEN_10170; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10172 = 8'hbc == io_state_in_11 ? 8'hed : _GEN_10171; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10173 = 8'hbd == io_state_in_11 ? 8'he0 : _GEN_10172; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10174 = 8'hbe == io_state_in_11 ? 8'hf7 : _GEN_10173; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10175 = 8'hbf == io_state_in_11 ? 8'hfa : _GEN_10174; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10176 = 8'hc0 == io_state_in_11 ? 8'hb7 : _GEN_10175; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10177 = 8'hc1 == io_state_in_11 ? 8'hba : _GEN_10176; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10178 = 8'hc2 == io_state_in_11 ? 8'had : _GEN_10177; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10179 = 8'hc3 == io_state_in_11 ? 8'ha0 : _GEN_10178; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10180 = 8'hc4 == io_state_in_11 ? 8'h83 : _GEN_10179; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10181 = 8'hc5 == io_state_in_11 ? 8'h8e : _GEN_10180; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10182 = 8'hc6 == io_state_in_11 ? 8'h99 : _GEN_10181; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10183 = 8'hc7 == io_state_in_11 ? 8'h94 : _GEN_10182; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10184 = 8'hc8 == io_state_in_11 ? 8'hdf : _GEN_10183; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10185 = 8'hc9 == io_state_in_11 ? 8'hd2 : _GEN_10184; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10186 = 8'hca == io_state_in_11 ? 8'hc5 : _GEN_10185; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10187 = 8'hcb == io_state_in_11 ? 8'hc8 : _GEN_10186; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10188 = 8'hcc == io_state_in_11 ? 8'heb : _GEN_10187; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10189 = 8'hcd == io_state_in_11 ? 8'he6 : _GEN_10188; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10190 = 8'hce == io_state_in_11 ? 8'hf1 : _GEN_10189; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10191 = 8'hcf == io_state_in_11 ? 8'hfc : _GEN_10190; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10192 = 8'hd0 == io_state_in_11 ? 8'h67 : _GEN_10191; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10193 = 8'hd1 == io_state_in_11 ? 8'h6a : _GEN_10192; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10194 = 8'hd2 == io_state_in_11 ? 8'h7d : _GEN_10193; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10195 = 8'hd3 == io_state_in_11 ? 8'h70 : _GEN_10194; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10196 = 8'hd4 == io_state_in_11 ? 8'h53 : _GEN_10195; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10197 = 8'hd5 == io_state_in_11 ? 8'h5e : _GEN_10196; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10198 = 8'hd6 == io_state_in_11 ? 8'h49 : _GEN_10197; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10199 = 8'hd7 == io_state_in_11 ? 8'h44 : _GEN_10198; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10200 = 8'hd8 == io_state_in_11 ? 8'hf : _GEN_10199; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10201 = 8'hd9 == io_state_in_11 ? 8'h2 : _GEN_10200; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10202 = 8'hda == io_state_in_11 ? 8'h15 : _GEN_10201; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10203 = 8'hdb == io_state_in_11 ? 8'h18 : _GEN_10202; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10204 = 8'hdc == io_state_in_11 ? 8'h3b : _GEN_10203; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10205 = 8'hdd == io_state_in_11 ? 8'h36 : _GEN_10204; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10206 = 8'hde == io_state_in_11 ? 8'h21 : _GEN_10205; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10207 = 8'hdf == io_state_in_11 ? 8'h2c : _GEN_10206; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10208 = 8'he0 == io_state_in_11 ? 8'hc : _GEN_10207; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10209 = 8'he1 == io_state_in_11 ? 8'h1 : _GEN_10208; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10210 = 8'he2 == io_state_in_11 ? 8'h16 : _GEN_10209; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10211 = 8'he3 == io_state_in_11 ? 8'h1b : _GEN_10210; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10212 = 8'he4 == io_state_in_11 ? 8'h38 : _GEN_10211; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10213 = 8'he5 == io_state_in_11 ? 8'h35 : _GEN_10212; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10214 = 8'he6 == io_state_in_11 ? 8'h22 : _GEN_10213; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10215 = 8'he7 == io_state_in_11 ? 8'h2f : _GEN_10214; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10216 = 8'he8 == io_state_in_11 ? 8'h64 : _GEN_10215; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10217 = 8'he9 == io_state_in_11 ? 8'h69 : _GEN_10216; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10218 = 8'hea == io_state_in_11 ? 8'h7e : _GEN_10217; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10219 = 8'heb == io_state_in_11 ? 8'h73 : _GEN_10218; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10220 = 8'hec == io_state_in_11 ? 8'h50 : _GEN_10219; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10221 = 8'hed == io_state_in_11 ? 8'h5d : _GEN_10220; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10222 = 8'hee == io_state_in_11 ? 8'h4a : _GEN_10221; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10223 = 8'hef == io_state_in_11 ? 8'h47 : _GEN_10222; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10224 = 8'hf0 == io_state_in_11 ? 8'hdc : _GEN_10223; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10225 = 8'hf1 == io_state_in_11 ? 8'hd1 : _GEN_10224; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10226 = 8'hf2 == io_state_in_11 ? 8'hc6 : _GEN_10225; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10227 = 8'hf3 == io_state_in_11 ? 8'hcb : _GEN_10226; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10228 = 8'hf4 == io_state_in_11 ? 8'he8 : _GEN_10227; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10229 = 8'hf5 == io_state_in_11 ? 8'he5 : _GEN_10228; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10230 = 8'hf6 == io_state_in_11 ? 8'hf2 : _GEN_10229; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10231 = 8'hf7 == io_state_in_11 ? 8'hff : _GEN_10230; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10232 = 8'hf8 == io_state_in_11 ? 8'hb4 : _GEN_10231; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10233 = 8'hf9 == io_state_in_11 ? 8'hb9 : _GEN_10232; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10234 = 8'hfa == io_state_in_11 ? 8'hae : _GEN_10233; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10235 = 8'hfb == io_state_in_11 ? 8'ha3 : _GEN_10234; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10236 = 8'hfc == io_state_in_11 ? 8'h80 : _GEN_10235; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10237 = 8'hfd == io_state_in_11 ? 8'h8d : _GEN_10236; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10238 = 8'hfe == io_state_in_11 ? 8'h9a : _GEN_10237; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10239 = 8'hff == io_state_in_11 ? 8'h97 : _GEN_10238; // @[InvMixColumns.scala 137:{90,90}]
  wire [7:0] _GEN_10241 = 8'h1 == io_state_in_8 ? 8'hd : 8'h0; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10242 = 8'h2 == io_state_in_8 ? 8'h1a : _GEN_10241; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10243 = 8'h3 == io_state_in_8 ? 8'h17 : _GEN_10242; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10244 = 8'h4 == io_state_in_8 ? 8'h34 : _GEN_10243; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10245 = 8'h5 == io_state_in_8 ? 8'h39 : _GEN_10244; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10246 = 8'h6 == io_state_in_8 ? 8'h2e : _GEN_10245; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10247 = 8'h7 == io_state_in_8 ? 8'h23 : _GEN_10246; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10248 = 8'h8 == io_state_in_8 ? 8'h68 : _GEN_10247; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10249 = 8'h9 == io_state_in_8 ? 8'h65 : _GEN_10248; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10250 = 8'ha == io_state_in_8 ? 8'h72 : _GEN_10249; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10251 = 8'hb == io_state_in_8 ? 8'h7f : _GEN_10250; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10252 = 8'hc == io_state_in_8 ? 8'h5c : _GEN_10251; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10253 = 8'hd == io_state_in_8 ? 8'h51 : _GEN_10252; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10254 = 8'he == io_state_in_8 ? 8'h46 : _GEN_10253; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10255 = 8'hf == io_state_in_8 ? 8'h4b : _GEN_10254; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10256 = 8'h10 == io_state_in_8 ? 8'hd0 : _GEN_10255; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10257 = 8'h11 == io_state_in_8 ? 8'hdd : _GEN_10256; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10258 = 8'h12 == io_state_in_8 ? 8'hca : _GEN_10257; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10259 = 8'h13 == io_state_in_8 ? 8'hc7 : _GEN_10258; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10260 = 8'h14 == io_state_in_8 ? 8'he4 : _GEN_10259; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10261 = 8'h15 == io_state_in_8 ? 8'he9 : _GEN_10260; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10262 = 8'h16 == io_state_in_8 ? 8'hfe : _GEN_10261; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10263 = 8'h17 == io_state_in_8 ? 8'hf3 : _GEN_10262; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10264 = 8'h18 == io_state_in_8 ? 8'hb8 : _GEN_10263; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10265 = 8'h19 == io_state_in_8 ? 8'hb5 : _GEN_10264; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10266 = 8'h1a == io_state_in_8 ? 8'ha2 : _GEN_10265; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10267 = 8'h1b == io_state_in_8 ? 8'haf : _GEN_10266; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10268 = 8'h1c == io_state_in_8 ? 8'h8c : _GEN_10267; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10269 = 8'h1d == io_state_in_8 ? 8'h81 : _GEN_10268; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10270 = 8'h1e == io_state_in_8 ? 8'h96 : _GEN_10269; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10271 = 8'h1f == io_state_in_8 ? 8'h9b : _GEN_10270; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10272 = 8'h20 == io_state_in_8 ? 8'hbb : _GEN_10271; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10273 = 8'h21 == io_state_in_8 ? 8'hb6 : _GEN_10272; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10274 = 8'h22 == io_state_in_8 ? 8'ha1 : _GEN_10273; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10275 = 8'h23 == io_state_in_8 ? 8'hac : _GEN_10274; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10276 = 8'h24 == io_state_in_8 ? 8'h8f : _GEN_10275; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10277 = 8'h25 == io_state_in_8 ? 8'h82 : _GEN_10276; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10278 = 8'h26 == io_state_in_8 ? 8'h95 : _GEN_10277; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10279 = 8'h27 == io_state_in_8 ? 8'h98 : _GEN_10278; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10280 = 8'h28 == io_state_in_8 ? 8'hd3 : _GEN_10279; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10281 = 8'h29 == io_state_in_8 ? 8'hde : _GEN_10280; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10282 = 8'h2a == io_state_in_8 ? 8'hc9 : _GEN_10281; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10283 = 8'h2b == io_state_in_8 ? 8'hc4 : _GEN_10282; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10284 = 8'h2c == io_state_in_8 ? 8'he7 : _GEN_10283; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10285 = 8'h2d == io_state_in_8 ? 8'hea : _GEN_10284; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10286 = 8'h2e == io_state_in_8 ? 8'hfd : _GEN_10285; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10287 = 8'h2f == io_state_in_8 ? 8'hf0 : _GEN_10286; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10288 = 8'h30 == io_state_in_8 ? 8'h6b : _GEN_10287; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10289 = 8'h31 == io_state_in_8 ? 8'h66 : _GEN_10288; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10290 = 8'h32 == io_state_in_8 ? 8'h71 : _GEN_10289; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10291 = 8'h33 == io_state_in_8 ? 8'h7c : _GEN_10290; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10292 = 8'h34 == io_state_in_8 ? 8'h5f : _GEN_10291; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10293 = 8'h35 == io_state_in_8 ? 8'h52 : _GEN_10292; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10294 = 8'h36 == io_state_in_8 ? 8'h45 : _GEN_10293; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10295 = 8'h37 == io_state_in_8 ? 8'h48 : _GEN_10294; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10296 = 8'h38 == io_state_in_8 ? 8'h3 : _GEN_10295; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10297 = 8'h39 == io_state_in_8 ? 8'he : _GEN_10296; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10298 = 8'h3a == io_state_in_8 ? 8'h19 : _GEN_10297; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10299 = 8'h3b == io_state_in_8 ? 8'h14 : _GEN_10298; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10300 = 8'h3c == io_state_in_8 ? 8'h37 : _GEN_10299; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10301 = 8'h3d == io_state_in_8 ? 8'h3a : _GEN_10300; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10302 = 8'h3e == io_state_in_8 ? 8'h2d : _GEN_10301; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10303 = 8'h3f == io_state_in_8 ? 8'h20 : _GEN_10302; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10304 = 8'h40 == io_state_in_8 ? 8'h6d : _GEN_10303; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10305 = 8'h41 == io_state_in_8 ? 8'h60 : _GEN_10304; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10306 = 8'h42 == io_state_in_8 ? 8'h77 : _GEN_10305; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10307 = 8'h43 == io_state_in_8 ? 8'h7a : _GEN_10306; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10308 = 8'h44 == io_state_in_8 ? 8'h59 : _GEN_10307; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10309 = 8'h45 == io_state_in_8 ? 8'h54 : _GEN_10308; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10310 = 8'h46 == io_state_in_8 ? 8'h43 : _GEN_10309; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10311 = 8'h47 == io_state_in_8 ? 8'h4e : _GEN_10310; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10312 = 8'h48 == io_state_in_8 ? 8'h5 : _GEN_10311; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10313 = 8'h49 == io_state_in_8 ? 8'h8 : _GEN_10312; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10314 = 8'h4a == io_state_in_8 ? 8'h1f : _GEN_10313; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10315 = 8'h4b == io_state_in_8 ? 8'h12 : _GEN_10314; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10316 = 8'h4c == io_state_in_8 ? 8'h31 : _GEN_10315; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10317 = 8'h4d == io_state_in_8 ? 8'h3c : _GEN_10316; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10318 = 8'h4e == io_state_in_8 ? 8'h2b : _GEN_10317; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10319 = 8'h4f == io_state_in_8 ? 8'h26 : _GEN_10318; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10320 = 8'h50 == io_state_in_8 ? 8'hbd : _GEN_10319; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10321 = 8'h51 == io_state_in_8 ? 8'hb0 : _GEN_10320; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10322 = 8'h52 == io_state_in_8 ? 8'ha7 : _GEN_10321; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10323 = 8'h53 == io_state_in_8 ? 8'haa : _GEN_10322; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10324 = 8'h54 == io_state_in_8 ? 8'h89 : _GEN_10323; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10325 = 8'h55 == io_state_in_8 ? 8'h84 : _GEN_10324; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10326 = 8'h56 == io_state_in_8 ? 8'h93 : _GEN_10325; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10327 = 8'h57 == io_state_in_8 ? 8'h9e : _GEN_10326; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10328 = 8'h58 == io_state_in_8 ? 8'hd5 : _GEN_10327; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10329 = 8'h59 == io_state_in_8 ? 8'hd8 : _GEN_10328; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10330 = 8'h5a == io_state_in_8 ? 8'hcf : _GEN_10329; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10331 = 8'h5b == io_state_in_8 ? 8'hc2 : _GEN_10330; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10332 = 8'h5c == io_state_in_8 ? 8'he1 : _GEN_10331; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10333 = 8'h5d == io_state_in_8 ? 8'hec : _GEN_10332; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10334 = 8'h5e == io_state_in_8 ? 8'hfb : _GEN_10333; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10335 = 8'h5f == io_state_in_8 ? 8'hf6 : _GEN_10334; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10336 = 8'h60 == io_state_in_8 ? 8'hd6 : _GEN_10335; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10337 = 8'h61 == io_state_in_8 ? 8'hdb : _GEN_10336; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10338 = 8'h62 == io_state_in_8 ? 8'hcc : _GEN_10337; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10339 = 8'h63 == io_state_in_8 ? 8'hc1 : _GEN_10338; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10340 = 8'h64 == io_state_in_8 ? 8'he2 : _GEN_10339; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10341 = 8'h65 == io_state_in_8 ? 8'hef : _GEN_10340; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10342 = 8'h66 == io_state_in_8 ? 8'hf8 : _GEN_10341; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10343 = 8'h67 == io_state_in_8 ? 8'hf5 : _GEN_10342; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10344 = 8'h68 == io_state_in_8 ? 8'hbe : _GEN_10343; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10345 = 8'h69 == io_state_in_8 ? 8'hb3 : _GEN_10344; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10346 = 8'h6a == io_state_in_8 ? 8'ha4 : _GEN_10345; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10347 = 8'h6b == io_state_in_8 ? 8'ha9 : _GEN_10346; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10348 = 8'h6c == io_state_in_8 ? 8'h8a : _GEN_10347; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10349 = 8'h6d == io_state_in_8 ? 8'h87 : _GEN_10348; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10350 = 8'h6e == io_state_in_8 ? 8'h90 : _GEN_10349; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10351 = 8'h6f == io_state_in_8 ? 8'h9d : _GEN_10350; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10352 = 8'h70 == io_state_in_8 ? 8'h6 : _GEN_10351; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10353 = 8'h71 == io_state_in_8 ? 8'hb : _GEN_10352; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10354 = 8'h72 == io_state_in_8 ? 8'h1c : _GEN_10353; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10355 = 8'h73 == io_state_in_8 ? 8'h11 : _GEN_10354; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10356 = 8'h74 == io_state_in_8 ? 8'h32 : _GEN_10355; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10357 = 8'h75 == io_state_in_8 ? 8'h3f : _GEN_10356; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10358 = 8'h76 == io_state_in_8 ? 8'h28 : _GEN_10357; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10359 = 8'h77 == io_state_in_8 ? 8'h25 : _GEN_10358; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10360 = 8'h78 == io_state_in_8 ? 8'h6e : _GEN_10359; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10361 = 8'h79 == io_state_in_8 ? 8'h63 : _GEN_10360; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10362 = 8'h7a == io_state_in_8 ? 8'h74 : _GEN_10361; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10363 = 8'h7b == io_state_in_8 ? 8'h79 : _GEN_10362; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10364 = 8'h7c == io_state_in_8 ? 8'h5a : _GEN_10363; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10365 = 8'h7d == io_state_in_8 ? 8'h57 : _GEN_10364; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10366 = 8'h7e == io_state_in_8 ? 8'h40 : _GEN_10365; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10367 = 8'h7f == io_state_in_8 ? 8'h4d : _GEN_10366; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10368 = 8'h80 == io_state_in_8 ? 8'hda : _GEN_10367; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10369 = 8'h81 == io_state_in_8 ? 8'hd7 : _GEN_10368; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10370 = 8'h82 == io_state_in_8 ? 8'hc0 : _GEN_10369; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10371 = 8'h83 == io_state_in_8 ? 8'hcd : _GEN_10370; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10372 = 8'h84 == io_state_in_8 ? 8'hee : _GEN_10371; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10373 = 8'h85 == io_state_in_8 ? 8'he3 : _GEN_10372; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10374 = 8'h86 == io_state_in_8 ? 8'hf4 : _GEN_10373; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10375 = 8'h87 == io_state_in_8 ? 8'hf9 : _GEN_10374; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10376 = 8'h88 == io_state_in_8 ? 8'hb2 : _GEN_10375; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10377 = 8'h89 == io_state_in_8 ? 8'hbf : _GEN_10376; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10378 = 8'h8a == io_state_in_8 ? 8'ha8 : _GEN_10377; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10379 = 8'h8b == io_state_in_8 ? 8'ha5 : _GEN_10378; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10380 = 8'h8c == io_state_in_8 ? 8'h86 : _GEN_10379; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10381 = 8'h8d == io_state_in_8 ? 8'h8b : _GEN_10380; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10382 = 8'h8e == io_state_in_8 ? 8'h9c : _GEN_10381; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10383 = 8'h8f == io_state_in_8 ? 8'h91 : _GEN_10382; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10384 = 8'h90 == io_state_in_8 ? 8'ha : _GEN_10383; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10385 = 8'h91 == io_state_in_8 ? 8'h7 : _GEN_10384; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10386 = 8'h92 == io_state_in_8 ? 8'h10 : _GEN_10385; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10387 = 8'h93 == io_state_in_8 ? 8'h1d : _GEN_10386; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10388 = 8'h94 == io_state_in_8 ? 8'h3e : _GEN_10387; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10389 = 8'h95 == io_state_in_8 ? 8'h33 : _GEN_10388; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10390 = 8'h96 == io_state_in_8 ? 8'h24 : _GEN_10389; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10391 = 8'h97 == io_state_in_8 ? 8'h29 : _GEN_10390; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10392 = 8'h98 == io_state_in_8 ? 8'h62 : _GEN_10391; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10393 = 8'h99 == io_state_in_8 ? 8'h6f : _GEN_10392; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10394 = 8'h9a == io_state_in_8 ? 8'h78 : _GEN_10393; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10395 = 8'h9b == io_state_in_8 ? 8'h75 : _GEN_10394; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10396 = 8'h9c == io_state_in_8 ? 8'h56 : _GEN_10395; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10397 = 8'h9d == io_state_in_8 ? 8'h5b : _GEN_10396; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10398 = 8'h9e == io_state_in_8 ? 8'h4c : _GEN_10397; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10399 = 8'h9f == io_state_in_8 ? 8'h41 : _GEN_10398; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10400 = 8'ha0 == io_state_in_8 ? 8'h61 : _GEN_10399; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10401 = 8'ha1 == io_state_in_8 ? 8'h6c : _GEN_10400; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10402 = 8'ha2 == io_state_in_8 ? 8'h7b : _GEN_10401; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10403 = 8'ha3 == io_state_in_8 ? 8'h76 : _GEN_10402; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10404 = 8'ha4 == io_state_in_8 ? 8'h55 : _GEN_10403; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10405 = 8'ha5 == io_state_in_8 ? 8'h58 : _GEN_10404; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10406 = 8'ha6 == io_state_in_8 ? 8'h4f : _GEN_10405; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10407 = 8'ha7 == io_state_in_8 ? 8'h42 : _GEN_10406; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10408 = 8'ha8 == io_state_in_8 ? 8'h9 : _GEN_10407; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10409 = 8'ha9 == io_state_in_8 ? 8'h4 : _GEN_10408; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10410 = 8'haa == io_state_in_8 ? 8'h13 : _GEN_10409; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10411 = 8'hab == io_state_in_8 ? 8'h1e : _GEN_10410; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10412 = 8'hac == io_state_in_8 ? 8'h3d : _GEN_10411; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10413 = 8'had == io_state_in_8 ? 8'h30 : _GEN_10412; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10414 = 8'hae == io_state_in_8 ? 8'h27 : _GEN_10413; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10415 = 8'haf == io_state_in_8 ? 8'h2a : _GEN_10414; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10416 = 8'hb0 == io_state_in_8 ? 8'hb1 : _GEN_10415; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10417 = 8'hb1 == io_state_in_8 ? 8'hbc : _GEN_10416; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10418 = 8'hb2 == io_state_in_8 ? 8'hab : _GEN_10417; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10419 = 8'hb3 == io_state_in_8 ? 8'ha6 : _GEN_10418; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10420 = 8'hb4 == io_state_in_8 ? 8'h85 : _GEN_10419; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10421 = 8'hb5 == io_state_in_8 ? 8'h88 : _GEN_10420; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10422 = 8'hb6 == io_state_in_8 ? 8'h9f : _GEN_10421; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10423 = 8'hb7 == io_state_in_8 ? 8'h92 : _GEN_10422; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10424 = 8'hb8 == io_state_in_8 ? 8'hd9 : _GEN_10423; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10425 = 8'hb9 == io_state_in_8 ? 8'hd4 : _GEN_10424; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10426 = 8'hba == io_state_in_8 ? 8'hc3 : _GEN_10425; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10427 = 8'hbb == io_state_in_8 ? 8'hce : _GEN_10426; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10428 = 8'hbc == io_state_in_8 ? 8'hed : _GEN_10427; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10429 = 8'hbd == io_state_in_8 ? 8'he0 : _GEN_10428; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10430 = 8'hbe == io_state_in_8 ? 8'hf7 : _GEN_10429; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10431 = 8'hbf == io_state_in_8 ? 8'hfa : _GEN_10430; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10432 = 8'hc0 == io_state_in_8 ? 8'hb7 : _GEN_10431; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10433 = 8'hc1 == io_state_in_8 ? 8'hba : _GEN_10432; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10434 = 8'hc2 == io_state_in_8 ? 8'had : _GEN_10433; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10435 = 8'hc3 == io_state_in_8 ? 8'ha0 : _GEN_10434; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10436 = 8'hc4 == io_state_in_8 ? 8'h83 : _GEN_10435; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10437 = 8'hc5 == io_state_in_8 ? 8'h8e : _GEN_10436; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10438 = 8'hc6 == io_state_in_8 ? 8'h99 : _GEN_10437; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10439 = 8'hc7 == io_state_in_8 ? 8'h94 : _GEN_10438; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10440 = 8'hc8 == io_state_in_8 ? 8'hdf : _GEN_10439; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10441 = 8'hc9 == io_state_in_8 ? 8'hd2 : _GEN_10440; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10442 = 8'hca == io_state_in_8 ? 8'hc5 : _GEN_10441; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10443 = 8'hcb == io_state_in_8 ? 8'hc8 : _GEN_10442; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10444 = 8'hcc == io_state_in_8 ? 8'heb : _GEN_10443; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10445 = 8'hcd == io_state_in_8 ? 8'he6 : _GEN_10444; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10446 = 8'hce == io_state_in_8 ? 8'hf1 : _GEN_10445; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10447 = 8'hcf == io_state_in_8 ? 8'hfc : _GEN_10446; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10448 = 8'hd0 == io_state_in_8 ? 8'h67 : _GEN_10447; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10449 = 8'hd1 == io_state_in_8 ? 8'h6a : _GEN_10448; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10450 = 8'hd2 == io_state_in_8 ? 8'h7d : _GEN_10449; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10451 = 8'hd3 == io_state_in_8 ? 8'h70 : _GEN_10450; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10452 = 8'hd4 == io_state_in_8 ? 8'h53 : _GEN_10451; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10453 = 8'hd5 == io_state_in_8 ? 8'h5e : _GEN_10452; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10454 = 8'hd6 == io_state_in_8 ? 8'h49 : _GEN_10453; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10455 = 8'hd7 == io_state_in_8 ? 8'h44 : _GEN_10454; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10456 = 8'hd8 == io_state_in_8 ? 8'hf : _GEN_10455; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10457 = 8'hd9 == io_state_in_8 ? 8'h2 : _GEN_10456; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10458 = 8'hda == io_state_in_8 ? 8'h15 : _GEN_10457; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10459 = 8'hdb == io_state_in_8 ? 8'h18 : _GEN_10458; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10460 = 8'hdc == io_state_in_8 ? 8'h3b : _GEN_10459; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10461 = 8'hdd == io_state_in_8 ? 8'h36 : _GEN_10460; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10462 = 8'hde == io_state_in_8 ? 8'h21 : _GEN_10461; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10463 = 8'hdf == io_state_in_8 ? 8'h2c : _GEN_10462; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10464 = 8'he0 == io_state_in_8 ? 8'hc : _GEN_10463; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10465 = 8'he1 == io_state_in_8 ? 8'h1 : _GEN_10464; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10466 = 8'he2 == io_state_in_8 ? 8'h16 : _GEN_10465; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10467 = 8'he3 == io_state_in_8 ? 8'h1b : _GEN_10466; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10468 = 8'he4 == io_state_in_8 ? 8'h38 : _GEN_10467; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10469 = 8'he5 == io_state_in_8 ? 8'h35 : _GEN_10468; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10470 = 8'he6 == io_state_in_8 ? 8'h22 : _GEN_10469; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10471 = 8'he7 == io_state_in_8 ? 8'h2f : _GEN_10470; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10472 = 8'he8 == io_state_in_8 ? 8'h64 : _GEN_10471; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10473 = 8'he9 == io_state_in_8 ? 8'h69 : _GEN_10472; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10474 = 8'hea == io_state_in_8 ? 8'h7e : _GEN_10473; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10475 = 8'heb == io_state_in_8 ? 8'h73 : _GEN_10474; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10476 = 8'hec == io_state_in_8 ? 8'h50 : _GEN_10475; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10477 = 8'hed == io_state_in_8 ? 8'h5d : _GEN_10476; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10478 = 8'hee == io_state_in_8 ? 8'h4a : _GEN_10477; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10479 = 8'hef == io_state_in_8 ? 8'h47 : _GEN_10478; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10480 = 8'hf0 == io_state_in_8 ? 8'hdc : _GEN_10479; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10481 = 8'hf1 == io_state_in_8 ? 8'hd1 : _GEN_10480; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10482 = 8'hf2 == io_state_in_8 ? 8'hc6 : _GEN_10481; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10483 = 8'hf3 == io_state_in_8 ? 8'hcb : _GEN_10482; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10484 = 8'hf4 == io_state_in_8 ? 8'he8 : _GEN_10483; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10485 = 8'hf5 == io_state_in_8 ? 8'he5 : _GEN_10484; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10486 = 8'hf6 == io_state_in_8 ? 8'hf2 : _GEN_10485; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10487 = 8'hf7 == io_state_in_8 ? 8'hff : _GEN_10486; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10488 = 8'hf8 == io_state_in_8 ? 8'hb4 : _GEN_10487; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10489 = 8'hf9 == io_state_in_8 ? 8'hb9 : _GEN_10488; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10490 = 8'hfa == io_state_in_8 ? 8'hae : _GEN_10489; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10491 = 8'hfb == io_state_in_8 ? 8'ha3 : _GEN_10490; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10492 = 8'hfc == io_state_in_8 ? 8'h80 : _GEN_10491; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10493 = 8'hfd == io_state_in_8 ? 8'h8d : _GEN_10492; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10494 = 8'hfe == io_state_in_8 ? 8'h9a : _GEN_10493; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10495 = 8'hff == io_state_in_8 ? 8'h97 : _GEN_10494; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10497 = 8'h1 == io_state_in_9 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10498 = 8'h2 == io_state_in_9 ? 8'h12 : _GEN_10497; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10499 = 8'h3 == io_state_in_9 ? 8'h1b : _GEN_10498; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10500 = 8'h4 == io_state_in_9 ? 8'h24 : _GEN_10499; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10501 = 8'h5 == io_state_in_9 ? 8'h2d : _GEN_10500; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10502 = 8'h6 == io_state_in_9 ? 8'h36 : _GEN_10501; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10503 = 8'h7 == io_state_in_9 ? 8'h3f : _GEN_10502; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10504 = 8'h8 == io_state_in_9 ? 8'h48 : _GEN_10503; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10505 = 8'h9 == io_state_in_9 ? 8'h41 : _GEN_10504; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10506 = 8'ha == io_state_in_9 ? 8'h5a : _GEN_10505; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10507 = 8'hb == io_state_in_9 ? 8'h53 : _GEN_10506; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10508 = 8'hc == io_state_in_9 ? 8'h6c : _GEN_10507; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10509 = 8'hd == io_state_in_9 ? 8'h65 : _GEN_10508; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10510 = 8'he == io_state_in_9 ? 8'h7e : _GEN_10509; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10511 = 8'hf == io_state_in_9 ? 8'h77 : _GEN_10510; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10512 = 8'h10 == io_state_in_9 ? 8'h90 : _GEN_10511; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10513 = 8'h11 == io_state_in_9 ? 8'h99 : _GEN_10512; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10514 = 8'h12 == io_state_in_9 ? 8'h82 : _GEN_10513; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10515 = 8'h13 == io_state_in_9 ? 8'h8b : _GEN_10514; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10516 = 8'h14 == io_state_in_9 ? 8'hb4 : _GEN_10515; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10517 = 8'h15 == io_state_in_9 ? 8'hbd : _GEN_10516; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10518 = 8'h16 == io_state_in_9 ? 8'ha6 : _GEN_10517; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10519 = 8'h17 == io_state_in_9 ? 8'haf : _GEN_10518; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10520 = 8'h18 == io_state_in_9 ? 8'hd8 : _GEN_10519; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10521 = 8'h19 == io_state_in_9 ? 8'hd1 : _GEN_10520; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10522 = 8'h1a == io_state_in_9 ? 8'hca : _GEN_10521; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10523 = 8'h1b == io_state_in_9 ? 8'hc3 : _GEN_10522; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10524 = 8'h1c == io_state_in_9 ? 8'hfc : _GEN_10523; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10525 = 8'h1d == io_state_in_9 ? 8'hf5 : _GEN_10524; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10526 = 8'h1e == io_state_in_9 ? 8'hee : _GEN_10525; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10527 = 8'h1f == io_state_in_9 ? 8'he7 : _GEN_10526; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10528 = 8'h20 == io_state_in_9 ? 8'h3b : _GEN_10527; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10529 = 8'h21 == io_state_in_9 ? 8'h32 : _GEN_10528; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10530 = 8'h22 == io_state_in_9 ? 8'h29 : _GEN_10529; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10531 = 8'h23 == io_state_in_9 ? 8'h20 : _GEN_10530; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10532 = 8'h24 == io_state_in_9 ? 8'h1f : _GEN_10531; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10533 = 8'h25 == io_state_in_9 ? 8'h16 : _GEN_10532; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10534 = 8'h26 == io_state_in_9 ? 8'hd : _GEN_10533; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10535 = 8'h27 == io_state_in_9 ? 8'h4 : _GEN_10534; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10536 = 8'h28 == io_state_in_9 ? 8'h73 : _GEN_10535; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10537 = 8'h29 == io_state_in_9 ? 8'h7a : _GEN_10536; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10538 = 8'h2a == io_state_in_9 ? 8'h61 : _GEN_10537; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10539 = 8'h2b == io_state_in_9 ? 8'h68 : _GEN_10538; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10540 = 8'h2c == io_state_in_9 ? 8'h57 : _GEN_10539; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10541 = 8'h2d == io_state_in_9 ? 8'h5e : _GEN_10540; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10542 = 8'h2e == io_state_in_9 ? 8'h45 : _GEN_10541; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10543 = 8'h2f == io_state_in_9 ? 8'h4c : _GEN_10542; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10544 = 8'h30 == io_state_in_9 ? 8'hab : _GEN_10543; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10545 = 8'h31 == io_state_in_9 ? 8'ha2 : _GEN_10544; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10546 = 8'h32 == io_state_in_9 ? 8'hb9 : _GEN_10545; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10547 = 8'h33 == io_state_in_9 ? 8'hb0 : _GEN_10546; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10548 = 8'h34 == io_state_in_9 ? 8'h8f : _GEN_10547; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10549 = 8'h35 == io_state_in_9 ? 8'h86 : _GEN_10548; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10550 = 8'h36 == io_state_in_9 ? 8'h9d : _GEN_10549; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10551 = 8'h37 == io_state_in_9 ? 8'h94 : _GEN_10550; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10552 = 8'h38 == io_state_in_9 ? 8'he3 : _GEN_10551; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10553 = 8'h39 == io_state_in_9 ? 8'hea : _GEN_10552; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10554 = 8'h3a == io_state_in_9 ? 8'hf1 : _GEN_10553; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10555 = 8'h3b == io_state_in_9 ? 8'hf8 : _GEN_10554; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10556 = 8'h3c == io_state_in_9 ? 8'hc7 : _GEN_10555; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10557 = 8'h3d == io_state_in_9 ? 8'hce : _GEN_10556; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10558 = 8'h3e == io_state_in_9 ? 8'hd5 : _GEN_10557; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10559 = 8'h3f == io_state_in_9 ? 8'hdc : _GEN_10558; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10560 = 8'h40 == io_state_in_9 ? 8'h76 : _GEN_10559; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10561 = 8'h41 == io_state_in_9 ? 8'h7f : _GEN_10560; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10562 = 8'h42 == io_state_in_9 ? 8'h64 : _GEN_10561; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10563 = 8'h43 == io_state_in_9 ? 8'h6d : _GEN_10562; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10564 = 8'h44 == io_state_in_9 ? 8'h52 : _GEN_10563; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10565 = 8'h45 == io_state_in_9 ? 8'h5b : _GEN_10564; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10566 = 8'h46 == io_state_in_9 ? 8'h40 : _GEN_10565; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10567 = 8'h47 == io_state_in_9 ? 8'h49 : _GEN_10566; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10568 = 8'h48 == io_state_in_9 ? 8'h3e : _GEN_10567; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10569 = 8'h49 == io_state_in_9 ? 8'h37 : _GEN_10568; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10570 = 8'h4a == io_state_in_9 ? 8'h2c : _GEN_10569; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10571 = 8'h4b == io_state_in_9 ? 8'h25 : _GEN_10570; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10572 = 8'h4c == io_state_in_9 ? 8'h1a : _GEN_10571; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10573 = 8'h4d == io_state_in_9 ? 8'h13 : _GEN_10572; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10574 = 8'h4e == io_state_in_9 ? 8'h8 : _GEN_10573; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10575 = 8'h4f == io_state_in_9 ? 8'h1 : _GEN_10574; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10576 = 8'h50 == io_state_in_9 ? 8'he6 : _GEN_10575; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10577 = 8'h51 == io_state_in_9 ? 8'hef : _GEN_10576; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10578 = 8'h52 == io_state_in_9 ? 8'hf4 : _GEN_10577; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10579 = 8'h53 == io_state_in_9 ? 8'hfd : _GEN_10578; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10580 = 8'h54 == io_state_in_9 ? 8'hc2 : _GEN_10579; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10581 = 8'h55 == io_state_in_9 ? 8'hcb : _GEN_10580; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10582 = 8'h56 == io_state_in_9 ? 8'hd0 : _GEN_10581; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10583 = 8'h57 == io_state_in_9 ? 8'hd9 : _GEN_10582; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10584 = 8'h58 == io_state_in_9 ? 8'hae : _GEN_10583; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10585 = 8'h59 == io_state_in_9 ? 8'ha7 : _GEN_10584; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10586 = 8'h5a == io_state_in_9 ? 8'hbc : _GEN_10585; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10587 = 8'h5b == io_state_in_9 ? 8'hb5 : _GEN_10586; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10588 = 8'h5c == io_state_in_9 ? 8'h8a : _GEN_10587; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10589 = 8'h5d == io_state_in_9 ? 8'h83 : _GEN_10588; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10590 = 8'h5e == io_state_in_9 ? 8'h98 : _GEN_10589; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10591 = 8'h5f == io_state_in_9 ? 8'h91 : _GEN_10590; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10592 = 8'h60 == io_state_in_9 ? 8'h4d : _GEN_10591; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10593 = 8'h61 == io_state_in_9 ? 8'h44 : _GEN_10592; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10594 = 8'h62 == io_state_in_9 ? 8'h5f : _GEN_10593; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10595 = 8'h63 == io_state_in_9 ? 8'h56 : _GEN_10594; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10596 = 8'h64 == io_state_in_9 ? 8'h69 : _GEN_10595; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10597 = 8'h65 == io_state_in_9 ? 8'h60 : _GEN_10596; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10598 = 8'h66 == io_state_in_9 ? 8'h7b : _GEN_10597; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10599 = 8'h67 == io_state_in_9 ? 8'h72 : _GEN_10598; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10600 = 8'h68 == io_state_in_9 ? 8'h5 : _GEN_10599; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10601 = 8'h69 == io_state_in_9 ? 8'hc : _GEN_10600; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10602 = 8'h6a == io_state_in_9 ? 8'h17 : _GEN_10601; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10603 = 8'h6b == io_state_in_9 ? 8'h1e : _GEN_10602; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10604 = 8'h6c == io_state_in_9 ? 8'h21 : _GEN_10603; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10605 = 8'h6d == io_state_in_9 ? 8'h28 : _GEN_10604; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10606 = 8'h6e == io_state_in_9 ? 8'h33 : _GEN_10605; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10607 = 8'h6f == io_state_in_9 ? 8'h3a : _GEN_10606; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10608 = 8'h70 == io_state_in_9 ? 8'hdd : _GEN_10607; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10609 = 8'h71 == io_state_in_9 ? 8'hd4 : _GEN_10608; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10610 = 8'h72 == io_state_in_9 ? 8'hcf : _GEN_10609; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10611 = 8'h73 == io_state_in_9 ? 8'hc6 : _GEN_10610; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10612 = 8'h74 == io_state_in_9 ? 8'hf9 : _GEN_10611; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10613 = 8'h75 == io_state_in_9 ? 8'hf0 : _GEN_10612; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10614 = 8'h76 == io_state_in_9 ? 8'heb : _GEN_10613; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10615 = 8'h77 == io_state_in_9 ? 8'he2 : _GEN_10614; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10616 = 8'h78 == io_state_in_9 ? 8'h95 : _GEN_10615; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10617 = 8'h79 == io_state_in_9 ? 8'h9c : _GEN_10616; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10618 = 8'h7a == io_state_in_9 ? 8'h87 : _GEN_10617; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10619 = 8'h7b == io_state_in_9 ? 8'h8e : _GEN_10618; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10620 = 8'h7c == io_state_in_9 ? 8'hb1 : _GEN_10619; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10621 = 8'h7d == io_state_in_9 ? 8'hb8 : _GEN_10620; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10622 = 8'h7e == io_state_in_9 ? 8'ha3 : _GEN_10621; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10623 = 8'h7f == io_state_in_9 ? 8'haa : _GEN_10622; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10624 = 8'h80 == io_state_in_9 ? 8'hec : _GEN_10623; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10625 = 8'h81 == io_state_in_9 ? 8'he5 : _GEN_10624; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10626 = 8'h82 == io_state_in_9 ? 8'hfe : _GEN_10625; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10627 = 8'h83 == io_state_in_9 ? 8'hf7 : _GEN_10626; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10628 = 8'h84 == io_state_in_9 ? 8'hc8 : _GEN_10627; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10629 = 8'h85 == io_state_in_9 ? 8'hc1 : _GEN_10628; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10630 = 8'h86 == io_state_in_9 ? 8'hda : _GEN_10629; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10631 = 8'h87 == io_state_in_9 ? 8'hd3 : _GEN_10630; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10632 = 8'h88 == io_state_in_9 ? 8'ha4 : _GEN_10631; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10633 = 8'h89 == io_state_in_9 ? 8'had : _GEN_10632; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10634 = 8'h8a == io_state_in_9 ? 8'hb6 : _GEN_10633; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10635 = 8'h8b == io_state_in_9 ? 8'hbf : _GEN_10634; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10636 = 8'h8c == io_state_in_9 ? 8'h80 : _GEN_10635; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10637 = 8'h8d == io_state_in_9 ? 8'h89 : _GEN_10636; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10638 = 8'h8e == io_state_in_9 ? 8'h92 : _GEN_10637; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10639 = 8'h8f == io_state_in_9 ? 8'h9b : _GEN_10638; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10640 = 8'h90 == io_state_in_9 ? 8'h7c : _GEN_10639; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10641 = 8'h91 == io_state_in_9 ? 8'h75 : _GEN_10640; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10642 = 8'h92 == io_state_in_9 ? 8'h6e : _GEN_10641; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10643 = 8'h93 == io_state_in_9 ? 8'h67 : _GEN_10642; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10644 = 8'h94 == io_state_in_9 ? 8'h58 : _GEN_10643; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10645 = 8'h95 == io_state_in_9 ? 8'h51 : _GEN_10644; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10646 = 8'h96 == io_state_in_9 ? 8'h4a : _GEN_10645; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10647 = 8'h97 == io_state_in_9 ? 8'h43 : _GEN_10646; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10648 = 8'h98 == io_state_in_9 ? 8'h34 : _GEN_10647; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10649 = 8'h99 == io_state_in_9 ? 8'h3d : _GEN_10648; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10650 = 8'h9a == io_state_in_9 ? 8'h26 : _GEN_10649; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10651 = 8'h9b == io_state_in_9 ? 8'h2f : _GEN_10650; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10652 = 8'h9c == io_state_in_9 ? 8'h10 : _GEN_10651; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10653 = 8'h9d == io_state_in_9 ? 8'h19 : _GEN_10652; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10654 = 8'h9e == io_state_in_9 ? 8'h2 : _GEN_10653; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10655 = 8'h9f == io_state_in_9 ? 8'hb : _GEN_10654; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10656 = 8'ha0 == io_state_in_9 ? 8'hd7 : _GEN_10655; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10657 = 8'ha1 == io_state_in_9 ? 8'hde : _GEN_10656; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10658 = 8'ha2 == io_state_in_9 ? 8'hc5 : _GEN_10657; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10659 = 8'ha3 == io_state_in_9 ? 8'hcc : _GEN_10658; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10660 = 8'ha4 == io_state_in_9 ? 8'hf3 : _GEN_10659; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10661 = 8'ha5 == io_state_in_9 ? 8'hfa : _GEN_10660; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10662 = 8'ha6 == io_state_in_9 ? 8'he1 : _GEN_10661; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10663 = 8'ha7 == io_state_in_9 ? 8'he8 : _GEN_10662; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10664 = 8'ha8 == io_state_in_9 ? 8'h9f : _GEN_10663; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10665 = 8'ha9 == io_state_in_9 ? 8'h96 : _GEN_10664; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10666 = 8'haa == io_state_in_9 ? 8'h8d : _GEN_10665; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10667 = 8'hab == io_state_in_9 ? 8'h84 : _GEN_10666; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10668 = 8'hac == io_state_in_9 ? 8'hbb : _GEN_10667; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10669 = 8'had == io_state_in_9 ? 8'hb2 : _GEN_10668; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10670 = 8'hae == io_state_in_9 ? 8'ha9 : _GEN_10669; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10671 = 8'haf == io_state_in_9 ? 8'ha0 : _GEN_10670; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10672 = 8'hb0 == io_state_in_9 ? 8'h47 : _GEN_10671; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10673 = 8'hb1 == io_state_in_9 ? 8'h4e : _GEN_10672; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10674 = 8'hb2 == io_state_in_9 ? 8'h55 : _GEN_10673; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10675 = 8'hb3 == io_state_in_9 ? 8'h5c : _GEN_10674; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10676 = 8'hb4 == io_state_in_9 ? 8'h63 : _GEN_10675; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10677 = 8'hb5 == io_state_in_9 ? 8'h6a : _GEN_10676; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10678 = 8'hb6 == io_state_in_9 ? 8'h71 : _GEN_10677; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10679 = 8'hb7 == io_state_in_9 ? 8'h78 : _GEN_10678; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10680 = 8'hb8 == io_state_in_9 ? 8'hf : _GEN_10679; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10681 = 8'hb9 == io_state_in_9 ? 8'h6 : _GEN_10680; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10682 = 8'hba == io_state_in_9 ? 8'h1d : _GEN_10681; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10683 = 8'hbb == io_state_in_9 ? 8'h14 : _GEN_10682; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10684 = 8'hbc == io_state_in_9 ? 8'h2b : _GEN_10683; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10685 = 8'hbd == io_state_in_9 ? 8'h22 : _GEN_10684; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10686 = 8'hbe == io_state_in_9 ? 8'h39 : _GEN_10685; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10687 = 8'hbf == io_state_in_9 ? 8'h30 : _GEN_10686; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10688 = 8'hc0 == io_state_in_9 ? 8'h9a : _GEN_10687; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10689 = 8'hc1 == io_state_in_9 ? 8'h93 : _GEN_10688; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10690 = 8'hc2 == io_state_in_9 ? 8'h88 : _GEN_10689; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10691 = 8'hc3 == io_state_in_9 ? 8'h81 : _GEN_10690; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10692 = 8'hc4 == io_state_in_9 ? 8'hbe : _GEN_10691; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10693 = 8'hc5 == io_state_in_9 ? 8'hb7 : _GEN_10692; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10694 = 8'hc6 == io_state_in_9 ? 8'hac : _GEN_10693; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10695 = 8'hc7 == io_state_in_9 ? 8'ha5 : _GEN_10694; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10696 = 8'hc8 == io_state_in_9 ? 8'hd2 : _GEN_10695; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10697 = 8'hc9 == io_state_in_9 ? 8'hdb : _GEN_10696; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10698 = 8'hca == io_state_in_9 ? 8'hc0 : _GEN_10697; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10699 = 8'hcb == io_state_in_9 ? 8'hc9 : _GEN_10698; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10700 = 8'hcc == io_state_in_9 ? 8'hf6 : _GEN_10699; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10701 = 8'hcd == io_state_in_9 ? 8'hff : _GEN_10700; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10702 = 8'hce == io_state_in_9 ? 8'he4 : _GEN_10701; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10703 = 8'hcf == io_state_in_9 ? 8'hed : _GEN_10702; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10704 = 8'hd0 == io_state_in_9 ? 8'ha : _GEN_10703; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10705 = 8'hd1 == io_state_in_9 ? 8'h3 : _GEN_10704; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10706 = 8'hd2 == io_state_in_9 ? 8'h18 : _GEN_10705; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10707 = 8'hd3 == io_state_in_9 ? 8'h11 : _GEN_10706; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10708 = 8'hd4 == io_state_in_9 ? 8'h2e : _GEN_10707; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10709 = 8'hd5 == io_state_in_9 ? 8'h27 : _GEN_10708; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10710 = 8'hd6 == io_state_in_9 ? 8'h3c : _GEN_10709; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10711 = 8'hd7 == io_state_in_9 ? 8'h35 : _GEN_10710; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10712 = 8'hd8 == io_state_in_9 ? 8'h42 : _GEN_10711; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10713 = 8'hd9 == io_state_in_9 ? 8'h4b : _GEN_10712; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10714 = 8'hda == io_state_in_9 ? 8'h50 : _GEN_10713; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10715 = 8'hdb == io_state_in_9 ? 8'h59 : _GEN_10714; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10716 = 8'hdc == io_state_in_9 ? 8'h66 : _GEN_10715; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10717 = 8'hdd == io_state_in_9 ? 8'h6f : _GEN_10716; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10718 = 8'hde == io_state_in_9 ? 8'h74 : _GEN_10717; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10719 = 8'hdf == io_state_in_9 ? 8'h7d : _GEN_10718; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10720 = 8'he0 == io_state_in_9 ? 8'ha1 : _GEN_10719; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10721 = 8'he1 == io_state_in_9 ? 8'ha8 : _GEN_10720; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10722 = 8'he2 == io_state_in_9 ? 8'hb3 : _GEN_10721; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10723 = 8'he3 == io_state_in_9 ? 8'hba : _GEN_10722; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10724 = 8'he4 == io_state_in_9 ? 8'h85 : _GEN_10723; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10725 = 8'he5 == io_state_in_9 ? 8'h8c : _GEN_10724; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10726 = 8'he6 == io_state_in_9 ? 8'h97 : _GEN_10725; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10727 = 8'he7 == io_state_in_9 ? 8'h9e : _GEN_10726; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10728 = 8'he8 == io_state_in_9 ? 8'he9 : _GEN_10727; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10729 = 8'he9 == io_state_in_9 ? 8'he0 : _GEN_10728; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10730 = 8'hea == io_state_in_9 ? 8'hfb : _GEN_10729; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10731 = 8'heb == io_state_in_9 ? 8'hf2 : _GEN_10730; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10732 = 8'hec == io_state_in_9 ? 8'hcd : _GEN_10731; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10733 = 8'hed == io_state_in_9 ? 8'hc4 : _GEN_10732; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10734 = 8'hee == io_state_in_9 ? 8'hdf : _GEN_10733; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10735 = 8'hef == io_state_in_9 ? 8'hd6 : _GEN_10734; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10736 = 8'hf0 == io_state_in_9 ? 8'h31 : _GEN_10735; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10737 = 8'hf1 == io_state_in_9 ? 8'h38 : _GEN_10736; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10738 = 8'hf2 == io_state_in_9 ? 8'h23 : _GEN_10737; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10739 = 8'hf3 == io_state_in_9 ? 8'h2a : _GEN_10738; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10740 = 8'hf4 == io_state_in_9 ? 8'h15 : _GEN_10739; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10741 = 8'hf5 == io_state_in_9 ? 8'h1c : _GEN_10740; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10742 = 8'hf6 == io_state_in_9 ? 8'h7 : _GEN_10741; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10743 = 8'hf7 == io_state_in_9 ? 8'he : _GEN_10742; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10744 = 8'hf8 == io_state_in_9 ? 8'h79 : _GEN_10743; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10745 = 8'hf9 == io_state_in_9 ? 8'h70 : _GEN_10744; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10746 = 8'hfa == io_state_in_9 ? 8'h6b : _GEN_10745; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10747 = 8'hfb == io_state_in_9 ? 8'h62 : _GEN_10746; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10748 = 8'hfc == io_state_in_9 ? 8'h5d : _GEN_10747; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10749 = 8'hfd == io_state_in_9 ? 8'h54 : _GEN_10748; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10750 = 8'hfe == io_state_in_9 ? 8'h4f : _GEN_10749; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_10751 = 8'hff == io_state_in_9 ? 8'h46 : _GEN_10750; // @[InvMixColumns.scala 138:{42,42}]
  wire [7:0] _tmp_state_10_T = _GEN_10495 ^ _GEN_10751; // @[InvMixColumns.scala 138:42]
  wire [7:0] _GEN_10753 = 8'h1 == io_state_in_10 ? 8'he : 8'h0; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10754 = 8'h2 == io_state_in_10 ? 8'h1c : _GEN_10753; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10755 = 8'h3 == io_state_in_10 ? 8'h12 : _GEN_10754; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10756 = 8'h4 == io_state_in_10 ? 8'h38 : _GEN_10755; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10757 = 8'h5 == io_state_in_10 ? 8'h36 : _GEN_10756; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10758 = 8'h6 == io_state_in_10 ? 8'h24 : _GEN_10757; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10759 = 8'h7 == io_state_in_10 ? 8'h2a : _GEN_10758; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10760 = 8'h8 == io_state_in_10 ? 8'h70 : _GEN_10759; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10761 = 8'h9 == io_state_in_10 ? 8'h7e : _GEN_10760; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10762 = 8'ha == io_state_in_10 ? 8'h6c : _GEN_10761; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10763 = 8'hb == io_state_in_10 ? 8'h62 : _GEN_10762; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10764 = 8'hc == io_state_in_10 ? 8'h48 : _GEN_10763; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10765 = 8'hd == io_state_in_10 ? 8'h46 : _GEN_10764; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10766 = 8'he == io_state_in_10 ? 8'h54 : _GEN_10765; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10767 = 8'hf == io_state_in_10 ? 8'h5a : _GEN_10766; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10768 = 8'h10 == io_state_in_10 ? 8'he0 : _GEN_10767; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10769 = 8'h11 == io_state_in_10 ? 8'hee : _GEN_10768; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10770 = 8'h12 == io_state_in_10 ? 8'hfc : _GEN_10769; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10771 = 8'h13 == io_state_in_10 ? 8'hf2 : _GEN_10770; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10772 = 8'h14 == io_state_in_10 ? 8'hd8 : _GEN_10771; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10773 = 8'h15 == io_state_in_10 ? 8'hd6 : _GEN_10772; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10774 = 8'h16 == io_state_in_10 ? 8'hc4 : _GEN_10773; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10775 = 8'h17 == io_state_in_10 ? 8'hca : _GEN_10774; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10776 = 8'h18 == io_state_in_10 ? 8'h90 : _GEN_10775; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10777 = 8'h19 == io_state_in_10 ? 8'h9e : _GEN_10776; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10778 = 8'h1a == io_state_in_10 ? 8'h8c : _GEN_10777; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10779 = 8'h1b == io_state_in_10 ? 8'h82 : _GEN_10778; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10780 = 8'h1c == io_state_in_10 ? 8'ha8 : _GEN_10779; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10781 = 8'h1d == io_state_in_10 ? 8'ha6 : _GEN_10780; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10782 = 8'h1e == io_state_in_10 ? 8'hb4 : _GEN_10781; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10783 = 8'h1f == io_state_in_10 ? 8'hba : _GEN_10782; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10784 = 8'h20 == io_state_in_10 ? 8'hdb : _GEN_10783; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10785 = 8'h21 == io_state_in_10 ? 8'hd5 : _GEN_10784; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10786 = 8'h22 == io_state_in_10 ? 8'hc7 : _GEN_10785; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10787 = 8'h23 == io_state_in_10 ? 8'hc9 : _GEN_10786; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10788 = 8'h24 == io_state_in_10 ? 8'he3 : _GEN_10787; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10789 = 8'h25 == io_state_in_10 ? 8'hed : _GEN_10788; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10790 = 8'h26 == io_state_in_10 ? 8'hff : _GEN_10789; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10791 = 8'h27 == io_state_in_10 ? 8'hf1 : _GEN_10790; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10792 = 8'h28 == io_state_in_10 ? 8'hab : _GEN_10791; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10793 = 8'h29 == io_state_in_10 ? 8'ha5 : _GEN_10792; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10794 = 8'h2a == io_state_in_10 ? 8'hb7 : _GEN_10793; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10795 = 8'h2b == io_state_in_10 ? 8'hb9 : _GEN_10794; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10796 = 8'h2c == io_state_in_10 ? 8'h93 : _GEN_10795; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10797 = 8'h2d == io_state_in_10 ? 8'h9d : _GEN_10796; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10798 = 8'h2e == io_state_in_10 ? 8'h8f : _GEN_10797; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10799 = 8'h2f == io_state_in_10 ? 8'h81 : _GEN_10798; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10800 = 8'h30 == io_state_in_10 ? 8'h3b : _GEN_10799; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10801 = 8'h31 == io_state_in_10 ? 8'h35 : _GEN_10800; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10802 = 8'h32 == io_state_in_10 ? 8'h27 : _GEN_10801; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10803 = 8'h33 == io_state_in_10 ? 8'h29 : _GEN_10802; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10804 = 8'h34 == io_state_in_10 ? 8'h3 : _GEN_10803; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10805 = 8'h35 == io_state_in_10 ? 8'hd : _GEN_10804; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10806 = 8'h36 == io_state_in_10 ? 8'h1f : _GEN_10805; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10807 = 8'h37 == io_state_in_10 ? 8'h11 : _GEN_10806; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10808 = 8'h38 == io_state_in_10 ? 8'h4b : _GEN_10807; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10809 = 8'h39 == io_state_in_10 ? 8'h45 : _GEN_10808; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10810 = 8'h3a == io_state_in_10 ? 8'h57 : _GEN_10809; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10811 = 8'h3b == io_state_in_10 ? 8'h59 : _GEN_10810; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10812 = 8'h3c == io_state_in_10 ? 8'h73 : _GEN_10811; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10813 = 8'h3d == io_state_in_10 ? 8'h7d : _GEN_10812; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10814 = 8'h3e == io_state_in_10 ? 8'h6f : _GEN_10813; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10815 = 8'h3f == io_state_in_10 ? 8'h61 : _GEN_10814; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10816 = 8'h40 == io_state_in_10 ? 8'had : _GEN_10815; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10817 = 8'h41 == io_state_in_10 ? 8'ha3 : _GEN_10816; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10818 = 8'h42 == io_state_in_10 ? 8'hb1 : _GEN_10817; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10819 = 8'h43 == io_state_in_10 ? 8'hbf : _GEN_10818; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10820 = 8'h44 == io_state_in_10 ? 8'h95 : _GEN_10819; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10821 = 8'h45 == io_state_in_10 ? 8'h9b : _GEN_10820; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10822 = 8'h46 == io_state_in_10 ? 8'h89 : _GEN_10821; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10823 = 8'h47 == io_state_in_10 ? 8'h87 : _GEN_10822; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10824 = 8'h48 == io_state_in_10 ? 8'hdd : _GEN_10823; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10825 = 8'h49 == io_state_in_10 ? 8'hd3 : _GEN_10824; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10826 = 8'h4a == io_state_in_10 ? 8'hc1 : _GEN_10825; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10827 = 8'h4b == io_state_in_10 ? 8'hcf : _GEN_10826; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10828 = 8'h4c == io_state_in_10 ? 8'he5 : _GEN_10827; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10829 = 8'h4d == io_state_in_10 ? 8'heb : _GEN_10828; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10830 = 8'h4e == io_state_in_10 ? 8'hf9 : _GEN_10829; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10831 = 8'h4f == io_state_in_10 ? 8'hf7 : _GEN_10830; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10832 = 8'h50 == io_state_in_10 ? 8'h4d : _GEN_10831; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10833 = 8'h51 == io_state_in_10 ? 8'h43 : _GEN_10832; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10834 = 8'h52 == io_state_in_10 ? 8'h51 : _GEN_10833; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10835 = 8'h53 == io_state_in_10 ? 8'h5f : _GEN_10834; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10836 = 8'h54 == io_state_in_10 ? 8'h75 : _GEN_10835; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10837 = 8'h55 == io_state_in_10 ? 8'h7b : _GEN_10836; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10838 = 8'h56 == io_state_in_10 ? 8'h69 : _GEN_10837; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10839 = 8'h57 == io_state_in_10 ? 8'h67 : _GEN_10838; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10840 = 8'h58 == io_state_in_10 ? 8'h3d : _GEN_10839; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10841 = 8'h59 == io_state_in_10 ? 8'h33 : _GEN_10840; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10842 = 8'h5a == io_state_in_10 ? 8'h21 : _GEN_10841; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10843 = 8'h5b == io_state_in_10 ? 8'h2f : _GEN_10842; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10844 = 8'h5c == io_state_in_10 ? 8'h5 : _GEN_10843; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10845 = 8'h5d == io_state_in_10 ? 8'hb : _GEN_10844; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10846 = 8'h5e == io_state_in_10 ? 8'h19 : _GEN_10845; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10847 = 8'h5f == io_state_in_10 ? 8'h17 : _GEN_10846; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10848 = 8'h60 == io_state_in_10 ? 8'h76 : _GEN_10847; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10849 = 8'h61 == io_state_in_10 ? 8'h78 : _GEN_10848; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10850 = 8'h62 == io_state_in_10 ? 8'h6a : _GEN_10849; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10851 = 8'h63 == io_state_in_10 ? 8'h64 : _GEN_10850; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10852 = 8'h64 == io_state_in_10 ? 8'h4e : _GEN_10851; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10853 = 8'h65 == io_state_in_10 ? 8'h40 : _GEN_10852; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10854 = 8'h66 == io_state_in_10 ? 8'h52 : _GEN_10853; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10855 = 8'h67 == io_state_in_10 ? 8'h5c : _GEN_10854; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10856 = 8'h68 == io_state_in_10 ? 8'h6 : _GEN_10855; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10857 = 8'h69 == io_state_in_10 ? 8'h8 : _GEN_10856; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10858 = 8'h6a == io_state_in_10 ? 8'h1a : _GEN_10857; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10859 = 8'h6b == io_state_in_10 ? 8'h14 : _GEN_10858; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10860 = 8'h6c == io_state_in_10 ? 8'h3e : _GEN_10859; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10861 = 8'h6d == io_state_in_10 ? 8'h30 : _GEN_10860; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10862 = 8'h6e == io_state_in_10 ? 8'h22 : _GEN_10861; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10863 = 8'h6f == io_state_in_10 ? 8'h2c : _GEN_10862; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10864 = 8'h70 == io_state_in_10 ? 8'h96 : _GEN_10863; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10865 = 8'h71 == io_state_in_10 ? 8'h98 : _GEN_10864; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10866 = 8'h72 == io_state_in_10 ? 8'h8a : _GEN_10865; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10867 = 8'h73 == io_state_in_10 ? 8'h84 : _GEN_10866; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10868 = 8'h74 == io_state_in_10 ? 8'hae : _GEN_10867; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10869 = 8'h75 == io_state_in_10 ? 8'ha0 : _GEN_10868; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10870 = 8'h76 == io_state_in_10 ? 8'hb2 : _GEN_10869; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10871 = 8'h77 == io_state_in_10 ? 8'hbc : _GEN_10870; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10872 = 8'h78 == io_state_in_10 ? 8'he6 : _GEN_10871; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10873 = 8'h79 == io_state_in_10 ? 8'he8 : _GEN_10872; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10874 = 8'h7a == io_state_in_10 ? 8'hfa : _GEN_10873; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10875 = 8'h7b == io_state_in_10 ? 8'hf4 : _GEN_10874; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10876 = 8'h7c == io_state_in_10 ? 8'hde : _GEN_10875; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10877 = 8'h7d == io_state_in_10 ? 8'hd0 : _GEN_10876; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10878 = 8'h7e == io_state_in_10 ? 8'hc2 : _GEN_10877; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10879 = 8'h7f == io_state_in_10 ? 8'hcc : _GEN_10878; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10880 = 8'h80 == io_state_in_10 ? 8'h41 : _GEN_10879; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10881 = 8'h81 == io_state_in_10 ? 8'h4f : _GEN_10880; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10882 = 8'h82 == io_state_in_10 ? 8'h5d : _GEN_10881; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10883 = 8'h83 == io_state_in_10 ? 8'h53 : _GEN_10882; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10884 = 8'h84 == io_state_in_10 ? 8'h79 : _GEN_10883; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10885 = 8'h85 == io_state_in_10 ? 8'h77 : _GEN_10884; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10886 = 8'h86 == io_state_in_10 ? 8'h65 : _GEN_10885; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10887 = 8'h87 == io_state_in_10 ? 8'h6b : _GEN_10886; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10888 = 8'h88 == io_state_in_10 ? 8'h31 : _GEN_10887; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10889 = 8'h89 == io_state_in_10 ? 8'h3f : _GEN_10888; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10890 = 8'h8a == io_state_in_10 ? 8'h2d : _GEN_10889; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10891 = 8'h8b == io_state_in_10 ? 8'h23 : _GEN_10890; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10892 = 8'h8c == io_state_in_10 ? 8'h9 : _GEN_10891; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10893 = 8'h8d == io_state_in_10 ? 8'h7 : _GEN_10892; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10894 = 8'h8e == io_state_in_10 ? 8'h15 : _GEN_10893; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10895 = 8'h8f == io_state_in_10 ? 8'h1b : _GEN_10894; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10896 = 8'h90 == io_state_in_10 ? 8'ha1 : _GEN_10895; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10897 = 8'h91 == io_state_in_10 ? 8'haf : _GEN_10896; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10898 = 8'h92 == io_state_in_10 ? 8'hbd : _GEN_10897; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10899 = 8'h93 == io_state_in_10 ? 8'hb3 : _GEN_10898; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10900 = 8'h94 == io_state_in_10 ? 8'h99 : _GEN_10899; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10901 = 8'h95 == io_state_in_10 ? 8'h97 : _GEN_10900; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10902 = 8'h96 == io_state_in_10 ? 8'h85 : _GEN_10901; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10903 = 8'h97 == io_state_in_10 ? 8'h8b : _GEN_10902; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10904 = 8'h98 == io_state_in_10 ? 8'hd1 : _GEN_10903; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10905 = 8'h99 == io_state_in_10 ? 8'hdf : _GEN_10904; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10906 = 8'h9a == io_state_in_10 ? 8'hcd : _GEN_10905; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10907 = 8'h9b == io_state_in_10 ? 8'hc3 : _GEN_10906; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10908 = 8'h9c == io_state_in_10 ? 8'he9 : _GEN_10907; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10909 = 8'h9d == io_state_in_10 ? 8'he7 : _GEN_10908; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10910 = 8'h9e == io_state_in_10 ? 8'hf5 : _GEN_10909; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10911 = 8'h9f == io_state_in_10 ? 8'hfb : _GEN_10910; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10912 = 8'ha0 == io_state_in_10 ? 8'h9a : _GEN_10911; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10913 = 8'ha1 == io_state_in_10 ? 8'h94 : _GEN_10912; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10914 = 8'ha2 == io_state_in_10 ? 8'h86 : _GEN_10913; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10915 = 8'ha3 == io_state_in_10 ? 8'h88 : _GEN_10914; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10916 = 8'ha4 == io_state_in_10 ? 8'ha2 : _GEN_10915; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10917 = 8'ha5 == io_state_in_10 ? 8'hac : _GEN_10916; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10918 = 8'ha6 == io_state_in_10 ? 8'hbe : _GEN_10917; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10919 = 8'ha7 == io_state_in_10 ? 8'hb0 : _GEN_10918; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10920 = 8'ha8 == io_state_in_10 ? 8'hea : _GEN_10919; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10921 = 8'ha9 == io_state_in_10 ? 8'he4 : _GEN_10920; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10922 = 8'haa == io_state_in_10 ? 8'hf6 : _GEN_10921; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10923 = 8'hab == io_state_in_10 ? 8'hf8 : _GEN_10922; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10924 = 8'hac == io_state_in_10 ? 8'hd2 : _GEN_10923; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10925 = 8'had == io_state_in_10 ? 8'hdc : _GEN_10924; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10926 = 8'hae == io_state_in_10 ? 8'hce : _GEN_10925; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10927 = 8'haf == io_state_in_10 ? 8'hc0 : _GEN_10926; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10928 = 8'hb0 == io_state_in_10 ? 8'h7a : _GEN_10927; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10929 = 8'hb1 == io_state_in_10 ? 8'h74 : _GEN_10928; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10930 = 8'hb2 == io_state_in_10 ? 8'h66 : _GEN_10929; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10931 = 8'hb3 == io_state_in_10 ? 8'h68 : _GEN_10930; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10932 = 8'hb4 == io_state_in_10 ? 8'h42 : _GEN_10931; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10933 = 8'hb5 == io_state_in_10 ? 8'h4c : _GEN_10932; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10934 = 8'hb6 == io_state_in_10 ? 8'h5e : _GEN_10933; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10935 = 8'hb7 == io_state_in_10 ? 8'h50 : _GEN_10934; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10936 = 8'hb8 == io_state_in_10 ? 8'ha : _GEN_10935; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10937 = 8'hb9 == io_state_in_10 ? 8'h4 : _GEN_10936; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10938 = 8'hba == io_state_in_10 ? 8'h16 : _GEN_10937; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10939 = 8'hbb == io_state_in_10 ? 8'h18 : _GEN_10938; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10940 = 8'hbc == io_state_in_10 ? 8'h32 : _GEN_10939; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10941 = 8'hbd == io_state_in_10 ? 8'h3c : _GEN_10940; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10942 = 8'hbe == io_state_in_10 ? 8'h2e : _GEN_10941; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10943 = 8'hbf == io_state_in_10 ? 8'h20 : _GEN_10942; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10944 = 8'hc0 == io_state_in_10 ? 8'hec : _GEN_10943; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10945 = 8'hc1 == io_state_in_10 ? 8'he2 : _GEN_10944; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10946 = 8'hc2 == io_state_in_10 ? 8'hf0 : _GEN_10945; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10947 = 8'hc3 == io_state_in_10 ? 8'hfe : _GEN_10946; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10948 = 8'hc4 == io_state_in_10 ? 8'hd4 : _GEN_10947; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10949 = 8'hc5 == io_state_in_10 ? 8'hda : _GEN_10948; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10950 = 8'hc6 == io_state_in_10 ? 8'hc8 : _GEN_10949; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10951 = 8'hc7 == io_state_in_10 ? 8'hc6 : _GEN_10950; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10952 = 8'hc8 == io_state_in_10 ? 8'h9c : _GEN_10951; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10953 = 8'hc9 == io_state_in_10 ? 8'h92 : _GEN_10952; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10954 = 8'hca == io_state_in_10 ? 8'h80 : _GEN_10953; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10955 = 8'hcb == io_state_in_10 ? 8'h8e : _GEN_10954; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10956 = 8'hcc == io_state_in_10 ? 8'ha4 : _GEN_10955; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10957 = 8'hcd == io_state_in_10 ? 8'haa : _GEN_10956; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10958 = 8'hce == io_state_in_10 ? 8'hb8 : _GEN_10957; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10959 = 8'hcf == io_state_in_10 ? 8'hb6 : _GEN_10958; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10960 = 8'hd0 == io_state_in_10 ? 8'hc : _GEN_10959; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10961 = 8'hd1 == io_state_in_10 ? 8'h2 : _GEN_10960; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10962 = 8'hd2 == io_state_in_10 ? 8'h10 : _GEN_10961; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10963 = 8'hd3 == io_state_in_10 ? 8'h1e : _GEN_10962; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10964 = 8'hd4 == io_state_in_10 ? 8'h34 : _GEN_10963; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10965 = 8'hd5 == io_state_in_10 ? 8'h3a : _GEN_10964; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10966 = 8'hd6 == io_state_in_10 ? 8'h28 : _GEN_10965; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10967 = 8'hd7 == io_state_in_10 ? 8'h26 : _GEN_10966; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10968 = 8'hd8 == io_state_in_10 ? 8'h7c : _GEN_10967; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10969 = 8'hd9 == io_state_in_10 ? 8'h72 : _GEN_10968; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10970 = 8'hda == io_state_in_10 ? 8'h60 : _GEN_10969; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10971 = 8'hdb == io_state_in_10 ? 8'h6e : _GEN_10970; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10972 = 8'hdc == io_state_in_10 ? 8'h44 : _GEN_10971; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10973 = 8'hdd == io_state_in_10 ? 8'h4a : _GEN_10972; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10974 = 8'hde == io_state_in_10 ? 8'h58 : _GEN_10973; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10975 = 8'hdf == io_state_in_10 ? 8'h56 : _GEN_10974; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10976 = 8'he0 == io_state_in_10 ? 8'h37 : _GEN_10975; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10977 = 8'he1 == io_state_in_10 ? 8'h39 : _GEN_10976; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10978 = 8'he2 == io_state_in_10 ? 8'h2b : _GEN_10977; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10979 = 8'he3 == io_state_in_10 ? 8'h25 : _GEN_10978; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10980 = 8'he4 == io_state_in_10 ? 8'hf : _GEN_10979; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10981 = 8'he5 == io_state_in_10 ? 8'h1 : _GEN_10980; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10982 = 8'he6 == io_state_in_10 ? 8'h13 : _GEN_10981; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10983 = 8'he7 == io_state_in_10 ? 8'h1d : _GEN_10982; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10984 = 8'he8 == io_state_in_10 ? 8'h47 : _GEN_10983; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10985 = 8'he9 == io_state_in_10 ? 8'h49 : _GEN_10984; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10986 = 8'hea == io_state_in_10 ? 8'h5b : _GEN_10985; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10987 = 8'heb == io_state_in_10 ? 8'h55 : _GEN_10986; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10988 = 8'hec == io_state_in_10 ? 8'h7f : _GEN_10987; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10989 = 8'hed == io_state_in_10 ? 8'h71 : _GEN_10988; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10990 = 8'hee == io_state_in_10 ? 8'h63 : _GEN_10989; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10991 = 8'hef == io_state_in_10 ? 8'h6d : _GEN_10990; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10992 = 8'hf0 == io_state_in_10 ? 8'hd7 : _GEN_10991; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10993 = 8'hf1 == io_state_in_10 ? 8'hd9 : _GEN_10992; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10994 = 8'hf2 == io_state_in_10 ? 8'hcb : _GEN_10993; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10995 = 8'hf3 == io_state_in_10 ? 8'hc5 : _GEN_10994; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10996 = 8'hf4 == io_state_in_10 ? 8'hef : _GEN_10995; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10997 = 8'hf5 == io_state_in_10 ? 8'he1 : _GEN_10996; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10998 = 8'hf6 == io_state_in_10 ? 8'hf3 : _GEN_10997; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_10999 = 8'hf7 == io_state_in_10 ? 8'hfd : _GEN_10998; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11000 = 8'hf8 == io_state_in_10 ? 8'ha7 : _GEN_10999; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11001 = 8'hf9 == io_state_in_10 ? 8'ha9 : _GEN_11000; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11002 = 8'hfa == io_state_in_10 ? 8'hbb : _GEN_11001; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11003 = 8'hfb == io_state_in_10 ? 8'hb5 : _GEN_11002; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11004 = 8'hfc == io_state_in_10 ? 8'h9f : _GEN_11003; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11005 = 8'hfd == io_state_in_10 ? 8'h91 : _GEN_11004; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11006 = 8'hfe == io_state_in_10 ? 8'h83 : _GEN_11005; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _GEN_11007 = 8'hff == io_state_in_10 ? 8'h8d : _GEN_11006; // @[InvMixColumns.scala 138:{66,66}]
  wire [7:0] _tmp_state_10_T_1 = _tmp_state_10_T ^ _GEN_11007; // @[InvMixColumns.scala 138:66]
  wire [7:0] _GEN_11009 = 8'h1 == io_state_in_11 ? 8'hb : 8'h0; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11010 = 8'h2 == io_state_in_11 ? 8'h16 : _GEN_11009; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11011 = 8'h3 == io_state_in_11 ? 8'h1d : _GEN_11010; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11012 = 8'h4 == io_state_in_11 ? 8'h2c : _GEN_11011; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11013 = 8'h5 == io_state_in_11 ? 8'h27 : _GEN_11012; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11014 = 8'h6 == io_state_in_11 ? 8'h3a : _GEN_11013; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11015 = 8'h7 == io_state_in_11 ? 8'h31 : _GEN_11014; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11016 = 8'h8 == io_state_in_11 ? 8'h58 : _GEN_11015; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11017 = 8'h9 == io_state_in_11 ? 8'h53 : _GEN_11016; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11018 = 8'ha == io_state_in_11 ? 8'h4e : _GEN_11017; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11019 = 8'hb == io_state_in_11 ? 8'h45 : _GEN_11018; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11020 = 8'hc == io_state_in_11 ? 8'h74 : _GEN_11019; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11021 = 8'hd == io_state_in_11 ? 8'h7f : _GEN_11020; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11022 = 8'he == io_state_in_11 ? 8'h62 : _GEN_11021; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11023 = 8'hf == io_state_in_11 ? 8'h69 : _GEN_11022; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11024 = 8'h10 == io_state_in_11 ? 8'hb0 : _GEN_11023; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11025 = 8'h11 == io_state_in_11 ? 8'hbb : _GEN_11024; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11026 = 8'h12 == io_state_in_11 ? 8'ha6 : _GEN_11025; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11027 = 8'h13 == io_state_in_11 ? 8'had : _GEN_11026; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11028 = 8'h14 == io_state_in_11 ? 8'h9c : _GEN_11027; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11029 = 8'h15 == io_state_in_11 ? 8'h97 : _GEN_11028; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11030 = 8'h16 == io_state_in_11 ? 8'h8a : _GEN_11029; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11031 = 8'h17 == io_state_in_11 ? 8'h81 : _GEN_11030; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11032 = 8'h18 == io_state_in_11 ? 8'he8 : _GEN_11031; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11033 = 8'h19 == io_state_in_11 ? 8'he3 : _GEN_11032; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11034 = 8'h1a == io_state_in_11 ? 8'hfe : _GEN_11033; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11035 = 8'h1b == io_state_in_11 ? 8'hf5 : _GEN_11034; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11036 = 8'h1c == io_state_in_11 ? 8'hc4 : _GEN_11035; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11037 = 8'h1d == io_state_in_11 ? 8'hcf : _GEN_11036; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11038 = 8'h1e == io_state_in_11 ? 8'hd2 : _GEN_11037; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11039 = 8'h1f == io_state_in_11 ? 8'hd9 : _GEN_11038; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11040 = 8'h20 == io_state_in_11 ? 8'h7b : _GEN_11039; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11041 = 8'h21 == io_state_in_11 ? 8'h70 : _GEN_11040; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11042 = 8'h22 == io_state_in_11 ? 8'h6d : _GEN_11041; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11043 = 8'h23 == io_state_in_11 ? 8'h66 : _GEN_11042; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11044 = 8'h24 == io_state_in_11 ? 8'h57 : _GEN_11043; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11045 = 8'h25 == io_state_in_11 ? 8'h5c : _GEN_11044; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11046 = 8'h26 == io_state_in_11 ? 8'h41 : _GEN_11045; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11047 = 8'h27 == io_state_in_11 ? 8'h4a : _GEN_11046; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11048 = 8'h28 == io_state_in_11 ? 8'h23 : _GEN_11047; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11049 = 8'h29 == io_state_in_11 ? 8'h28 : _GEN_11048; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11050 = 8'h2a == io_state_in_11 ? 8'h35 : _GEN_11049; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11051 = 8'h2b == io_state_in_11 ? 8'h3e : _GEN_11050; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11052 = 8'h2c == io_state_in_11 ? 8'hf : _GEN_11051; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11053 = 8'h2d == io_state_in_11 ? 8'h4 : _GEN_11052; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11054 = 8'h2e == io_state_in_11 ? 8'h19 : _GEN_11053; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11055 = 8'h2f == io_state_in_11 ? 8'h12 : _GEN_11054; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11056 = 8'h30 == io_state_in_11 ? 8'hcb : _GEN_11055; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11057 = 8'h31 == io_state_in_11 ? 8'hc0 : _GEN_11056; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11058 = 8'h32 == io_state_in_11 ? 8'hdd : _GEN_11057; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11059 = 8'h33 == io_state_in_11 ? 8'hd6 : _GEN_11058; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11060 = 8'h34 == io_state_in_11 ? 8'he7 : _GEN_11059; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11061 = 8'h35 == io_state_in_11 ? 8'hec : _GEN_11060; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11062 = 8'h36 == io_state_in_11 ? 8'hf1 : _GEN_11061; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11063 = 8'h37 == io_state_in_11 ? 8'hfa : _GEN_11062; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11064 = 8'h38 == io_state_in_11 ? 8'h93 : _GEN_11063; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11065 = 8'h39 == io_state_in_11 ? 8'h98 : _GEN_11064; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11066 = 8'h3a == io_state_in_11 ? 8'h85 : _GEN_11065; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11067 = 8'h3b == io_state_in_11 ? 8'h8e : _GEN_11066; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11068 = 8'h3c == io_state_in_11 ? 8'hbf : _GEN_11067; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11069 = 8'h3d == io_state_in_11 ? 8'hb4 : _GEN_11068; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11070 = 8'h3e == io_state_in_11 ? 8'ha9 : _GEN_11069; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11071 = 8'h3f == io_state_in_11 ? 8'ha2 : _GEN_11070; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11072 = 8'h40 == io_state_in_11 ? 8'hf6 : _GEN_11071; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11073 = 8'h41 == io_state_in_11 ? 8'hfd : _GEN_11072; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11074 = 8'h42 == io_state_in_11 ? 8'he0 : _GEN_11073; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11075 = 8'h43 == io_state_in_11 ? 8'heb : _GEN_11074; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11076 = 8'h44 == io_state_in_11 ? 8'hda : _GEN_11075; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11077 = 8'h45 == io_state_in_11 ? 8'hd1 : _GEN_11076; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11078 = 8'h46 == io_state_in_11 ? 8'hcc : _GEN_11077; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11079 = 8'h47 == io_state_in_11 ? 8'hc7 : _GEN_11078; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11080 = 8'h48 == io_state_in_11 ? 8'hae : _GEN_11079; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11081 = 8'h49 == io_state_in_11 ? 8'ha5 : _GEN_11080; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11082 = 8'h4a == io_state_in_11 ? 8'hb8 : _GEN_11081; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11083 = 8'h4b == io_state_in_11 ? 8'hb3 : _GEN_11082; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11084 = 8'h4c == io_state_in_11 ? 8'h82 : _GEN_11083; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11085 = 8'h4d == io_state_in_11 ? 8'h89 : _GEN_11084; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11086 = 8'h4e == io_state_in_11 ? 8'h94 : _GEN_11085; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11087 = 8'h4f == io_state_in_11 ? 8'h9f : _GEN_11086; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11088 = 8'h50 == io_state_in_11 ? 8'h46 : _GEN_11087; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11089 = 8'h51 == io_state_in_11 ? 8'h4d : _GEN_11088; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11090 = 8'h52 == io_state_in_11 ? 8'h50 : _GEN_11089; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11091 = 8'h53 == io_state_in_11 ? 8'h5b : _GEN_11090; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11092 = 8'h54 == io_state_in_11 ? 8'h6a : _GEN_11091; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11093 = 8'h55 == io_state_in_11 ? 8'h61 : _GEN_11092; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11094 = 8'h56 == io_state_in_11 ? 8'h7c : _GEN_11093; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11095 = 8'h57 == io_state_in_11 ? 8'h77 : _GEN_11094; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11096 = 8'h58 == io_state_in_11 ? 8'h1e : _GEN_11095; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11097 = 8'h59 == io_state_in_11 ? 8'h15 : _GEN_11096; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11098 = 8'h5a == io_state_in_11 ? 8'h8 : _GEN_11097; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11099 = 8'h5b == io_state_in_11 ? 8'h3 : _GEN_11098; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11100 = 8'h5c == io_state_in_11 ? 8'h32 : _GEN_11099; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11101 = 8'h5d == io_state_in_11 ? 8'h39 : _GEN_11100; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11102 = 8'h5e == io_state_in_11 ? 8'h24 : _GEN_11101; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11103 = 8'h5f == io_state_in_11 ? 8'h2f : _GEN_11102; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11104 = 8'h60 == io_state_in_11 ? 8'h8d : _GEN_11103; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11105 = 8'h61 == io_state_in_11 ? 8'h86 : _GEN_11104; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11106 = 8'h62 == io_state_in_11 ? 8'h9b : _GEN_11105; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11107 = 8'h63 == io_state_in_11 ? 8'h90 : _GEN_11106; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11108 = 8'h64 == io_state_in_11 ? 8'ha1 : _GEN_11107; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11109 = 8'h65 == io_state_in_11 ? 8'haa : _GEN_11108; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11110 = 8'h66 == io_state_in_11 ? 8'hb7 : _GEN_11109; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11111 = 8'h67 == io_state_in_11 ? 8'hbc : _GEN_11110; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11112 = 8'h68 == io_state_in_11 ? 8'hd5 : _GEN_11111; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11113 = 8'h69 == io_state_in_11 ? 8'hde : _GEN_11112; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11114 = 8'h6a == io_state_in_11 ? 8'hc3 : _GEN_11113; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11115 = 8'h6b == io_state_in_11 ? 8'hc8 : _GEN_11114; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11116 = 8'h6c == io_state_in_11 ? 8'hf9 : _GEN_11115; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11117 = 8'h6d == io_state_in_11 ? 8'hf2 : _GEN_11116; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11118 = 8'h6e == io_state_in_11 ? 8'hef : _GEN_11117; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11119 = 8'h6f == io_state_in_11 ? 8'he4 : _GEN_11118; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11120 = 8'h70 == io_state_in_11 ? 8'h3d : _GEN_11119; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11121 = 8'h71 == io_state_in_11 ? 8'h36 : _GEN_11120; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11122 = 8'h72 == io_state_in_11 ? 8'h2b : _GEN_11121; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11123 = 8'h73 == io_state_in_11 ? 8'h20 : _GEN_11122; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11124 = 8'h74 == io_state_in_11 ? 8'h11 : _GEN_11123; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11125 = 8'h75 == io_state_in_11 ? 8'h1a : _GEN_11124; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11126 = 8'h76 == io_state_in_11 ? 8'h7 : _GEN_11125; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11127 = 8'h77 == io_state_in_11 ? 8'hc : _GEN_11126; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11128 = 8'h78 == io_state_in_11 ? 8'h65 : _GEN_11127; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11129 = 8'h79 == io_state_in_11 ? 8'h6e : _GEN_11128; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11130 = 8'h7a == io_state_in_11 ? 8'h73 : _GEN_11129; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11131 = 8'h7b == io_state_in_11 ? 8'h78 : _GEN_11130; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11132 = 8'h7c == io_state_in_11 ? 8'h49 : _GEN_11131; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11133 = 8'h7d == io_state_in_11 ? 8'h42 : _GEN_11132; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11134 = 8'h7e == io_state_in_11 ? 8'h5f : _GEN_11133; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11135 = 8'h7f == io_state_in_11 ? 8'h54 : _GEN_11134; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11136 = 8'h80 == io_state_in_11 ? 8'hf7 : _GEN_11135; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11137 = 8'h81 == io_state_in_11 ? 8'hfc : _GEN_11136; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11138 = 8'h82 == io_state_in_11 ? 8'he1 : _GEN_11137; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11139 = 8'h83 == io_state_in_11 ? 8'hea : _GEN_11138; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11140 = 8'h84 == io_state_in_11 ? 8'hdb : _GEN_11139; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11141 = 8'h85 == io_state_in_11 ? 8'hd0 : _GEN_11140; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11142 = 8'h86 == io_state_in_11 ? 8'hcd : _GEN_11141; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11143 = 8'h87 == io_state_in_11 ? 8'hc6 : _GEN_11142; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11144 = 8'h88 == io_state_in_11 ? 8'haf : _GEN_11143; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11145 = 8'h89 == io_state_in_11 ? 8'ha4 : _GEN_11144; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11146 = 8'h8a == io_state_in_11 ? 8'hb9 : _GEN_11145; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11147 = 8'h8b == io_state_in_11 ? 8'hb2 : _GEN_11146; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11148 = 8'h8c == io_state_in_11 ? 8'h83 : _GEN_11147; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11149 = 8'h8d == io_state_in_11 ? 8'h88 : _GEN_11148; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11150 = 8'h8e == io_state_in_11 ? 8'h95 : _GEN_11149; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11151 = 8'h8f == io_state_in_11 ? 8'h9e : _GEN_11150; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11152 = 8'h90 == io_state_in_11 ? 8'h47 : _GEN_11151; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11153 = 8'h91 == io_state_in_11 ? 8'h4c : _GEN_11152; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11154 = 8'h92 == io_state_in_11 ? 8'h51 : _GEN_11153; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11155 = 8'h93 == io_state_in_11 ? 8'h5a : _GEN_11154; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11156 = 8'h94 == io_state_in_11 ? 8'h6b : _GEN_11155; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11157 = 8'h95 == io_state_in_11 ? 8'h60 : _GEN_11156; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11158 = 8'h96 == io_state_in_11 ? 8'h7d : _GEN_11157; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11159 = 8'h97 == io_state_in_11 ? 8'h76 : _GEN_11158; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11160 = 8'h98 == io_state_in_11 ? 8'h1f : _GEN_11159; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11161 = 8'h99 == io_state_in_11 ? 8'h14 : _GEN_11160; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11162 = 8'h9a == io_state_in_11 ? 8'h9 : _GEN_11161; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11163 = 8'h9b == io_state_in_11 ? 8'h2 : _GEN_11162; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11164 = 8'h9c == io_state_in_11 ? 8'h33 : _GEN_11163; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11165 = 8'h9d == io_state_in_11 ? 8'h38 : _GEN_11164; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11166 = 8'h9e == io_state_in_11 ? 8'h25 : _GEN_11165; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11167 = 8'h9f == io_state_in_11 ? 8'h2e : _GEN_11166; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11168 = 8'ha0 == io_state_in_11 ? 8'h8c : _GEN_11167; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11169 = 8'ha1 == io_state_in_11 ? 8'h87 : _GEN_11168; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11170 = 8'ha2 == io_state_in_11 ? 8'h9a : _GEN_11169; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11171 = 8'ha3 == io_state_in_11 ? 8'h91 : _GEN_11170; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11172 = 8'ha4 == io_state_in_11 ? 8'ha0 : _GEN_11171; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11173 = 8'ha5 == io_state_in_11 ? 8'hab : _GEN_11172; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11174 = 8'ha6 == io_state_in_11 ? 8'hb6 : _GEN_11173; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11175 = 8'ha7 == io_state_in_11 ? 8'hbd : _GEN_11174; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11176 = 8'ha8 == io_state_in_11 ? 8'hd4 : _GEN_11175; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11177 = 8'ha9 == io_state_in_11 ? 8'hdf : _GEN_11176; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11178 = 8'haa == io_state_in_11 ? 8'hc2 : _GEN_11177; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11179 = 8'hab == io_state_in_11 ? 8'hc9 : _GEN_11178; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11180 = 8'hac == io_state_in_11 ? 8'hf8 : _GEN_11179; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11181 = 8'had == io_state_in_11 ? 8'hf3 : _GEN_11180; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11182 = 8'hae == io_state_in_11 ? 8'hee : _GEN_11181; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11183 = 8'haf == io_state_in_11 ? 8'he5 : _GEN_11182; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11184 = 8'hb0 == io_state_in_11 ? 8'h3c : _GEN_11183; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11185 = 8'hb1 == io_state_in_11 ? 8'h37 : _GEN_11184; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11186 = 8'hb2 == io_state_in_11 ? 8'h2a : _GEN_11185; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11187 = 8'hb3 == io_state_in_11 ? 8'h21 : _GEN_11186; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11188 = 8'hb4 == io_state_in_11 ? 8'h10 : _GEN_11187; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11189 = 8'hb5 == io_state_in_11 ? 8'h1b : _GEN_11188; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11190 = 8'hb6 == io_state_in_11 ? 8'h6 : _GEN_11189; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11191 = 8'hb7 == io_state_in_11 ? 8'hd : _GEN_11190; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11192 = 8'hb8 == io_state_in_11 ? 8'h64 : _GEN_11191; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11193 = 8'hb9 == io_state_in_11 ? 8'h6f : _GEN_11192; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11194 = 8'hba == io_state_in_11 ? 8'h72 : _GEN_11193; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11195 = 8'hbb == io_state_in_11 ? 8'h79 : _GEN_11194; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11196 = 8'hbc == io_state_in_11 ? 8'h48 : _GEN_11195; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11197 = 8'hbd == io_state_in_11 ? 8'h43 : _GEN_11196; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11198 = 8'hbe == io_state_in_11 ? 8'h5e : _GEN_11197; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11199 = 8'hbf == io_state_in_11 ? 8'h55 : _GEN_11198; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11200 = 8'hc0 == io_state_in_11 ? 8'h1 : _GEN_11199; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11201 = 8'hc1 == io_state_in_11 ? 8'ha : _GEN_11200; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11202 = 8'hc2 == io_state_in_11 ? 8'h17 : _GEN_11201; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11203 = 8'hc3 == io_state_in_11 ? 8'h1c : _GEN_11202; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11204 = 8'hc4 == io_state_in_11 ? 8'h2d : _GEN_11203; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11205 = 8'hc5 == io_state_in_11 ? 8'h26 : _GEN_11204; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11206 = 8'hc6 == io_state_in_11 ? 8'h3b : _GEN_11205; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11207 = 8'hc7 == io_state_in_11 ? 8'h30 : _GEN_11206; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11208 = 8'hc8 == io_state_in_11 ? 8'h59 : _GEN_11207; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11209 = 8'hc9 == io_state_in_11 ? 8'h52 : _GEN_11208; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11210 = 8'hca == io_state_in_11 ? 8'h4f : _GEN_11209; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11211 = 8'hcb == io_state_in_11 ? 8'h44 : _GEN_11210; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11212 = 8'hcc == io_state_in_11 ? 8'h75 : _GEN_11211; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11213 = 8'hcd == io_state_in_11 ? 8'h7e : _GEN_11212; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11214 = 8'hce == io_state_in_11 ? 8'h63 : _GEN_11213; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11215 = 8'hcf == io_state_in_11 ? 8'h68 : _GEN_11214; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11216 = 8'hd0 == io_state_in_11 ? 8'hb1 : _GEN_11215; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11217 = 8'hd1 == io_state_in_11 ? 8'hba : _GEN_11216; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11218 = 8'hd2 == io_state_in_11 ? 8'ha7 : _GEN_11217; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11219 = 8'hd3 == io_state_in_11 ? 8'hac : _GEN_11218; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11220 = 8'hd4 == io_state_in_11 ? 8'h9d : _GEN_11219; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11221 = 8'hd5 == io_state_in_11 ? 8'h96 : _GEN_11220; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11222 = 8'hd6 == io_state_in_11 ? 8'h8b : _GEN_11221; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11223 = 8'hd7 == io_state_in_11 ? 8'h80 : _GEN_11222; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11224 = 8'hd8 == io_state_in_11 ? 8'he9 : _GEN_11223; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11225 = 8'hd9 == io_state_in_11 ? 8'he2 : _GEN_11224; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11226 = 8'hda == io_state_in_11 ? 8'hff : _GEN_11225; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11227 = 8'hdb == io_state_in_11 ? 8'hf4 : _GEN_11226; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11228 = 8'hdc == io_state_in_11 ? 8'hc5 : _GEN_11227; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11229 = 8'hdd == io_state_in_11 ? 8'hce : _GEN_11228; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11230 = 8'hde == io_state_in_11 ? 8'hd3 : _GEN_11229; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11231 = 8'hdf == io_state_in_11 ? 8'hd8 : _GEN_11230; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11232 = 8'he0 == io_state_in_11 ? 8'h7a : _GEN_11231; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11233 = 8'he1 == io_state_in_11 ? 8'h71 : _GEN_11232; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11234 = 8'he2 == io_state_in_11 ? 8'h6c : _GEN_11233; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11235 = 8'he3 == io_state_in_11 ? 8'h67 : _GEN_11234; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11236 = 8'he4 == io_state_in_11 ? 8'h56 : _GEN_11235; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11237 = 8'he5 == io_state_in_11 ? 8'h5d : _GEN_11236; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11238 = 8'he6 == io_state_in_11 ? 8'h40 : _GEN_11237; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11239 = 8'he7 == io_state_in_11 ? 8'h4b : _GEN_11238; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11240 = 8'he8 == io_state_in_11 ? 8'h22 : _GEN_11239; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11241 = 8'he9 == io_state_in_11 ? 8'h29 : _GEN_11240; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11242 = 8'hea == io_state_in_11 ? 8'h34 : _GEN_11241; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11243 = 8'heb == io_state_in_11 ? 8'h3f : _GEN_11242; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11244 = 8'hec == io_state_in_11 ? 8'he : _GEN_11243; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11245 = 8'hed == io_state_in_11 ? 8'h5 : _GEN_11244; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11246 = 8'hee == io_state_in_11 ? 8'h18 : _GEN_11245; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11247 = 8'hef == io_state_in_11 ? 8'h13 : _GEN_11246; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11248 = 8'hf0 == io_state_in_11 ? 8'hca : _GEN_11247; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11249 = 8'hf1 == io_state_in_11 ? 8'hc1 : _GEN_11248; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11250 = 8'hf2 == io_state_in_11 ? 8'hdc : _GEN_11249; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11251 = 8'hf3 == io_state_in_11 ? 8'hd7 : _GEN_11250; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11252 = 8'hf4 == io_state_in_11 ? 8'he6 : _GEN_11251; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11253 = 8'hf5 == io_state_in_11 ? 8'hed : _GEN_11252; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11254 = 8'hf6 == io_state_in_11 ? 8'hf0 : _GEN_11253; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11255 = 8'hf7 == io_state_in_11 ? 8'hfb : _GEN_11254; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11256 = 8'hf8 == io_state_in_11 ? 8'h92 : _GEN_11255; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11257 = 8'hf9 == io_state_in_11 ? 8'h99 : _GEN_11256; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11258 = 8'hfa == io_state_in_11 ? 8'h84 : _GEN_11257; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11259 = 8'hfb == io_state_in_11 ? 8'h8f : _GEN_11258; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11260 = 8'hfc == io_state_in_11 ? 8'hbe : _GEN_11259; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11261 = 8'hfd == io_state_in_11 ? 8'hb5 : _GEN_11260; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11262 = 8'hfe == io_state_in_11 ? 8'ha8 : _GEN_11261; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11263 = 8'hff == io_state_in_11 ? 8'ha3 : _GEN_11262; // @[InvMixColumns.scala 138:{91,91}]
  wire [7:0] _GEN_11265 = 8'h1 == io_state_in_8 ? 8'hb : 8'h0; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11266 = 8'h2 == io_state_in_8 ? 8'h16 : _GEN_11265; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11267 = 8'h3 == io_state_in_8 ? 8'h1d : _GEN_11266; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11268 = 8'h4 == io_state_in_8 ? 8'h2c : _GEN_11267; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11269 = 8'h5 == io_state_in_8 ? 8'h27 : _GEN_11268; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11270 = 8'h6 == io_state_in_8 ? 8'h3a : _GEN_11269; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11271 = 8'h7 == io_state_in_8 ? 8'h31 : _GEN_11270; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11272 = 8'h8 == io_state_in_8 ? 8'h58 : _GEN_11271; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11273 = 8'h9 == io_state_in_8 ? 8'h53 : _GEN_11272; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11274 = 8'ha == io_state_in_8 ? 8'h4e : _GEN_11273; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11275 = 8'hb == io_state_in_8 ? 8'h45 : _GEN_11274; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11276 = 8'hc == io_state_in_8 ? 8'h74 : _GEN_11275; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11277 = 8'hd == io_state_in_8 ? 8'h7f : _GEN_11276; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11278 = 8'he == io_state_in_8 ? 8'h62 : _GEN_11277; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11279 = 8'hf == io_state_in_8 ? 8'h69 : _GEN_11278; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11280 = 8'h10 == io_state_in_8 ? 8'hb0 : _GEN_11279; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11281 = 8'h11 == io_state_in_8 ? 8'hbb : _GEN_11280; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11282 = 8'h12 == io_state_in_8 ? 8'ha6 : _GEN_11281; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11283 = 8'h13 == io_state_in_8 ? 8'had : _GEN_11282; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11284 = 8'h14 == io_state_in_8 ? 8'h9c : _GEN_11283; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11285 = 8'h15 == io_state_in_8 ? 8'h97 : _GEN_11284; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11286 = 8'h16 == io_state_in_8 ? 8'h8a : _GEN_11285; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11287 = 8'h17 == io_state_in_8 ? 8'h81 : _GEN_11286; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11288 = 8'h18 == io_state_in_8 ? 8'he8 : _GEN_11287; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11289 = 8'h19 == io_state_in_8 ? 8'he3 : _GEN_11288; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11290 = 8'h1a == io_state_in_8 ? 8'hfe : _GEN_11289; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11291 = 8'h1b == io_state_in_8 ? 8'hf5 : _GEN_11290; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11292 = 8'h1c == io_state_in_8 ? 8'hc4 : _GEN_11291; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11293 = 8'h1d == io_state_in_8 ? 8'hcf : _GEN_11292; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11294 = 8'h1e == io_state_in_8 ? 8'hd2 : _GEN_11293; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11295 = 8'h1f == io_state_in_8 ? 8'hd9 : _GEN_11294; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11296 = 8'h20 == io_state_in_8 ? 8'h7b : _GEN_11295; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11297 = 8'h21 == io_state_in_8 ? 8'h70 : _GEN_11296; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11298 = 8'h22 == io_state_in_8 ? 8'h6d : _GEN_11297; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11299 = 8'h23 == io_state_in_8 ? 8'h66 : _GEN_11298; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11300 = 8'h24 == io_state_in_8 ? 8'h57 : _GEN_11299; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11301 = 8'h25 == io_state_in_8 ? 8'h5c : _GEN_11300; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11302 = 8'h26 == io_state_in_8 ? 8'h41 : _GEN_11301; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11303 = 8'h27 == io_state_in_8 ? 8'h4a : _GEN_11302; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11304 = 8'h28 == io_state_in_8 ? 8'h23 : _GEN_11303; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11305 = 8'h29 == io_state_in_8 ? 8'h28 : _GEN_11304; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11306 = 8'h2a == io_state_in_8 ? 8'h35 : _GEN_11305; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11307 = 8'h2b == io_state_in_8 ? 8'h3e : _GEN_11306; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11308 = 8'h2c == io_state_in_8 ? 8'hf : _GEN_11307; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11309 = 8'h2d == io_state_in_8 ? 8'h4 : _GEN_11308; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11310 = 8'h2e == io_state_in_8 ? 8'h19 : _GEN_11309; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11311 = 8'h2f == io_state_in_8 ? 8'h12 : _GEN_11310; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11312 = 8'h30 == io_state_in_8 ? 8'hcb : _GEN_11311; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11313 = 8'h31 == io_state_in_8 ? 8'hc0 : _GEN_11312; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11314 = 8'h32 == io_state_in_8 ? 8'hdd : _GEN_11313; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11315 = 8'h33 == io_state_in_8 ? 8'hd6 : _GEN_11314; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11316 = 8'h34 == io_state_in_8 ? 8'he7 : _GEN_11315; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11317 = 8'h35 == io_state_in_8 ? 8'hec : _GEN_11316; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11318 = 8'h36 == io_state_in_8 ? 8'hf1 : _GEN_11317; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11319 = 8'h37 == io_state_in_8 ? 8'hfa : _GEN_11318; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11320 = 8'h38 == io_state_in_8 ? 8'h93 : _GEN_11319; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11321 = 8'h39 == io_state_in_8 ? 8'h98 : _GEN_11320; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11322 = 8'h3a == io_state_in_8 ? 8'h85 : _GEN_11321; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11323 = 8'h3b == io_state_in_8 ? 8'h8e : _GEN_11322; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11324 = 8'h3c == io_state_in_8 ? 8'hbf : _GEN_11323; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11325 = 8'h3d == io_state_in_8 ? 8'hb4 : _GEN_11324; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11326 = 8'h3e == io_state_in_8 ? 8'ha9 : _GEN_11325; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11327 = 8'h3f == io_state_in_8 ? 8'ha2 : _GEN_11326; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11328 = 8'h40 == io_state_in_8 ? 8'hf6 : _GEN_11327; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11329 = 8'h41 == io_state_in_8 ? 8'hfd : _GEN_11328; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11330 = 8'h42 == io_state_in_8 ? 8'he0 : _GEN_11329; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11331 = 8'h43 == io_state_in_8 ? 8'heb : _GEN_11330; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11332 = 8'h44 == io_state_in_8 ? 8'hda : _GEN_11331; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11333 = 8'h45 == io_state_in_8 ? 8'hd1 : _GEN_11332; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11334 = 8'h46 == io_state_in_8 ? 8'hcc : _GEN_11333; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11335 = 8'h47 == io_state_in_8 ? 8'hc7 : _GEN_11334; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11336 = 8'h48 == io_state_in_8 ? 8'hae : _GEN_11335; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11337 = 8'h49 == io_state_in_8 ? 8'ha5 : _GEN_11336; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11338 = 8'h4a == io_state_in_8 ? 8'hb8 : _GEN_11337; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11339 = 8'h4b == io_state_in_8 ? 8'hb3 : _GEN_11338; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11340 = 8'h4c == io_state_in_8 ? 8'h82 : _GEN_11339; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11341 = 8'h4d == io_state_in_8 ? 8'h89 : _GEN_11340; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11342 = 8'h4e == io_state_in_8 ? 8'h94 : _GEN_11341; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11343 = 8'h4f == io_state_in_8 ? 8'h9f : _GEN_11342; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11344 = 8'h50 == io_state_in_8 ? 8'h46 : _GEN_11343; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11345 = 8'h51 == io_state_in_8 ? 8'h4d : _GEN_11344; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11346 = 8'h52 == io_state_in_8 ? 8'h50 : _GEN_11345; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11347 = 8'h53 == io_state_in_8 ? 8'h5b : _GEN_11346; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11348 = 8'h54 == io_state_in_8 ? 8'h6a : _GEN_11347; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11349 = 8'h55 == io_state_in_8 ? 8'h61 : _GEN_11348; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11350 = 8'h56 == io_state_in_8 ? 8'h7c : _GEN_11349; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11351 = 8'h57 == io_state_in_8 ? 8'h77 : _GEN_11350; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11352 = 8'h58 == io_state_in_8 ? 8'h1e : _GEN_11351; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11353 = 8'h59 == io_state_in_8 ? 8'h15 : _GEN_11352; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11354 = 8'h5a == io_state_in_8 ? 8'h8 : _GEN_11353; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11355 = 8'h5b == io_state_in_8 ? 8'h3 : _GEN_11354; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11356 = 8'h5c == io_state_in_8 ? 8'h32 : _GEN_11355; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11357 = 8'h5d == io_state_in_8 ? 8'h39 : _GEN_11356; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11358 = 8'h5e == io_state_in_8 ? 8'h24 : _GEN_11357; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11359 = 8'h5f == io_state_in_8 ? 8'h2f : _GEN_11358; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11360 = 8'h60 == io_state_in_8 ? 8'h8d : _GEN_11359; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11361 = 8'h61 == io_state_in_8 ? 8'h86 : _GEN_11360; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11362 = 8'h62 == io_state_in_8 ? 8'h9b : _GEN_11361; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11363 = 8'h63 == io_state_in_8 ? 8'h90 : _GEN_11362; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11364 = 8'h64 == io_state_in_8 ? 8'ha1 : _GEN_11363; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11365 = 8'h65 == io_state_in_8 ? 8'haa : _GEN_11364; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11366 = 8'h66 == io_state_in_8 ? 8'hb7 : _GEN_11365; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11367 = 8'h67 == io_state_in_8 ? 8'hbc : _GEN_11366; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11368 = 8'h68 == io_state_in_8 ? 8'hd5 : _GEN_11367; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11369 = 8'h69 == io_state_in_8 ? 8'hde : _GEN_11368; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11370 = 8'h6a == io_state_in_8 ? 8'hc3 : _GEN_11369; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11371 = 8'h6b == io_state_in_8 ? 8'hc8 : _GEN_11370; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11372 = 8'h6c == io_state_in_8 ? 8'hf9 : _GEN_11371; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11373 = 8'h6d == io_state_in_8 ? 8'hf2 : _GEN_11372; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11374 = 8'h6e == io_state_in_8 ? 8'hef : _GEN_11373; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11375 = 8'h6f == io_state_in_8 ? 8'he4 : _GEN_11374; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11376 = 8'h70 == io_state_in_8 ? 8'h3d : _GEN_11375; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11377 = 8'h71 == io_state_in_8 ? 8'h36 : _GEN_11376; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11378 = 8'h72 == io_state_in_8 ? 8'h2b : _GEN_11377; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11379 = 8'h73 == io_state_in_8 ? 8'h20 : _GEN_11378; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11380 = 8'h74 == io_state_in_8 ? 8'h11 : _GEN_11379; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11381 = 8'h75 == io_state_in_8 ? 8'h1a : _GEN_11380; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11382 = 8'h76 == io_state_in_8 ? 8'h7 : _GEN_11381; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11383 = 8'h77 == io_state_in_8 ? 8'hc : _GEN_11382; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11384 = 8'h78 == io_state_in_8 ? 8'h65 : _GEN_11383; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11385 = 8'h79 == io_state_in_8 ? 8'h6e : _GEN_11384; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11386 = 8'h7a == io_state_in_8 ? 8'h73 : _GEN_11385; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11387 = 8'h7b == io_state_in_8 ? 8'h78 : _GEN_11386; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11388 = 8'h7c == io_state_in_8 ? 8'h49 : _GEN_11387; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11389 = 8'h7d == io_state_in_8 ? 8'h42 : _GEN_11388; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11390 = 8'h7e == io_state_in_8 ? 8'h5f : _GEN_11389; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11391 = 8'h7f == io_state_in_8 ? 8'h54 : _GEN_11390; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11392 = 8'h80 == io_state_in_8 ? 8'hf7 : _GEN_11391; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11393 = 8'h81 == io_state_in_8 ? 8'hfc : _GEN_11392; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11394 = 8'h82 == io_state_in_8 ? 8'he1 : _GEN_11393; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11395 = 8'h83 == io_state_in_8 ? 8'hea : _GEN_11394; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11396 = 8'h84 == io_state_in_8 ? 8'hdb : _GEN_11395; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11397 = 8'h85 == io_state_in_8 ? 8'hd0 : _GEN_11396; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11398 = 8'h86 == io_state_in_8 ? 8'hcd : _GEN_11397; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11399 = 8'h87 == io_state_in_8 ? 8'hc6 : _GEN_11398; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11400 = 8'h88 == io_state_in_8 ? 8'haf : _GEN_11399; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11401 = 8'h89 == io_state_in_8 ? 8'ha4 : _GEN_11400; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11402 = 8'h8a == io_state_in_8 ? 8'hb9 : _GEN_11401; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11403 = 8'h8b == io_state_in_8 ? 8'hb2 : _GEN_11402; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11404 = 8'h8c == io_state_in_8 ? 8'h83 : _GEN_11403; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11405 = 8'h8d == io_state_in_8 ? 8'h88 : _GEN_11404; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11406 = 8'h8e == io_state_in_8 ? 8'h95 : _GEN_11405; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11407 = 8'h8f == io_state_in_8 ? 8'h9e : _GEN_11406; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11408 = 8'h90 == io_state_in_8 ? 8'h47 : _GEN_11407; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11409 = 8'h91 == io_state_in_8 ? 8'h4c : _GEN_11408; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11410 = 8'h92 == io_state_in_8 ? 8'h51 : _GEN_11409; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11411 = 8'h93 == io_state_in_8 ? 8'h5a : _GEN_11410; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11412 = 8'h94 == io_state_in_8 ? 8'h6b : _GEN_11411; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11413 = 8'h95 == io_state_in_8 ? 8'h60 : _GEN_11412; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11414 = 8'h96 == io_state_in_8 ? 8'h7d : _GEN_11413; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11415 = 8'h97 == io_state_in_8 ? 8'h76 : _GEN_11414; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11416 = 8'h98 == io_state_in_8 ? 8'h1f : _GEN_11415; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11417 = 8'h99 == io_state_in_8 ? 8'h14 : _GEN_11416; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11418 = 8'h9a == io_state_in_8 ? 8'h9 : _GEN_11417; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11419 = 8'h9b == io_state_in_8 ? 8'h2 : _GEN_11418; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11420 = 8'h9c == io_state_in_8 ? 8'h33 : _GEN_11419; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11421 = 8'h9d == io_state_in_8 ? 8'h38 : _GEN_11420; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11422 = 8'h9e == io_state_in_8 ? 8'h25 : _GEN_11421; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11423 = 8'h9f == io_state_in_8 ? 8'h2e : _GEN_11422; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11424 = 8'ha0 == io_state_in_8 ? 8'h8c : _GEN_11423; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11425 = 8'ha1 == io_state_in_8 ? 8'h87 : _GEN_11424; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11426 = 8'ha2 == io_state_in_8 ? 8'h9a : _GEN_11425; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11427 = 8'ha3 == io_state_in_8 ? 8'h91 : _GEN_11426; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11428 = 8'ha4 == io_state_in_8 ? 8'ha0 : _GEN_11427; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11429 = 8'ha5 == io_state_in_8 ? 8'hab : _GEN_11428; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11430 = 8'ha6 == io_state_in_8 ? 8'hb6 : _GEN_11429; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11431 = 8'ha7 == io_state_in_8 ? 8'hbd : _GEN_11430; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11432 = 8'ha8 == io_state_in_8 ? 8'hd4 : _GEN_11431; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11433 = 8'ha9 == io_state_in_8 ? 8'hdf : _GEN_11432; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11434 = 8'haa == io_state_in_8 ? 8'hc2 : _GEN_11433; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11435 = 8'hab == io_state_in_8 ? 8'hc9 : _GEN_11434; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11436 = 8'hac == io_state_in_8 ? 8'hf8 : _GEN_11435; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11437 = 8'had == io_state_in_8 ? 8'hf3 : _GEN_11436; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11438 = 8'hae == io_state_in_8 ? 8'hee : _GEN_11437; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11439 = 8'haf == io_state_in_8 ? 8'he5 : _GEN_11438; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11440 = 8'hb0 == io_state_in_8 ? 8'h3c : _GEN_11439; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11441 = 8'hb1 == io_state_in_8 ? 8'h37 : _GEN_11440; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11442 = 8'hb2 == io_state_in_8 ? 8'h2a : _GEN_11441; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11443 = 8'hb3 == io_state_in_8 ? 8'h21 : _GEN_11442; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11444 = 8'hb4 == io_state_in_8 ? 8'h10 : _GEN_11443; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11445 = 8'hb5 == io_state_in_8 ? 8'h1b : _GEN_11444; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11446 = 8'hb6 == io_state_in_8 ? 8'h6 : _GEN_11445; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11447 = 8'hb7 == io_state_in_8 ? 8'hd : _GEN_11446; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11448 = 8'hb8 == io_state_in_8 ? 8'h64 : _GEN_11447; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11449 = 8'hb9 == io_state_in_8 ? 8'h6f : _GEN_11448; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11450 = 8'hba == io_state_in_8 ? 8'h72 : _GEN_11449; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11451 = 8'hbb == io_state_in_8 ? 8'h79 : _GEN_11450; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11452 = 8'hbc == io_state_in_8 ? 8'h48 : _GEN_11451; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11453 = 8'hbd == io_state_in_8 ? 8'h43 : _GEN_11452; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11454 = 8'hbe == io_state_in_8 ? 8'h5e : _GEN_11453; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11455 = 8'hbf == io_state_in_8 ? 8'h55 : _GEN_11454; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11456 = 8'hc0 == io_state_in_8 ? 8'h1 : _GEN_11455; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11457 = 8'hc1 == io_state_in_8 ? 8'ha : _GEN_11456; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11458 = 8'hc2 == io_state_in_8 ? 8'h17 : _GEN_11457; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11459 = 8'hc3 == io_state_in_8 ? 8'h1c : _GEN_11458; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11460 = 8'hc4 == io_state_in_8 ? 8'h2d : _GEN_11459; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11461 = 8'hc5 == io_state_in_8 ? 8'h26 : _GEN_11460; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11462 = 8'hc6 == io_state_in_8 ? 8'h3b : _GEN_11461; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11463 = 8'hc7 == io_state_in_8 ? 8'h30 : _GEN_11462; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11464 = 8'hc8 == io_state_in_8 ? 8'h59 : _GEN_11463; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11465 = 8'hc9 == io_state_in_8 ? 8'h52 : _GEN_11464; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11466 = 8'hca == io_state_in_8 ? 8'h4f : _GEN_11465; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11467 = 8'hcb == io_state_in_8 ? 8'h44 : _GEN_11466; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11468 = 8'hcc == io_state_in_8 ? 8'h75 : _GEN_11467; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11469 = 8'hcd == io_state_in_8 ? 8'h7e : _GEN_11468; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11470 = 8'hce == io_state_in_8 ? 8'h63 : _GEN_11469; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11471 = 8'hcf == io_state_in_8 ? 8'h68 : _GEN_11470; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11472 = 8'hd0 == io_state_in_8 ? 8'hb1 : _GEN_11471; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11473 = 8'hd1 == io_state_in_8 ? 8'hba : _GEN_11472; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11474 = 8'hd2 == io_state_in_8 ? 8'ha7 : _GEN_11473; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11475 = 8'hd3 == io_state_in_8 ? 8'hac : _GEN_11474; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11476 = 8'hd4 == io_state_in_8 ? 8'h9d : _GEN_11475; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11477 = 8'hd5 == io_state_in_8 ? 8'h96 : _GEN_11476; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11478 = 8'hd6 == io_state_in_8 ? 8'h8b : _GEN_11477; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11479 = 8'hd7 == io_state_in_8 ? 8'h80 : _GEN_11478; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11480 = 8'hd8 == io_state_in_8 ? 8'he9 : _GEN_11479; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11481 = 8'hd9 == io_state_in_8 ? 8'he2 : _GEN_11480; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11482 = 8'hda == io_state_in_8 ? 8'hff : _GEN_11481; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11483 = 8'hdb == io_state_in_8 ? 8'hf4 : _GEN_11482; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11484 = 8'hdc == io_state_in_8 ? 8'hc5 : _GEN_11483; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11485 = 8'hdd == io_state_in_8 ? 8'hce : _GEN_11484; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11486 = 8'hde == io_state_in_8 ? 8'hd3 : _GEN_11485; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11487 = 8'hdf == io_state_in_8 ? 8'hd8 : _GEN_11486; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11488 = 8'he0 == io_state_in_8 ? 8'h7a : _GEN_11487; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11489 = 8'he1 == io_state_in_8 ? 8'h71 : _GEN_11488; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11490 = 8'he2 == io_state_in_8 ? 8'h6c : _GEN_11489; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11491 = 8'he3 == io_state_in_8 ? 8'h67 : _GEN_11490; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11492 = 8'he4 == io_state_in_8 ? 8'h56 : _GEN_11491; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11493 = 8'he5 == io_state_in_8 ? 8'h5d : _GEN_11492; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11494 = 8'he6 == io_state_in_8 ? 8'h40 : _GEN_11493; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11495 = 8'he7 == io_state_in_8 ? 8'h4b : _GEN_11494; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11496 = 8'he8 == io_state_in_8 ? 8'h22 : _GEN_11495; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11497 = 8'he9 == io_state_in_8 ? 8'h29 : _GEN_11496; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11498 = 8'hea == io_state_in_8 ? 8'h34 : _GEN_11497; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11499 = 8'heb == io_state_in_8 ? 8'h3f : _GEN_11498; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11500 = 8'hec == io_state_in_8 ? 8'he : _GEN_11499; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11501 = 8'hed == io_state_in_8 ? 8'h5 : _GEN_11500; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11502 = 8'hee == io_state_in_8 ? 8'h18 : _GEN_11501; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11503 = 8'hef == io_state_in_8 ? 8'h13 : _GEN_11502; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11504 = 8'hf0 == io_state_in_8 ? 8'hca : _GEN_11503; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11505 = 8'hf1 == io_state_in_8 ? 8'hc1 : _GEN_11504; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11506 = 8'hf2 == io_state_in_8 ? 8'hdc : _GEN_11505; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11507 = 8'hf3 == io_state_in_8 ? 8'hd7 : _GEN_11506; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11508 = 8'hf4 == io_state_in_8 ? 8'he6 : _GEN_11507; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11509 = 8'hf5 == io_state_in_8 ? 8'hed : _GEN_11508; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11510 = 8'hf6 == io_state_in_8 ? 8'hf0 : _GEN_11509; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11511 = 8'hf7 == io_state_in_8 ? 8'hfb : _GEN_11510; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11512 = 8'hf8 == io_state_in_8 ? 8'h92 : _GEN_11511; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11513 = 8'hf9 == io_state_in_8 ? 8'h99 : _GEN_11512; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11514 = 8'hfa == io_state_in_8 ? 8'h84 : _GEN_11513; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11515 = 8'hfb == io_state_in_8 ? 8'h8f : _GEN_11514; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11516 = 8'hfc == io_state_in_8 ? 8'hbe : _GEN_11515; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11517 = 8'hfd == io_state_in_8 ? 8'hb5 : _GEN_11516; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11518 = 8'hfe == io_state_in_8 ? 8'ha8 : _GEN_11517; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11519 = 8'hff == io_state_in_8 ? 8'ha3 : _GEN_11518; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11521 = 8'h1 == io_state_in_9 ? 8'hd : 8'h0; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11522 = 8'h2 == io_state_in_9 ? 8'h1a : _GEN_11521; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11523 = 8'h3 == io_state_in_9 ? 8'h17 : _GEN_11522; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11524 = 8'h4 == io_state_in_9 ? 8'h34 : _GEN_11523; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11525 = 8'h5 == io_state_in_9 ? 8'h39 : _GEN_11524; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11526 = 8'h6 == io_state_in_9 ? 8'h2e : _GEN_11525; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11527 = 8'h7 == io_state_in_9 ? 8'h23 : _GEN_11526; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11528 = 8'h8 == io_state_in_9 ? 8'h68 : _GEN_11527; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11529 = 8'h9 == io_state_in_9 ? 8'h65 : _GEN_11528; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11530 = 8'ha == io_state_in_9 ? 8'h72 : _GEN_11529; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11531 = 8'hb == io_state_in_9 ? 8'h7f : _GEN_11530; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11532 = 8'hc == io_state_in_9 ? 8'h5c : _GEN_11531; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11533 = 8'hd == io_state_in_9 ? 8'h51 : _GEN_11532; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11534 = 8'he == io_state_in_9 ? 8'h46 : _GEN_11533; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11535 = 8'hf == io_state_in_9 ? 8'h4b : _GEN_11534; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11536 = 8'h10 == io_state_in_9 ? 8'hd0 : _GEN_11535; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11537 = 8'h11 == io_state_in_9 ? 8'hdd : _GEN_11536; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11538 = 8'h12 == io_state_in_9 ? 8'hca : _GEN_11537; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11539 = 8'h13 == io_state_in_9 ? 8'hc7 : _GEN_11538; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11540 = 8'h14 == io_state_in_9 ? 8'he4 : _GEN_11539; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11541 = 8'h15 == io_state_in_9 ? 8'he9 : _GEN_11540; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11542 = 8'h16 == io_state_in_9 ? 8'hfe : _GEN_11541; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11543 = 8'h17 == io_state_in_9 ? 8'hf3 : _GEN_11542; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11544 = 8'h18 == io_state_in_9 ? 8'hb8 : _GEN_11543; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11545 = 8'h19 == io_state_in_9 ? 8'hb5 : _GEN_11544; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11546 = 8'h1a == io_state_in_9 ? 8'ha2 : _GEN_11545; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11547 = 8'h1b == io_state_in_9 ? 8'haf : _GEN_11546; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11548 = 8'h1c == io_state_in_9 ? 8'h8c : _GEN_11547; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11549 = 8'h1d == io_state_in_9 ? 8'h81 : _GEN_11548; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11550 = 8'h1e == io_state_in_9 ? 8'h96 : _GEN_11549; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11551 = 8'h1f == io_state_in_9 ? 8'h9b : _GEN_11550; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11552 = 8'h20 == io_state_in_9 ? 8'hbb : _GEN_11551; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11553 = 8'h21 == io_state_in_9 ? 8'hb6 : _GEN_11552; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11554 = 8'h22 == io_state_in_9 ? 8'ha1 : _GEN_11553; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11555 = 8'h23 == io_state_in_9 ? 8'hac : _GEN_11554; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11556 = 8'h24 == io_state_in_9 ? 8'h8f : _GEN_11555; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11557 = 8'h25 == io_state_in_9 ? 8'h82 : _GEN_11556; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11558 = 8'h26 == io_state_in_9 ? 8'h95 : _GEN_11557; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11559 = 8'h27 == io_state_in_9 ? 8'h98 : _GEN_11558; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11560 = 8'h28 == io_state_in_9 ? 8'hd3 : _GEN_11559; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11561 = 8'h29 == io_state_in_9 ? 8'hde : _GEN_11560; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11562 = 8'h2a == io_state_in_9 ? 8'hc9 : _GEN_11561; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11563 = 8'h2b == io_state_in_9 ? 8'hc4 : _GEN_11562; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11564 = 8'h2c == io_state_in_9 ? 8'he7 : _GEN_11563; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11565 = 8'h2d == io_state_in_9 ? 8'hea : _GEN_11564; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11566 = 8'h2e == io_state_in_9 ? 8'hfd : _GEN_11565; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11567 = 8'h2f == io_state_in_9 ? 8'hf0 : _GEN_11566; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11568 = 8'h30 == io_state_in_9 ? 8'h6b : _GEN_11567; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11569 = 8'h31 == io_state_in_9 ? 8'h66 : _GEN_11568; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11570 = 8'h32 == io_state_in_9 ? 8'h71 : _GEN_11569; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11571 = 8'h33 == io_state_in_9 ? 8'h7c : _GEN_11570; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11572 = 8'h34 == io_state_in_9 ? 8'h5f : _GEN_11571; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11573 = 8'h35 == io_state_in_9 ? 8'h52 : _GEN_11572; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11574 = 8'h36 == io_state_in_9 ? 8'h45 : _GEN_11573; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11575 = 8'h37 == io_state_in_9 ? 8'h48 : _GEN_11574; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11576 = 8'h38 == io_state_in_9 ? 8'h3 : _GEN_11575; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11577 = 8'h39 == io_state_in_9 ? 8'he : _GEN_11576; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11578 = 8'h3a == io_state_in_9 ? 8'h19 : _GEN_11577; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11579 = 8'h3b == io_state_in_9 ? 8'h14 : _GEN_11578; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11580 = 8'h3c == io_state_in_9 ? 8'h37 : _GEN_11579; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11581 = 8'h3d == io_state_in_9 ? 8'h3a : _GEN_11580; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11582 = 8'h3e == io_state_in_9 ? 8'h2d : _GEN_11581; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11583 = 8'h3f == io_state_in_9 ? 8'h20 : _GEN_11582; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11584 = 8'h40 == io_state_in_9 ? 8'h6d : _GEN_11583; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11585 = 8'h41 == io_state_in_9 ? 8'h60 : _GEN_11584; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11586 = 8'h42 == io_state_in_9 ? 8'h77 : _GEN_11585; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11587 = 8'h43 == io_state_in_9 ? 8'h7a : _GEN_11586; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11588 = 8'h44 == io_state_in_9 ? 8'h59 : _GEN_11587; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11589 = 8'h45 == io_state_in_9 ? 8'h54 : _GEN_11588; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11590 = 8'h46 == io_state_in_9 ? 8'h43 : _GEN_11589; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11591 = 8'h47 == io_state_in_9 ? 8'h4e : _GEN_11590; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11592 = 8'h48 == io_state_in_9 ? 8'h5 : _GEN_11591; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11593 = 8'h49 == io_state_in_9 ? 8'h8 : _GEN_11592; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11594 = 8'h4a == io_state_in_9 ? 8'h1f : _GEN_11593; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11595 = 8'h4b == io_state_in_9 ? 8'h12 : _GEN_11594; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11596 = 8'h4c == io_state_in_9 ? 8'h31 : _GEN_11595; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11597 = 8'h4d == io_state_in_9 ? 8'h3c : _GEN_11596; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11598 = 8'h4e == io_state_in_9 ? 8'h2b : _GEN_11597; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11599 = 8'h4f == io_state_in_9 ? 8'h26 : _GEN_11598; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11600 = 8'h50 == io_state_in_9 ? 8'hbd : _GEN_11599; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11601 = 8'h51 == io_state_in_9 ? 8'hb0 : _GEN_11600; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11602 = 8'h52 == io_state_in_9 ? 8'ha7 : _GEN_11601; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11603 = 8'h53 == io_state_in_9 ? 8'haa : _GEN_11602; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11604 = 8'h54 == io_state_in_9 ? 8'h89 : _GEN_11603; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11605 = 8'h55 == io_state_in_9 ? 8'h84 : _GEN_11604; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11606 = 8'h56 == io_state_in_9 ? 8'h93 : _GEN_11605; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11607 = 8'h57 == io_state_in_9 ? 8'h9e : _GEN_11606; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11608 = 8'h58 == io_state_in_9 ? 8'hd5 : _GEN_11607; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11609 = 8'h59 == io_state_in_9 ? 8'hd8 : _GEN_11608; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11610 = 8'h5a == io_state_in_9 ? 8'hcf : _GEN_11609; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11611 = 8'h5b == io_state_in_9 ? 8'hc2 : _GEN_11610; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11612 = 8'h5c == io_state_in_9 ? 8'he1 : _GEN_11611; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11613 = 8'h5d == io_state_in_9 ? 8'hec : _GEN_11612; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11614 = 8'h5e == io_state_in_9 ? 8'hfb : _GEN_11613; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11615 = 8'h5f == io_state_in_9 ? 8'hf6 : _GEN_11614; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11616 = 8'h60 == io_state_in_9 ? 8'hd6 : _GEN_11615; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11617 = 8'h61 == io_state_in_9 ? 8'hdb : _GEN_11616; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11618 = 8'h62 == io_state_in_9 ? 8'hcc : _GEN_11617; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11619 = 8'h63 == io_state_in_9 ? 8'hc1 : _GEN_11618; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11620 = 8'h64 == io_state_in_9 ? 8'he2 : _GEN_11619; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11621 = 8'h65 == io_state_in_9 ? 8'hef : _GEN_11620; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11622 = 8'h66 == io_state_in_9 ? 8'hf8 : _GEN_11621; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11623 = 8'h67 == io_state_in_9 ? 8'hf5 : _GEN_11622; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11624 = 8'h68 == io_state_in_9 ? 8'hbe : _GEN_11623; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11625 = 8'h69 == io_state_in_9 ? 8'hb3 : _GEN_11624; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11626 = 8'h6a == io_state_in_9 ? 8'ha4 : _GEN_11625; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11627 = 8'h6b == io_state_in_9 ? 8'ha9 : _GEN_11626; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11628 = 8'h6c == io_state_in_9 ? 8'h8a : _GEN_11627; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11629 = 8'h6d == io_state_in_9 ? 8'h87 : _GEN_11628; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11630 = 8'h6e == io_state_in_9 ? 8'h90 : _GEN_11629; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11631 = 8'h6f == io_state_in_9 ? 8'h9d : _GEN_11630; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11632 = 8'h70 == io_state_in_9 ? 8'h6 : _GEN_11631; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11633 = 8'h71 == io_state_in_9 ? 8'hb : _GEN_11632; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11634 = 8'h72 == io_state_in_9 ? 8'h1c : _GEN_11633; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11635 = 8'h73 == io_state_in_9 ? 8'h11 : _GEN_11634; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11636 = 8'h74 == io_state_in_9 ? 8'h32 : _GEN_11635; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11637 = 8'h75 == io_state_in_9 ? 8'h3f : _GEN_11636; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11638 = 8'h76 == io_state_in_9 ? 8'h28 : _GEN_11637; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11639 = 8'h77 == io_state_in_9 ? 8'h25 : _GEN_11638; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11640 = 8'h78 == io_state_in_9 ? 8'h6e : _GEN_11639; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11641 = 8'h79 == io_state_in_9 ? 8'h63 : _GEN_11640; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11642 = 8'h7a == io_state_in_9 ? 8'h74 : _GEN_11641; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11643 = 8'h7b == io_state_in_9 ? 8'h79 : _GEN_11642; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11644 = 8'h7c == io_state_in_9 ? 8'h5a : _GEN_11643; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11645 = 8'h7d == io_state_in_9 ? 8'h57 : _GEN_11644; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11646 = 8'h7e == io_state_in_9 ? 8'h40 : _GEN_11645; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11647 = 8'h7f == io_state_in_9 ? 8'h4d : _GEN_11646; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11648 = 8'h80 == io_state_in_9 ? 8'hda : _GEN_11647; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11649 = 8'h81 == io_state_in_9 ? 8'hd7 : _GEN_11648; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11650 = 8'h82 == io_state_in_9 ? 8'hc0 : _GEN_11649; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11651 = 8'h83 == io_state_in_9 ? 8'hcd : _GEN_11650; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11652 = 8'h84 == io_state_in_9 ? 8'hee : _GEN_11651; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11653 = 8'h85 == io_state_in_9 ? 8'he3 : _GEN_11652; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11654 = 8'h86 == io_state_in_9 ? 8'hf4 : _GEN_11653; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11655 = 8'h87 == io_state_in_9 ? 8'hf9 : _GEN_11654; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11656 = 8'h88 == io_state_in_9 ? 8'hb2 : _GEN_11655; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11657 = 8'h89 == io_state_in_9 ? 8'hbf : _GEN_11656; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11658 = 8'h8a == io_state_in_9 ? 8'ha8 : _GEN_11657; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11659 = 8'h8b == io_state_in_9 ? 8'ha5 : _GEN_11658; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11660 = 8'h8c == io_state_in_9 ? 8'h86 : _GEN_11659; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11661 = 8'h8d == io_state_in_9 ? 8'h8b : _GEN_11660; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11662 = 8'h8e == io_state_in_9 ? 8'h9c : _GEN_11661; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11663 = 8'h8f == io_state_in_9 ? 8'h91 : _GEN_11662; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11664 = 8'h90 == io_state_in_9 ? 8'ha : _GEN_11663; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11665 = 8'h91 == io_state_in_9 ? 8'h7 : _GEN_11664; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11666 = 8'h92 == io_state_in_9 ? 8'h10 : _GEN_11665; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11667 = 8'h93 == io_state_in_9 ? 8'h1d : _GEN_11666; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11668 = 8'h94 == io_state_in_9 ? 8'h3e : _GEN_11667; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11669 = 8'h95 == io_state_in_9 ? 8'h33 : _GEN_11668; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11670 = 8'h96 == io_state_in_9 ? 8'h24 : _GEN_11669; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11671 = 8'h97 == io_state_in_9 ? 8'h29 : _GEN_11670; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11672 = 8'h98 == io_state_in_9 ? 8'h62 : _GEN_11671; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11673 = 8'h99 == io_state_in_9 ? 8'h6f : _GEN_11672; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11674 = 8'h9a == io_state_in_9 ? 8'h78 : _GEN_11673; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11675 = 8'h9b == io_state_in_9 ? 8'h75 : _GEN_11674; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11676 = 8'h9c == io_state_in_9 ? 8'h56 : _GEN_11675; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11677 = 8'h9d == io_state_in_9 ? 8'h5b : _GEN_11676; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11678 = 8'h9e == io_state_in_9 ? 8'h4c : _GEN_11677; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11679 = 8'h9f == io_state_in_9 ? 8'h41 : _GEN_11678; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11680 = 8'ha0 == io_state_in_9 ? 8'h61 : _GEN_11679; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11681 = 8'ha1 == io_state_in_9 ? 8'h6c : _GEN_11680; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11682 = 8'ha2 == io_state_in_9 ? 8'h7b : _GEN_11681; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11683 = 8'ha3 == io_state_in_9 ? 8'h76 : _GEN_11682; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11684 = 8'ha4 == io_state_in_9 ? 8'h55 : _GEN_11683; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11685 = 8'ha5 == io_state_in_9 ? 8'h58 : _GEN_11684; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11686 = 8'ha6 == io_state_in_9 ? 8'h4f : _GEN_11685; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11687 = 8'ha7 == io_state_in_9 ? 8'h42 : _GEN_11686; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11688 = 8'ha8 == io_state_in_9 ? 8'h9 : _GEN_11687; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11689 = 8'ha9 == io_state_in_9 ? 8'h4 : _GEN_11688; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11690 = 8'haa == io_state_in_9 ? 8'h13 : _GEN_11689; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11691 = 8'hab == io_state_in_9 ? 8'h1e : _GEN_11690; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11692 = 8'hac == io_state_in_9 ? 8'h3d : _GEN_11691; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11693 = 8'had == io_state_in_9 ? 8'h30 : _GEN_11692; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11694 = 8'hae == io_state_in_9 ? 8'h27 : _GEN_11693; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11695 = 8'haf == io_state_in_9 ? 8'h2a : _GEN_11694; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11696 = 8'hb0 == io_state_in_9 ? 8'hb1 : _GEN_11695; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11697 = 8'hb1 == io_state_in_9 ? 8'hbc : _GEN_11696; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11698 = 8'hb2 == io_state_in_9 ? 8'hab : _GEN_11697; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11699 = 8'hb3 == io_state_in_9 ? 8'ha6 : _GEN_11698; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11700 = 8'hb4 == io_state_in_9 ? 8'h85 : _GEN_11699; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11701 = 8'hb5 == io_state_in_9 ? 8'h88 : _GEN_11700; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11702 = 8'hb6 == io_state_in_9 ? 8'h9f : _GEN_11701; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11703 = 8'hb7 == io_state_in_9 ? 8'h92 : _GEN_11702; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11704 = 8'hb8 == io_state_in_9 ? 8'hd9 : _GEN_11703; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11705 = 8'hb9 == io_state_in_9 ? 8'hd4 : _GEN_11704; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11706 = 8'hba == io_state_in_9 ? 8'hc3 : _GEN_11705; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11707 = 8'hbb == io_state_in_9 ? 8'hce : _GEN_11706; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11708 = 8'hbc == io_state_in_9 ? 8'hed : _GEN_11707; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11709 = 8'hbd == io_state_in_9 ? 8'he0 : _GEN_11708; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11710 = 8'hbe == io_state_in_9 ? 8'hf7 : _GEN_11709; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11711 = 8'hbf == io_state_in_9 ? 8'hfa : _GEN_11710; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11712 = 8'hc0 == io_state_in_9 ? 8'hb7 : _GEN_11711; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11713 = 8'hc1 == io_state_in_9 ? 8'hba : _GEN_11712; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11714 = 8'hc2 == io_state_in_9 ? 8'had : _GEN_11713; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11715 = 8'hc3 == io_state_in_9 ? 8'ha0 : _GEN_11714; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11716 = 8'hc4 == io_state_in_9 ? 8'h83 : _GEN_11715; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11717 = 8'hc5 == io_state_in_9 ? 8'h8e : _GEN_11716; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11718 = 8'hc6 == io_state_in_9 ? 8'h99 : _GEN_11717; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11719 = 8'hc7 == io_state_in_9 ? 8'h94 : _GEN_11718; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11720 = 8'hc8 == io_state_in_9 ? 8'hdf : _GEN_11719; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11721 = 8'hc9 == io_state_in_9 ? 8'hd2 : _GEN_11720; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11722 = 8'hca == io_state_in_9 ? 8'hc5 : _GEN_11721; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11723 = 8'hcb == io_state_in_9 ? 8'hc8 : _GEN_11722; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11724 = 8'hcc == io_state_in_9 ? 8'heb : _GEN_11723; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11725 = 8'hcd == io_state_in_9 ? 8'he6 : _GEN_11724; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11726 = 8'hce == io_state_in_9 ? 8'hf1 : _GEN_11725; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11727 = 8'hcf == io_state_in_9 ? 8'hfc : _GEN_11726; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11728 = 8'hd0 == io_state_in_9 ? 8'h67 : _GEN_11727; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11729 = 8'hd1 == io_state_in_9 ? 8'h6a : _GEN_11728; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11730 = 8'hd2 == io_state_in_9 ? 8'h7d : _GEN_11729; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11731 = 8'hd3 == io_state_in_9 ? 8'h70 : _GEN_11730; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11732 = 8'hd4 == io_state_in_9 ? 8'h53 : _GEN_11731; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11733 = 8'hd5 == io_state_in_9 ? 8'h5e : _GEN_11732; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11734 = 8'hd6 == io_state_in_9 ? 8'h49 : _GEN_11733; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11735 = 8'hd7 == io_state_in_9 ? 8'h44 : _GEN_11734; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11736 = 8'hd8 == io_state_in_9 ? 8'hf : _GEN_11735; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11737 = 8'hd9 == io_state_in_9 ? 8'h2 : _GEN_11736; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11738 = 8'hda == io_state_in_9 ? 8'h15 : _GEN_11737; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11739 = 8'hdb == io_state_in_9 ? 8'h18 : _GEN_11738; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11740 = 8'hdc == io_state_in_9 ? 8'h3b : _GEN_11739; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11741 = 8'hdd == io_state_in_9 ? 8'h36 : _GEN_11740; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11742 = 8'hde == io_state_in_9 ? 8'h21 : _GEN_11741; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11743 = 8'hdf == io_state_in_9 ? 8'h2c : _GEN_11742; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11744 = 8'he0 == io_state_in_9 ? 8'hc : _GEN_11743; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11745 = 8'he1 == io_state_in_9 ? 8'h1 : _GEN_11744; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11746 = 8'he2 == io_state_in_9 ? 8'h16 : _GEN_11745; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11747 = 8'he3 == io_state_in_9 ? 8'h1b : _GEN_11746; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11748 = 8'he4 == io_state_in_9 ? 8'h38 : _GEN_11747; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11749 = 8'he5 == io_state_in_9 ? 8'h35 : _GEN_11748; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11750 = 8'he6 == io_state_in_9 ? 8'h22 : _GEN_11749; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11751 = 8'he7 == io_state_in_9 ? 8'h2f : _GEN_11750; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11752 = 8'he8 == io_state_in_9 ? 8'h64 : _GEN_11751; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11753 = 8'he9 == io_state_in_9 ? 8'h69 : _GEN_11752; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11754 = 8'hea == io_state_in_9 ? 8'h7e : _GEN_11753; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11755 = 8'heb == io_state_in_9 ? 8'h73 : _GEN_11754; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11756 = 8'hec == io_state_in_9 ? 8'h50 : _GEN_11755; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11757 = 8'hed == io_state_in_9 ? 8'h5d : _GEN_11756; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11758 = 8'hee == io_state_in_9 ? 8'h4a : _GEN_11757; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11759 = 8'hef == io_state_in_9 ? 8'h47 : _GEN_11758; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11760 = 8'hf0 == io_state_in_9 ? 8'hdc : _GEN_11759; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11761 = 8'hf1 == io_state_in_9 ? 8'hd1 : _GEN_11760; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11762 = 8'hf2 == io_state_in_9 ? 8'hc6 : _GEN_11761; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11763 = 8'hf3 == io_state_in_9 ? 8'hcb : _GEN_11762; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11764 = 8'hf4 == io_state_in_9 ? 8'he8 : _GEN_11763; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11765 = 8'hf5 == io_state_in_9 ? 8'he5 : _GEN_11764; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11766 = 8'hf6 == io_state_in_9 ? 8'hf2 : _GEN_11765; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11767 = 8'hf7 == io_state_in_9 ? 8'hff : _GEN_11766; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11768 = 8'hf8 == io_state_in_9 ? 8'hb4 : _GEN_11767; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11769 = 8'hf9 == io_state_in_9 ? 8'hb9 : _GEN_11768; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11770 = 8'hfa == io_state_in_9 ? 8'hae : _GEN_11769; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11771 = 8'hfb == io_state_in_9 ? 8'ha3 : _GEN_11770; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11772 = 8'hfc == io_state_in_9 ? 8'h80 : _GEN_11771; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11773 = 8'hfd == io_state_in_9 ? 8'h8d : _GEN_11772; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11774 = 8'hfe == io_state_in_9 ? 8'h9a : _GEN_11773; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _GEN_11775 = 8'hff == io_state_in_9 ? 8'h97 : _GEN_11774; // @[InvMixColumns.scala 139:{42,42}]
  wire [7:0] _tmp_state_11_T = _GEN_11519 ^ _GEN_11775; // @[InvMixColumns.scala 139:42]
  wire [7:0] _GEN_11777 = 8'h1 == io_state_in_10 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11778 = 8'h2 == io_state_in_10 ? 8'h12 : _GEN_11777; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11779 = 8'h3 == io_state_in_10 ? 8'h1b : _GEN_11778; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11780 = 8'h4 == io_state_in_10 ? 8'h24 : _GEN_11779; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11781 = 8'h5 == io_state_in_10 ? 8'h2d : _GEN_11780; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11782 = 8'h6 == io_state_in_10 ? 8'h36 : _GEN_11781; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11783 = 8'h7 == io_state_in_10 ? 8'h3f : _GEN_11782; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11784 = 8'h8 == io_state_in_10 ? 8'h48 : _GEN_11783; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11785 = 8'h9 == io_state_in_10 ? 8'h41 : _GEN_11784; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11786 = 8'ha == io_state_in_10 ? 8'h5a : _GEN_11785; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11787 = 8'hb == io_state_in_10 ? 8'h53 : _GEN_11786; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11788 = 8'hc == io_state_in_10 ? 8'h6c : _GEN_11787; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11789 = 8'hd == io_state_in_10 ? 8'h65 : _GEN_11788; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11790 = 8'he == io_state_in_10 ? 8'h7e : _GEN_11789; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11791 = 8'hf == io_state_in_10 ? 8'h77 : _GEN_11790; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11792 = 8'h10 == io_state_in_10 ? 8'h90 : _GEN_11791; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11793 = 8'h11 == io_state_in_10 ? 8'h99 : _GEN_11792; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11794 = 8'h12 == io_state_in_10 ? 8'h82 : _GEN_11793; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11795 = 8'h13 == io_state_in_10 ? 8'h8b : _GEN_11794; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11796 = 8'h14 == io_state_in_10 ? 8'hb4 : _GEN_11795; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11797 = 8'h15 == io_state_in_10 ? 8'hbd : _GEN_11796; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11798 = 8'h16 == io_state_in_10 ? 8'ha6 : _GEN_11797; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11799 = 8'h17 == io_state_in_10 ? 8'haf : _GEN_11798; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11800 = 8'h18 == io_state_in_10 ? 8'hd8 : _GEN_11799; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11801 = 8'h19 == io_state_in_10 ? 8'hd1 : _GEN_11800; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11802 = 8'h1a == io_state_in_10 ? 8'hca : _GEN_11801; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11803 = 8'h1b == io_state_in_10 ? 8'hc3 : _GEN_11802; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11804 = 8'h1c == io_state_in_10 ? 8'hfc : _GEN_11803; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11805 = 8'h1d == io_state_in_10 ? 8'hf5 : _GEN_11804; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11806 = 8'h1e == io_state_in_10 ? 8'hee : _GEN_11805; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11807 = 8'h1f == io_state_in_10 ? 8'he7 : _GEN_11806; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11808 = 8'h20 == io_state_in_10 ? 8'h3b : _GEN_11807; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11809 = 8'h21 == io_state_in_10 ? 8'h32 : _GEN_11808; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11810 = 8'h22 == io_state_in_10 ? 8'h29 : _GEN_11809; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11811 = 8'h23 == io_state_in_10 ? 8'h20 : _GEN_11810; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11812 = 8'h24 == io_state_in_10 ? 8'h1f : _GEN_11811; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11813 = 8'h25 == io_state_in_10 ? 8'h16 : _GEN_11812; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11814 = 8'h26 == io_state_in_10 ? 8'hd : _GEN_11813; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11815 = 8'h27 == io_state_in_10 ? 8'h4 : _GEN_11814; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11816 = 8'h28 == io_state_in_10 ? 8'h73 : _GEN_11815; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11817 = 8'h29 == io_state_in_10 ? 8'h7a : _GEN_11816; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11818 = 8'h2a == io_state_in_10 ? 8'h61 : _GEN_11817; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11819 = 8'h2b == io_state_in_10 ? 8'h68 : _GEN_11818; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11820 = 8'h2c == io_state_in_10 ? 8'h57 : _GEN_11819; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11821 = 8'h2d == io_state_in_10 ? 8'h5e : _GEN_11820; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11822 = 8'h2e == io_state_in_10 ? 8'h45 : _GEN_11821; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11823 = 8'h2f == io_state_in_10 ? 8'h4c : _GEN_11822; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11824 = 8'h30 == io_state_in_10 ? 8'hab : _GEN_11823; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11825 = 8'h31 == io_state_in_10 ? 8'ha2 : _GEN_11824; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11826 = 8'h32 == io_state_in_10 ? 8'hb9 : _GEN_11825; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11827 = 8'h33 == io_state_in_10 ? 8'hb0 : _GEN_11826; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11828 = 8'h34 == io_state_in_10 ? 8'h8f : _GEN_11827; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11829 = 8'h35 == io_state_in_10 ? 8'h86 : _GEN_11828; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11830 = 8'h36 == io_state_in_10 ? 8'h9d : _GEN_11829; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11831 = 8'h37 == io_state_in_10 ? 8'h94 : _GEN_11830; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11832 = 8'h38 == io_state_in_10 ? 8'he3 : _GEN_11831; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11833 = 8'h39 == io_state_in_10 ? 8'hea : _GEN_11832; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11834 = 8'h3a == io_state_in_10 ? 8'hf1 : _GEN_11833; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11835 = 8'h3b == io_state_in_10 ? 8'hf8 : _GEN_11834; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11836 = 8'h3c == io_state_in_10 ? 8'hc7 : _GEN_11835; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11837 = 8'h3d == io_state_in_10 ? 8'hce : _GEN_11836; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11838 = 8'h3e == io_state_in_10 ? 8'hd5 : _GEN_11837; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11839 = 8'h3f == io_state_in_10 ? 8'hdc : _GEN_11838; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11840 = 8'h40 == io_state_in_10 ? 8'h76 : _GEN_11839; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11841 = 8'h41 == io_state_in_10 ? 8'h7f : _GEN_11840; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11842 = 8'h42 == io_state_in_10 ? 8'h64 : _GEN_11841; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11843 = 8'h43 == io_state_in_10 ? 8'h6d : _GEN_11842; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11844 = 8'h44 == io_state_in_10 ? 8'h52 : _GEN_11843; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11845 = 8'h45 == io_state_in_10 ? 8'h5b : _GEN_11844; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11846 = 8'h46 == io_state_in_10 ? 8'h40 : _GEN_11845; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11847 = 8'h47 == io_state_in_10 ? 8'h49 : _GEN_11846; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11848 = 8'h48 == io_state_in_10 ? 8'h3e : _GEN_11847; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11849 = 8'h49 == io_state_in_10 ? 8'h37 : _GEN_11848; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11850 = 8'h4a == io_state_in_10 ? 8'h2c : _GEN_11849; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11851 = 8'h4b == io_state_in_10 ? 8'h25 : _GEN_11850; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11852 = 8'h4c == io_state_in_10 ? 8'h1a : _GEN_11851; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11853 = 8'h4d == io_state_in_10 ? 8'h13 : _GEN_11852; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11854 = 8'h4e == io_state_in_10 ? 8'h8 : _GEN_11853; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11855 = 8'h4f == io_state_in_10 ? 8'h1 : _GEN_11854; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11856 = 8'h50 == io_state_in_10 ? 8'he6 : _GEN_11855; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11857 = 8'h51 == io_state_in_10 ? 8'hef : _GEN_11856; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11858 = 8'h52 == io_state_in_10 ? 8'hf4 : _GEN_11857; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11859 = 8'h53 == io_state_in_10 ? 8'hfd : _GEN_11858; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11860 = 8'h54 == io_state_in_10 ? 8'hc2 : _GEN_11859; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11861 = 8'h55 == io_state_in_10 ? 8'hcb : _GEN_11860; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11862 = 8'h56 == io_state_in_10 ? 8'hd0 : _GEN_11861; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11863 = 8'h57 == io_state_in_10 ? 8'hd9 : _GEN_11862; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11864 = 8'h58 == io_state_in_10 ? 8'hae : _GEN_11863; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11865 = 8'h59 == io_state_in_10 ? 8'ha7 : _GEN_11864; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11866 = 8'h5a == io_state_in_10 ? 8'hbc : _GEN_11865; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11867 = 8'h5b == io_state_in_10 ? 8'hb5 : _GEN_11866; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11868 = 8'h5c == io_state_in_10 ? 8'h8a : _GEN_11867; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11869 = 8'h5d == io_state_in_10 ? 8'h83 : _GEN_11868; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11870 = 8'h5e == io_state_in_10 ? 8'h98 : _GEN_11869; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11871 = 8'h5f == io_state_in_10 ? 8'h91 : _GEN_11870; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11872 = 8'h60 == io_state_in_10 ? 8'h4d : _GEN_11871; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11873 = 8'h61 == io_state_in_10 ? 8'h44 : _GEN_11872; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11874 = 8'h62 == io_state_in_10 ? 8'h5f : _GEN_11873; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11875 = 8'h63 == io_state_in_10 ? 8'h56 : _GEN_11874; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11876 = 8'h64 == io_state_in_10 ? 8'h69 : _GEN_11875; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11877 = 8'h65 == io_state_in_10 ? 8'h60 : _GEN_11876; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11878 = 8'h66 == io_state_in_10 ? 8'h7b : _GEN_11877; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11879 = 8'h67 == io_state_in_10 ? 8'h72 : _GEN_11878; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11880 = 8'h68 == io_state_in_10 ? 8'h5 : _GEN_11879; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11881 = 8'h69 == io_state_in_10 ? 8'hc : _GEN_11880; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11882 = 8'h6a == io_state_in_10 ? 8'h17 : _GEN_11881; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11883 = 8'h6b == io_state_in_10 ? 8'h1e : _GEN_11882; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11884 = 8'h6c == io_state_in_10 ? 8'h21 : _GEN_11883; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11885 = 8'h6d == io_state_in_10 ? 8'h28 : _GEN_11884; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11886 = 8'h6e == io_state_in_10 ? 8'h33 : _GEN_11885; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11887 = 8'h6f == io_state_in_10 ? 8'h3a : _GEN_11886; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11888 = 8'h70 == io_state_in_10 ? 8'hdd : _GEN_11887; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11889 = 8'h71 == io_state_in_10 ? 8'hd4 : _GEN_11888; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11890 = 8'h72 == io_state_in_10 ? 8'hcf : _GEN_11889; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11891 = 8'h73 == io_state_in_10 ? 8'hc6 : _GEN_11890; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11892 = 8'h74 == io_state_in_10 ? 8'hf9 : _GEN_11891; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11893 = 8'h75 == io_state_in_10 ? 8'hf0 : _GEN_11892; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11894 = 8'h76 == io_state_in_10 ? 8'heb : _GEN_11893; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11895 = 8'h77 == io_state_in_10 ? 8'he2 : _GEN_11894; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11896 = 8'h78 == io_state_in_10 ? 8'h95 : _GEN_11895; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11897 = 8'h79 == io_state_in_10 ? 8'h9c : _GEN_11896; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11898 = 8'h7a == io_state_in_10 ? 8'h87 : _GEN_11897; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11899 = 8'h7b == io_state_in_10 ? 8'h8e : _GEN_11898; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11900 = 8'h7c == io_state_in_10 ? 8'hb1 : _GEN_11899; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11901 = 8'h7d == io_state_in_10 ? 8'hb8 : _GEN_11900; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11902 = 8'h7e == io_state_in_10 ? 8'ha3 : _GEN_11901; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11903 = 8'h7f == io_state_in_10 ? 8'haa : _GEN_11902; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11904 = 8'h80 == io_state_in_10 ? 8'hec : _GEN_11903; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11905 = 8'h81 == io_state_in_10 ? 8'he5 : _GEN_11904; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11906 = 8'h82 == io_state_in_10 ? 8'hfe : _GEN_11905; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11907 = 8'h83 == io_state_in_10 ? 8'hf7 : _GEN_11906; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11908 = 8'h84 == io_state_in_10 ? 8'hc8 : _GEN_11907; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11909 = 8'h85 == io_state_in_10 ? 8'hc1 : _GEN_11908; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11910 = 8'h86 == io_state_in_10 ? 8'hda : _GEN_11909; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11911 = 8'h87 == io_state_in_10 ? 8'hd3 : _GEN_11910; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11912 = 8'h88 == io_state_in_10 ? 8'ha4 : _GEN_11911; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11913 = 8'h89 == io_state_in_10 ? 8'had : _GEN_11912; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11914 = 8'h8a == io_state_in_10 ? 8'hb6 : _GEN_11913; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11915 = 8'h8b == io_state_in_10 ? 8'hbf : _GEN_11914; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11916 = 8'h8c == io_state_in_10 ? 8'h80 : _GEN_11915; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11917 = 8'h8d == io_state_in_10 ? 8'h89 : _GEN_11916; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11918 = 8'h8e == io_state_in_10 ? 8'h92 : _GEN_11917; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11919 = 8'h8f == io_state_in_10 ? 8'h9b : _GEN_11918; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11920 = 8'h90 == io_state_in_10 ? 8'h7c : _GEN_11919; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11921 = 8'h91 == io_state_in_10 ? 8'h75 : _GEN_11920; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11922 = 8'h92 == io_state_in_10 ? 8'h6e : _GEN_11921; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11923 = 8'h93 == io_state_in_10 ? 8'h67 : _GEN_11922; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11924 = 8'h94 == io_state_in_10 ? 8'h58 : _GEN_11923; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11925 = 8'h95 == io_state_in_10 ? 8'h51 : _GEN_11924; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11926 = 8'h96 == io_state_in_10 ? 8'h4a : _GEN_11925; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11927 = 8'h97 == io_state_in_10 ? 8'h43 : _GEN_11926; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11928 = 8'h98 == io_state_in_10 ? 8'h34 : _GEN_11927; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11929 = 8'h99 == io_state_in_10 ? 8'h3d : _GEN_11928; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11930 = 8'h9a == io_state_in_10 ? 8'h26 : _GEN_11929; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11931 = 8'h9b == io_state_in_10 ? 8'h2f : _GEN_11930; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11932 = 8'h9c == io_state_in_10 ? 8'h10 : _GEN_11931; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11933 = 8'h9d == io_state_in_10 ? 8'h19 : _GEN_11932; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11934 = 8'h9e == io_state_in_10 ? 8'h2 : _GEN_11933; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11935 = 8'h9f == io_state_in_10 ? 8'hb : _GEN_11934; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11936 = 8'ha0 == io_state_in_10 ? 8'hd7 : _GEN_11935; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11937 = 8'ha1 == io_state_in_10 ? 8'hde : _GEN_11936; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11938 = 8'ha2 == io_state_in_10 ? 8'hc5 : _GEN_11937; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11939 = 8'ha3 == io_state_in_10 ? 8'hcc : _GEN_11938; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11940 = 8'ha4 == io_state_in_10 ? 8'hf3 : _GEN_11939; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11941 = 8'ha5 == io_state_in_10 ? 8'hfa : _GEN_11940; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11942 = 8'ha6 == io_state_in_10 ? 8'he1 : _GEN_11941; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11943 = 8'ha7 == io_state_in_10 ? 8'he8 : _GEN_11942; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11944 = 8'ha8 == io_state_in_10 ? 8'h9f : _GEN_11943; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11945 = 8'ha9 == io_state_in_10 ? 8'h96 : _GEN_11944; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11946 = 8'haa == io_state_in_10 ? 8'h8d : _GEN_11945; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11947 = 8'hab == io_state_in_10 ? 8'h84 : _GEN_11946; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11948 = 8'hac == io_state_in_10 ? 8'hbb : _GEN_11947; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11949 = 8'had == io_state_in_10 ? 8'hb2 : _GEN_11948; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11950 = 8'hae == io_state_in_10 ? 8'ha9 : _GEN_11949; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11951 = 8'haf == io_state_in_10 ? 8'ha0 : _GEN_11950; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11952 = 8'hb0 == io_state_in_10 ? 8'h47 : _GEN_11951; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11953 = 8'hb1 == io_state_in_10 ? 8'h4e : _GEN_11952; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11954 = 8'hb2 == io_state_in_10 ? 8'h55 : _GEN_11953; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11955 = 8'hb3 == io_state_in_10 ? 8'h5c : _GEN_11954; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11956 = 8'hb4 == io_state_in_10 ? 8'h63 : _GEN_11955; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11957 = 8'hb5 == io_state_in_10 ? 8'h6a : _GEN_11956; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11958 = 8'hb6 == io_state_in_10 ? 8'h71 : _GEN_11957; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11959 = 8'hb7 == io_state_in_10 ? 8'h78 : _GEN_11958; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11960 = 8'hb8 == io_state_in_10 ? 8'hf : _GEN_11959; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11961 = 8'hb9 == io_state_in_10 ? 8'h6 : _GEN_11960; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11962 = 8'hba == io_state_in_10 ? 8'h1d : _GEN_11961; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11963 = 8'hbb == io_state_in_10 ? 8'h14 : _GEN_11962; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11964 = 8'hbc == io_state_in_10 ? 8'h2b : _GEN_11963; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11965 = 8'hbd == io_state_in_10 ? 8'h22 : _GEN_11964; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11966 = 8'hbe == io_state_in_10 ? 8'h39 : _GEN_11965; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11967 = 8'hbf == io_state_in_10 ? 8'h30 : _GEN_11966; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11968 = 8'hc0 == io_state_in_10 ? 8'h9a : _GEN_11967; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11969 = 8'hc1 == io_state_in_10 ? 8'h93 : _GEN_11968; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11970 = 8'hc2 == io_state_in_10 ? 8'h88 : _GEN_11969; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11971 = 8'hc3 == io_state_in_10 ? 8'h81 : _GEN_11970; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11972 = 8'hc4 == io_state_in_10 ? 8'hbe : _GEN_11971; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11973 = 8'hc5 == io_state_in_10 ? 8'hb7 : _GEN_11972; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11974 = 8'hc6 == io_state_in_10 ? 8'hac : _GEN_11973; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11975 = 8'hc7 == io_state_in_10 ? 8'ha5 : _GEN_11974; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11976 = 8'hc8 == io_state_in_10 ? 8'hd2 : _GEN_11975; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11977 = 8'hc9 == io_state_in_10 ? 8'hdb : _GEN_11976; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11978 = 8'hca == io_state_in_10 ? 8'hc0 : _GEN_11977; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11979 = 8'hcb == io_state_in_10 ? 8'hc9 : _GEN_11978; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11980 = 8'hcc == io_state_in_10 ? 8'hf6 : _GEN_11979; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11981 = 8'hcd == io_state_in_10 ? 8'hff : _GEN_11980; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11982 = 8'hce == io_state_in_10 ? 8'he4 : _GEN_11981; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11983 = 8'hcf == io_state_in_10 ? 8'hed : _GEN_11982; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11984 = 8'hd0 == io_state_in_10 ? 8'ha : _GEN_11983; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11985 = 8'hd1 == io_state_in_10 ? 8'h3 : _GEN_11984; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11986 = 8'hd2 == io_state_in_10 ? 8'h18 : _GEN_11985; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11987 = 8'hd3 == io_state_in_10 ? 8'h11 : _GEN_11986; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11988 = 8'hd4 == io_state_in_10 ? 8'h2e : _GEN_11987; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11989 = 8'hd5 == io_state_in_10 ? 8'h27 : _GEN_11988; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11990 = 8'hd6 == io_state_in_10 ? 8'h3c : _GEN_11989; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11991 = 8'hd7 == io_state_in_10 ? 8'h35 : _GEN_11990; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11992 = 8'hd8 == io_state_in_10 ? 8'h42 : _GEN_11991; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11993 = 8'hd9 == io_state_in_10 ? 8'h4b : _GEN_11992; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11994 = 8'hda == io_state_in_10 ? 8'h50 : _GEN_11993; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11995 = 8'hdb == io_state_in_10 ? 8'h59 : _GEN_11994; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11996 = 8'hdc == io_state_in_10 ? 8'h66 : _GEN_11995; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11997 = 8'hdd == io_state_in_10 ? 8'h6f : _GEN_11996; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11998 = 8'hde == io_state_in_10 ? 8'h74 : _GEN_11997; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_11999 = 8'hdf == io_state_in_10 ? 8'h7d : _GEN_11998; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12000 = 8'he0 == io_state_in_10 ? 8'ha1 : _GEN_11999; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12001 = 8'he1 == io_state_in_10 ? 8'ha8 : _GEN_12000; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12002 = 8'he2 == io_state_in_10 ? 8'hb3 : _GEN_12001; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12003 = 8'he3 == io_state_in_10 ? 8'hba : _GEN_12002; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12004 = 8'he4 == io_state_in_10 ? 8'h85 : _GEN_12003; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12005 = 8'he5 == io_state_in_10 ? 8'h8c : _GEN_12004; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12006 = 8'he6 == io_state_in_10 ? 8'h97 : _GEN_12005; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12007 = 8'he7 == io_state_in_10 ? 8'h9e : _GEN_12006; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12008 = 8'he8 == io_state_in_10 ? 8'he9 : _GEN_12007; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12009 = 8'he9 == io_state_in_10 ? 8'he0 : _GEN_12008; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12010 = 8'hea == io_state_in_10 ? 8'hfb : _GEN_12009; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12011 = 8'heb == io_state_in_10 ? 8'hf2 : _GEN_12010; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12012 = 8'hec == io_state_in_10 ? 8'hcd : _GEN_12011; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12013 = 8'hed == io_state_in_10 ? 8'hc4 : _GEN_12012; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12014 = 8'hee == io_state_in_10 ? 8'hdf : _GEN_12013; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12015 = 8'hef == io_state_in_10 ? 8'hd6 : _GEN_12014; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12016 = 8'hf0 == io_state_in_10 ? 8'h31 : _GEN_12015; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12017 = 8'hf1 == io_state_in_10 ? 8'h38 : _GEN_12016; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12018 = 8'hf2 == io_state_in_10 ? 8'h23 : _GEN_12017; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12019 = 8'hf3 == io_state_in_10 ? 8'h2a : _GEN_12018; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12020 = 8'hf4 == io_state_in_10 ? 8'h15 : _GEN_12019; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12021 = 8'hf5 == io_state_in_10 ? 8'h1c : _GEN_12020; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12022 = 8'hf6 == io_state_in_10 ? 8'h7 : _GEN_12021; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12023 = 8'hf7 == io_state_in_10 ? 8'he : _GEN_12022; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12024 = 8'hf8 == io_state_in_10 ? 8'h79 : _GEN_12023; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12025 = 8'hf9 == io_state_in_10 ? 8'h70 : _GEN_12024; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12026 = 8'hfa == io_state_in_10 ? 8'h6b : _GEN_12025; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12027 = 8'hfb == io_state_in_10 ? 8'h62 : _GEN_12026; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12028 = 8'hfc == io_state_in_10 ? 8'h5d : _GEN_12027; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12029 = 8'hfd == io_state_in_10 ? 8'h54 : _GEN_12028; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12030 = 8'hfe == io_state_in_10 ? 8'h4f : _GEN_12029; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _GEN_12031 = 8'hff == io_state_in_10 ? 8'h46 : _GEN_12030; // @[InvMixColumns.scala 139:{66,66}]
  wire [7:0] _tmp_state_11_T_1 = _tmp_state_11_T ^ _GEN_12031; // @[InvMixColumns.scala 139:66]
  wire [7:0] _GEN_12033 = 8'h1 == io_state_in_11 ? 8'he : 8'h0; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12034 = 8'h2 == io_state_in_11 ? 8'h1c : _GEN_12033; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12035 = 8'h3 == io_state_in_11 ? 8'h12 : _GEN_12034; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12036 = 8'h4 == io_state_in_11 ? 8'h38 : _GEN_12035; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12037 = 8'h5 == io_state_in_11 ? 8'h36 : _GEN_12036; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12038 = 8'h6 == io_state_in_11 ? 8'h24 : _GEN_12037; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12039 = 8'h7 == io_state_in_11 ? 8'h2a : _GEN_12038; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12040 = 8'h8 == io_state_in_11 ? 8'h70 : _GEN_12039; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12041 = 8'h9 == io_state_in_11 ? 8'h7e : _GEN_12040; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12042 = 8'ha == io_state_in_11 ? 8'h6c : _GEN_12041; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12043 = 8'hb == io_state_in_11 ? 8'h62 : _GEN_12042; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12044 = 8'hc == io_state_in_11 ? 8'h48 : _GEN_12043; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12045 = 8'hd == io_state_in_11 ? 8'h46 : _GEN_12044; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12046 = 8'he == io_state_in_11 ? 8'h54 : _GEN_12045; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12047 = 8'hf == io_state_in_11 ? 8'h5a : _GEN_12046; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12048 = 8'h10 == io_state_in_11 ? 8'he0 : _GEN_12047; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12049 = 8'h11 == io_state_in_11 ? 8'hee : _GEN_12048; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12050 = 8'h12 == io_state_in_11 ? 8'hfc : _GEN_12049; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12051 = 8'h13 == io_state_in_11 ? 8'hf2 : _GEN_12050; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12052 = 8'h14 == io_state_in_11 ? 8'hd8 : _GEN_12051; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12053 = 8'h15 == io_state_in_11 ? 8'hd6 : _GEN_12052; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12054 = 8'h16 == io_state_in_11 ? 8'hc4 : _GEN_12053; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12055 = 8'h17 == io_state_in_11 ? 8'hca : _GEN_12054; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12056 = 8'h18 == io_state_in_11 ? 8'h90 : _GEN_12055; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12057 = 8'h19 == io_state_in_11 ? 8'h9e : _GEN_12056; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12058 = 8'h1a == io_state_in_11 ? 8'h8c : _GEN_12057; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12059 = 8'h1b == io_state_in_11 ? 8'h82 : _GEN_12058; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12060 = 8'h1c == io_state_in_11 ? 8'ha8 : _GEN_12059; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12061 = 8'h1d == io_state_in_11 ? 8'ha6 : _GEN_12060; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12062 = 8'h1e == io_state_in_11 ? 8'hb4 : _GEN_12061; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12063 = 8'h1f == io_state_in_11 ? 8'hba : _GEN_12062; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12064 = 8'h20 == io_state_in_11 ? 8'hdb : _GEN_12063; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12065 = 8'h21 == io_state_in_11 ? 8'hd5 : _GEN_12064; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12066 = 8'h22 == io_state_in_11 ? 8'hc7 : _GEN_12065; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12067 = 8'h23 == io_state_in_11 ? 8'hc9 : _GEN_12066; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12068 = 8'h24 == io_state_in_11 ? 8'he3 : _GEN_12067; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12069 = 8'h25 == io_state_in_11 ? 8'hed : _GEN_12068; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12070 = 8'h26 == io_state_in_11 ? 8'hff : _GEN_12069; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12071 = 8'h27 == io_state_in_11 ? 8'hf1 : _GEN_12070; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12072 = 8'h28 == io_state_in_11 ? 8'hab : _GEN_12071; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12073 = 8'h29 == io_state_in_11 ? 8'ha5 : _GEN_12072; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12074 = 8'h2a == io_state_in_11 ? 8'hb7 : _GEN_12073; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12075 = 8'h2b == io_state_in_11 ? 8'hb9 : _GEN_12074; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12076 = 8'h2c == io_state_in_11 ? 8'h93 : _GEN_12075; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12077 = 8'h2d == io_state_in_11 ? 8'h9d : _GEN_12076; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12078 = 8'h2e == io_state_in_11 ? 8'h8f : _GEN_12077; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12079 = 8'h2f == io_state_in_11 ? 8'h81 : _GEN_12078; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12080 = 8'h30 == io_state_in_11 ? 8'h3b : _GEN_12079; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12081 = 8'h31 == io_state_in_11 ? 8'h35 : _GEN_12080; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12082 = 8'h32 == io_state_in_11 ? 8'h27 : _GEN_12081; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12083 = 8'h33 == io_state_in_11 ? 8'h29 : _GEN_12082; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12084 = 8'h34 == io_state_in_11 ? 8'h3 : _GEN_12083; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12085 = 8'h35 == io_state_in_11 ? 8'hd : _GEN_12084; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12086 = 8'h36 == io_state_in_11 ? 8'h1f : _GEN_12085; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12087 = 8'h37 == io_state_in_11 ? 8'h11 : _GEN_12086; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12088 = 8'h38 == io_state_in_11 ? 8'h4b : _GEN_12087; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12089 = 8'h39 == io_state_in_11 ? 8'h45 : _GEN_12088; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12090 = 8'h3a == io_state_in_11 ? 8'h57 : _GEN_12089; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12091 = 8'h3b == io_state_in_11 ? 8'h59 : _GEN_12090; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12092 = 8'h3c == io_state_in_11 ? 8'h73 : _GEN_12091; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12093 = 8'h3d == io_state_in_11 ? 8'h7d : _GEN_12092; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12094 = 8'h3e == io_state_in_11 ? 8'h6f : _GEN_12093; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12095 = 8'h3f == io_state_in_11 ? 8'h61 : _GEN_12094; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12096 = 8'h40 == io_state_in_11 ? 8'had : _GEN_12095; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12097 = 8'h41 == io_state_in_11 ? 8'ha3 : _GEN_12096; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12098 = 8'h42 == io_state_in_11 ? 8'hb1 : _GEN_12097; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12099 = 8'h43 == io_state_in_11 ? 8'hbf : _GEN_12098; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12100 = 8'h44 == io_state_in_11 ? 8'h95 : _GEN_12099; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12101 = 8'h45 == io_state_in_11 ? 8'h9b : _GEN_12100; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12102 = 8'h46 == io_state_in_11 ? 8'h89 : _GEN_12101; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12103 = 8'h47 == io_state_in_11 ? 8'h87 : _GEN_12102; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12104 = 8'h48 == io_state_in_11 ? 8'hdd : _GEN_12103; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12105 = 8'h49 == io_state_in_11 ? 8'hd3 : _GEN_12104; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12106 = 8'h4a == io_state_in_11 ? 8'hc1 : _GEN_12105; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12107 = 8'h4b == io_state_in_11 ? 8'hcf : _GEN_12106; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12108 = 8'h4c == io_state_in_11 ? 8'he5 : _GEN_12107; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12109 = 8'h4d == io_state_in_11 ? 8'heb : _GEN_12108; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12110 = 8'h4e == io_state_in_11 ? 8'hf9 : _GEN_12109; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12111 = 8'h4f == io_state_in_11 ? 8'hf7 : _GEN_12110; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12112 = 8'h50 == io_state_in_11 ? 8'h4d : _GEN_12111; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12113 = 8'h51 == io_state_in_11 ? 8'h43 : _GEN_12112; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12114 = 8'h52 == io_state_in_11 ? 8'h51 : _GEN_12113; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12115 = 8'h53 == io_state_in_11 ? 8'h5f : _GEN_12114; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12116 = 8'h54 == io_state_in_11 ? 8'h75 : _GEN_12115; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12117 = 8'h55 == io_state_in_11 ? 8'h7b : _GEN_12116; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12118 = 8'h56 == io_state_in_11 ? 8'h69 : _GEN_12117; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12119 = 8'h57 == io_state_in_11 ? 8'h67 : _GEN_12118; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12120 = 8'h58 == io_state_in_11 ? 8'h3d : _GEN_12119; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12121 = 8'h59 == io_state_in_11 ? 8'h33 : _GEN_12120; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12122 = 8'h5a == io_state_in_11 ? 8'h21 : _GEN_12121; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12123 = 8'h5b == io_state_in_11 ? 8'h2f : _GEN_12122; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12124 = 8'h5c == io_state_in_11 ? 8'h5 : _GEN_12123; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12125 = 8'h5d == io_state_in_11 ? 8'hb : _GEN_12124; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12126 = 8'h5e == io_state_in_11 ? 8'h19 : _GEN_12125; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12127 = 8'h5f == io_state_in_11 ? 8'h17 : _GEN_12126; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12128 = 8'h60 == io_state_in_11 ? 8'h76 : _GEN_12127; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12129 = 8'h61 == io_state_in_11 ? 8'h78 : _GEN_12128; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12130 = 8'h62 == io_state_in_11 ? 8'h6a : _GEN_12129; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12131 = 8'h63 == io_state_in_11 ? 8'h64 : _GEN_12130; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12132 = 8'h64 == io_state_in_11 ? 8'h4e : _GEN_12131; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12133 = 8'h65 == io_state_in_11 ? 8'h40 : _GEN_12132; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12134 = 8'h66 == io_state_in_11 ? 8'h52 : _GEN_12133; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12135 = 8'h67 == io_state_in_11 ? 8'h5c : _GEN_12134; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12136 = 8'h68 == io_state_in_11 ? 8'h6 : _GEN_12135; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12137 = 8'h69 == io_state_in_11 ? 8'h8 : _GEN_12136; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12138 = 8'h6a == io_state_in_11 ? 8'h1a : _GEN_12137; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12139 = 8'h6b == io_state_in_11 ? 8'h14 : _GEN_12138; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12140 = 8'h6c == io_state_in_11 ? 8'h3e : _GEN_12139; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12141 = 8'h6d == io_state_in_11 ? 8'h30 : _GEN_12140; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12142 = 8'h6e == io_state_in_11 ? 8'h22 : _GEN_12141; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12143 = 8'h6f == io_state_in_11 ? 8'h2c : _GEN_12142; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12144 = 8'h70 == io_state_in_11 ? 8'h96 : _GEN_12143; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12145 = 8'h71 == io_state_in_11 ? 8'h98 : _GEN_12144; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12146 = 8'h72 == io_state_in_11 ? 8'h8a : _GEN_12145; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12147 = 8'h73 == io_state_in_11 ? 8'h84 : _GEN_12146; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12148 = 8'h74 == io_state_in_11 ? 8'hae : _GEN_12147; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12149 = 8'h75 == io_state_in_11 ? 8'ha0 : _GEN_12148; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12150 = 8'h76 == io_state_in_11 ? 8'hb2 : _GEN_12149; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12151 = 8'h77 == io_state_in_11 ? 8'hbc : _GEN_12150; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12152 = 8'h78 == io_state_in_11 ? 8'he6 : _GEN_12151; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12153 = 8'h79 == io_state_in_11 ? 8'he8 : _GEN_12152; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12154 = 8'h7a == io_state_in_11 ? 8'hfa : _GEN_12153; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12155 = 8'h7b == io_state_in_11 ? 8'hf4 : _GEN_12154; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12156 = 8'h7c == io_state_in_11 ? 8'hde : _GEN_12155; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12157 = 8'h7d == io_state_in_11 ? 8'hd0 : _GEN_12156; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12158 = 8'h7e == io_state_in_11 ? 8'hc2 : _GEN_12157; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12159 = 8'h7f == io_state_in_11 ? 8'hcc : _GEN_12158; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12160 = 8'h80 == io_state_in_11 ? 8'h41 : _GEN_12159; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12161 = 8'h81 == io_state_in_11 ? 8'h4f : _GEN_12160; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12162 = 8'h82 == io_state_in_11 ? 8'h5d : _GEN_12161; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12163 = 8'h83 == io_state_in_11 ? 8'h53 : _GEN_12162; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12164 = 8'h84 == io_state_in_11 ? 8'h79 : _GEN_12163; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12165 = 8'h85 == io_state_in_11 ? 8'h77 : _GEN_12164; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12166 = 8'h86 == io_state_in_11 ? 8'h65 : _GEN_12165; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12167 = 8'h87 == io_state_in_11 ? 8'h6b : _GEN_12166; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12168 = 8'h88 == io_state_in_11 ? 8'h31 : _GEN_12167; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12169 = 8'h89 == io_state_in_11 ? 8'h3f : _GEN_12168; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12170 = 8'h8a == io_state_in_11 ? 8'h2d : _GEN_12169; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12171 = 8'h8b == io_state_in_11 ? 8'h23 : _GEN_12170; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12172 = 8'h8c == io_state_in_11 ? 8'h9 : _GEN_12171; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12173 = 8'h8d == io_state_in_11 ? 8'h7 : _GEN_12172; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12174 = 8'h8e == io_state_in_11 ? 8'h15 : _GEN_12173; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12175 = 8'h8f == io_state_in_11 ? 8'h1b : _GEN_12174; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12176 = 8'h90 == io_state_in_11 ? 8'ha1 : _GEN_12175; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12177 = 8'h91 == io_state_in_11 ? 8'haf : _GEN_12176; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12178 = 8'h92 == io_state_in_11 ? 8'hbd : _GEN_12177; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12179 = 8'h93 == io_state_in_11 ? 8'hb3 : _GEN_12178; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12180 = 8'h94 == io_state_in_11 ? 8'h99 : _GEN_12179; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12181 = 8'h95 == io_state_in_11 ? 8'h97 : _GEN_12180; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12182 = 8'h96 == io_state_in_11 ? 8'h85 : _GEN_12181; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12183 = 8'h97 == io_state_in_11 ? 8'h8b : _GEN_12182; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12184 = 8'h98 == io_state_in_11 ? 8'hd1 : _GEN_12183; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12185 = 8'h99 == io_state_in_11 ? 8'hdf : _GEN_12184; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12186 = 8'h9a == io_state_in_11 ? 8'hcd : _GEN_12185; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12187 = 8'h9b == io_state_in_11 ? 8'hc3 : _GEN_12186; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12188 = 8'h9c == io_state_in_11 ? 8'he9 : _GEN_12187; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12189 = 8'h9d == io_state_in_11 ? 8'he7 : _GEN_12188; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12190 = 8'h9e == io_state_in_11 ? 8'hf5 : _GEN_12189; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12191 = 8'h9f == io_state_in_11 ? 8'hfb : _GEN_12190; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12192 = 8'ha0 == io_state_in_11 ? 8'h9a : _GEN_12191; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12193 = 8'ha1 == io_state_in_11 ? 8'h94 : _GEN_12192; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12194 = 8'ha2 == io_state_in_11 ? 8'h86 : _GEN_12193; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12195 = 8'ha3 == io_state_in_11 ? 8'h88 : _GEN_12194; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12196 = 8'ha4 == io_state_in_11 ? 8'ha2 : _GEN_12195; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12197 = 8'ha5 == io_state_in_11 ? 8'hac : _GEN_12196; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12198 = 8'ha6 == io_state_in_11 ? 8'hbe : _GEN_12197; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12199 = 8'ha7 == io_state_in_11 ? 8'hb0 : _GEN_12198; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12200 = 8'ha8 == io_state_in_11 ? 8'hea : _GEN_12199; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12201 = 8'ha9 == io_state_in_11 ? 8'he4 : _GEN_12200; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12202 = 8'haa == io_state_in_11 ? 8'hf6 : _GEN_12201; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12203 = 8'hab == io_state_in_11 ? 8'hf8 : _GEN_12202; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12204 = 8'hac == io_state_in_11 ? 8'hd2 : _GEN_12203; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12205 = 8'had == io_state_in_11 ? 8'hdc : _GEN_12204; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12206 = 8'hae == io_state_in_11 ? 8'hce : _GEN_12205; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12207 = 8'haf == io_state_in_11 ? 8'hc0 : _GEN_12206; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12208 = 8'hb0 == io_state_in_11 ? 8'h7a : _GEN_12207; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12209 = 8'hb1 == io_state_in_11 ? 8'h74 : _GEN_12208; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12210 = 8'hb2 == io_state_in_11 ? 8'h66 : _GEN_12209; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12211 = 8'hb3 == io_state_in_11 ? 8'h68 : _GEN_12210; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12212 = 8'hb4 == io_state_in_11 ? 8'h42 : _GEN_12211; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12213 = 8'hb5 == io_state_in_11 ? 8'h4c : _GEN_12212; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12214 = 8'hb6 == io_state_in_11 ? 8'h5e : _GEN_12213; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12215 = 8'hb7 == io_state_in_11 ? 8'h50 : _GEN_12214; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12216 = 8'hb8 == io_state_in_11 ? 8'ha : _GEN_12215; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12217 = 8'hb9 == io_state_in_11 ? 8'h4 : _GEN_12216; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12218 = 8'hba == io_state_in_11 ? 8'h16 : _GEN_12217; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12219 = 8'hbb == io_state_in_11 ? 8'h18 : _GEN_12218; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12220 = 8'hbc == io_state_in_11 ? 8'h32 : _GEN_12219; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12221 = 8'hbd == io_state_in_11 ? 8'h3c : _GEN_12220; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12222 = 8'hbe == io_state_in_11 ? 8'h2e : _GEN_12221; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12223 = 8'hbf == io_state_in_11 ? 8'h20 : _GEN_12222; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12224 = 8'hc0 == io_state_in_11 ? 8'hec : _GEN_12223; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12225 = 8'hc1 == io_state_in_11 ? 8'he2 : _GEN_12224; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12226 = 8'hc2 == io_state_in_11 ? 8'hf0 : _GEN_12225; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12227 = 8'hc3 == io_state_in_11 ? 8'hfe : _GEN_12226; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12228 = 8'hc4 == io_state_in_11 ? 8'hd4 : _GEN_12227; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12229 = 8'hc5 == io_state_in_11 ? 8'hda : _GEN_12228; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12230 = 8'hc6 == io_state_in_11 ? 8'hc8 : _GEN_12229; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12231 = 8'hc7 == io_state_in_11 ? 8'hc6 : _GEN_12230; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12232 = 8'hc8 == io_state_in_11 ? 8'h9c : _GEN_12231; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12233 = 8'hc9 == io_state_in_11 ? 8'h92 : _GEN_12232; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12234 = 8'hca == io_state_in_11 ? 8'h80 : _GEN_12233; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12235 = 8'hcb == io_state_in_11 ? 8'h8e : _GEN_12234; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12236 = 8'hcc == io_state_in_11 ? 8'ha4 : _GEN_12235; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12237 = 8'hcd == io_state_in_11 ? 8'haa : _GEN_12236; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12238 = 8'hce == io_state_in_11 ? 8'hb8 : _GEN_12237; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12239 = 8'hcf == io_state_in_11 ? 8'hb6 : _GEN_12238; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12240 = 8'hd0 == io_state_in_11 ? 8'hc : _GEN_12239; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12241 = 8'hd1 == io_state_in_11 ? 8'h2 : _GEN_12240; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12242 = 8'hd2 == io_state_in_11 ? 8'h10 : _GEN_12241; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12243 = 8'hd3 == io_state_in_11 ? 8'h1e : _GEN_12242; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12244 = 8'hd4 == io_state_in_11 ? 8'h34 : _GEN_12243; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12245 = 8'hd5 == io_state_in_11 ? 8'h3a : _GEN_12244; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12246 = 8'hd6 == io_state_in_11 ? 8'h28 : _GEN_12245; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12247 = 8'hd7 == io_state_in_11 ? 8'h26 : _GEN_12246; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12248 = 8'hd8 == io_state_in_11 ? 8'h7c : _GEN_12247; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12249 = 8'hd9 == io_state_in_11 ? 8'h72 : _GEN_12248; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12250 = 8'hda == io_state_in_11 ? 8'h60 : _GEN_12249; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12251 = 8'hdb == io_state_in_11 ? 8'h6e : _GEN_12250; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12252 = 8'hdc == io_state_in_11 ? 8'h44 : _GEN_12251; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12253 = 8'hdd == io_state_in_11 ? 8'h4a : _GEN_12252; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12254 = 8'hde == io_state_in_11 ? 8'h58 : _GEN_12253; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12255 = 8'hdf == io_state_in_11 ? 8'h56 : _GEN_12254; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12256 = 8'he0 == io_state_in_11 ? 8'h37 : _GEN_12255; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12257 = 8'he1 == io_state_in_11 ? 8'h39 : _GEN_12256; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12258 = 8'he2 == io_state_in_11 ? 8'h2b : _GEN_12257; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12259 = 8'he3 == io_state_in_11 ? 8'h25 : _GEN_12258; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12260 = 8'he4 == io_state_in_11 ? 8'hf : _GEN_12259; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12261 = 8'he5 == io_state_in_11 ? 8'h1 : _GEN_12260; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12262 = 8'he6 == io_state_in_11 ? 8'h13 : _GEN_12261; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12263 = 8'he7 == io_state_in_11 ? 8'h1d : _GEN_12262; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12264 = 8'he8 == io_state_in_11 ? 8'h47 : _GEN_12263; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12265 = 8'he9 == io_state_in_11 ? 8'h49 : _GEN_12264; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12266 = 8'hea == io_state_in_11 ? 8'h5b : _GEN_12265; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12267 = 8'heb == io_state_in_11 ? 8'h55 : _GEN_12266; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12268 = 8'hec == io_state_in_11 ? 8'h7f : _GEN_12267; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12269 = 8'hed == io_state_in_11 ? 8'h71 : _GEN_12268; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12270 = 8'hee == io_state_in_11 ? 8'h63 : _GEN_12269; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12271 = 8'hef == io_state_in_11 ? 8'h6d : _GEN_12270; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12272 = 8'hf0 == io_state_in_11 ? 8'hd7 : _GEN_12271; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12273 = 8'hf1 == io_state_in_11 ? 8'hd9 : _GEN_12272; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12274 = 8'hf2 == io_state_in_11 ? 8'hcb : _GEN_12273; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12275 = 8'hf3 == io_state_in_11 ? 8'hc5 : _GEN_12274; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12276 = 8'hf4 == io_state_in_11 ? 8'hef : _GEN_12275; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12277 = 8'hf5 == io_state_in_11 ? 8'he1 : _GEN_12276; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12278 = 8'hf6 == io_state_in_11 ? 8'hf3 : _GEN_12277; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12279 = 8'hf7 == io_state_in_11 ? 8'hfd : _GEN_12278; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12280 = 8'hf8 == io_state_in_11 ? 8'ha7 : _GEN_12279; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12281 = 8'hf9 == io_state_in_11 ? 8'ha9 : _GEN_12280; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12282 = 8'hfa == io_state_in_11 ? 8'hbb : _GEN_12281; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12283 = 8'hfb == io_state_in_11 ? 8'hb5 : _GEN_12282; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12284 = 8'hfc == io_state_in_11 ? 8'h9f : _GEN_12283; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12285 = 8'hfd == io_state_in_11 ? 8'h91 : _GEN_12284; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12286 = 8'hfe == io_state_in_11 ? 8'h83 : _GEN_12285; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12287 = 8'hff == io_state_in_11 ? 8'h8d : _GEN_12286; // @[InvMixColumns.scala 139:{91,91}]
  wire [7:0] _GEN_12289 = 8'h1 == io_state_in_12 ? 8'he : 8'h0; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12290 = 8'h2 == io_state_in_12 ? 8'h1c : _GEN_12289; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12291 = 8'h3 == io_state_in_12 ? 8'h12 : _GEN_12290; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12292 = 8'h4 == io_state_in_12 ? 8'h38 : _GEN_12291; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12293 = 8'h5 == io_state_in_12 ? 8'h36 : _GEN_12292; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12294 = 8'h6 == io_state_in_12 ? 8'h24 : _GEN_12293; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12295 = 8'h7 == io_state_in_12 ? 8'h2a : _GEN_12294; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12296 = 8'h8 == io_state_in_12 ? 8'h70 : _GEN_12295; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12297 = 8'h9 == io_state_in_12 ? 8'h7e : _GEN_12296; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12298 = 8'ha == io_state_in_12 ? 8'h6c : _GEN_12297; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12299 = 8'hb == io_state_in_12 ? 8'h62 : _GEN_12298; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12300 = 8'hc == io_state_in_12 ? 8'h48 : _GEN_12299; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12301 = 8'hd == io_state_in_12 ? 8'h46 : _GEN_12300; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12302 = 8'he == io_state_in_12 ? 8'h54 : _GEN_12301; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12303 = 8'hf == io_state_in_12 ? 8'h5a : _GEN_12302; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12304 = 8'h10 == io_state_in_12 ? 8'he0 : _GEN_12303; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12305 = 8'h11 == io_state_in_12 ? 8'hee : _GEN_12304; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12306 = 8'h12 == io_state_in_12 ? 8'hfc : _GEN_12305; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12307 = 8'h13 == io_state_in_12 ? 8'hf2 : _GEN_12306; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12308 = 8'h14 == io_state_in_12 ? 8'hd8 : _GEN_12307; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12309 = 8'h15 == io_state_in_12 ? 8'hd6 : _GEN_12308; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12310 = 8'h16 == io_state_in_12 ? 8'hc4 : _GEN_12309; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12311 = 8'h17 == io_state_in_12 ? 8'hca : _GEN_12310; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12312 = 8'h18 == io_state_in_12 ? 8'h90 : _GEN_12311; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12313 = 8'h19 == io_state_in_12 ? 8'h9e : _GEN_12312; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12314 = 8'h1a == io_state_in_12 ? 8'h8c : _GEN_12313; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12315 = 8'h1b == io_state_in_12 ? 8'h82 : _GEN_12314; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12316 = 8'h1c == io_state_in_12 ? 8'ha8 : _GEN_12315; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12317 = 8'h1d == io_state_in_12 ? 8'ha6 : _GEN_12316; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12318 = 8'h1e == io_state_in_12 ? 8'hb4 : _GEN_12317; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12319 = 8'h1f == io_state_in_12 ? 8'hba : _GEN_12318; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12320 = 8'h20 == io_state_in_12 ? 8'hdb : _GEN_12319; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12321 = 8'h21 == io_state_in_12 ? 8'hd5 : _GEN_12320; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12322 = 8'h22 == io_state_in_12 ? 8'hc7 : _GEN_12321; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12323 = 8'h23 == io_state_in_12 ? 8'hc9 : _GEN_12322; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12324 = 8'h24 == io_state_in_12 ? 8'he3 : _GEN_12323; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12325 = 8'h25 == io_state_in_12 ? 8'hed : _GEN_12324; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12326 = 8'h26 == io_state_in_12 ? 8'hff : _GEN_12325; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12327 = 8'h27 == io_state_in_12 ? 8'hf1 : _GEN_12326; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12328 = 8'h28 == io_state_in_12 ? 8'hab : _GEN_12327; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12329 = 8'h29 == io_state_in_12 ? 8'ha5 : _GEN_12328; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12330 = 8'h2a == io_state_in_12 ? 8'hb7 : _GEN_12329; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12331 = 8'h2b == io_state_in_12 ? 8'hb9 : _GEN_12330; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12332 = 8'h2c == io_state_in_12 ? 8'h93 : _GEN_12331; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12333 = 8'h2d == io_state_in_12 ? 8'h9d : _GEN_12332; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12334 = 8'h2e == io_state_in_12 ? 8'h8f : _GEN_12333; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12335 = 8'h2f == io_state_in_12 ? 8'h81 : _GEN_12334; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12336 = 8'h30 == io_state_in_12 ? 8'h3b : _GEN_12335; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12337 = 8'h31 == io_state_in_12 ? 8'h35 : _GEN_12336; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12338 = 8'h32 == io_state_in_12 ? 8'h27 : _GEN_12337; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12339 = 8'h33 == io_state_in_12 ? 8'h29 : _GEN_12338; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12340 = 8'h34 == io_state_in_12 ? 8'h3 : _GEN_12339; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12341 = 8'h35 == io_state_in_12 ? 8'hd : _GEN_12340; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12342 = 8'h36 == io_state_in_12 ? 8'h1f : _GEN_12341; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12343 = 8'h37 == io_state_in_12 ? 8'h11 : _GEN_12342; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12344 = 8'h38 == io_state_in_12 ? 8'h4b : _GEN_12343; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12345 = 8'h39 == io_state_in_12 ? 8'h45 : _GEN_12344; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12346 = 8'h3a == io_state_in_12 ? 8'h57 : _GEN_12345; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12347 = 8'h3b == io_state_in_12 ? 8'h59 : _GEN_12346; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12348 = 8'h3c == io_state_in_12 ? 8'h73 : _GEN_12347; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12349 = 8'h3d == io_state_in_12 ? 8'h7d : _GEN_12348; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12350 = 8'h3e == io_state_in_12 ? 8'h6f : _GEN_12349; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12351 = 8'h3f == io_state_in_12 ? 8'h61 : _GEN_12350; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12352 = 8'h40 == io_state_in_12 ? 8'had : _GEN_12351; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12353 = 8'h41 == io_state_in_12 ? 8'ha3 : _GEN_12352; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12354 = 8'h42 == io_state_in_12 ? 8'hb1 : _GEN_12353; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12355 = 8'h43 == io_state_in_12 ? 8'hbf : _GEN_12354; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12356 = 8'h44 == io_state_in_12 ? 8'h95 : _GEN_12355; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12357 = 8'h45 == io_state_in_12 ? 8'h9b : _GEN_12356; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12358 = 8'h46 == io_state_in_12 ? 8'h89 : _GEN_12357; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12359 = 8'h47 == io_state_in_12 ? 8'h87 : _GEN_12358; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12360 = 8'h48 == io_state_in_12 ? 8'hdd : _GEN_12359; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12361 = 8'h49 == io_state_in_12 ? 8'hd3 : _GEN_12360; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12362 = 8'h4a == io_state_in_12 ? 8'hc1 : _GEN_12361; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12363 = 8'h4b == io_state_in_12 ? 8'hcf : _GEN_12362; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12364 = 8'h4c == io_state_in_12 ? 8'he5 : _GEN_12363; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12365 = 8'h4d == io_state_in_12 ? 8'heb : _GEN_12364; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12366 = 8'h4e == io_state_in_12 ? 8'hf9 : _GEN_12365; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12367 = 8'h4f == io_state_in_12 ? 8'hf7 : _GEN_12366; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12368 = 8'h50 == io_state_in_12 ? 8'h4d : _GEN_12367; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12369 = 8'h51 == io_state_in_12 ? 8'h43 : _GEN_12368; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12370 = 8'h52 == io_state_in_12 ? 8'h51 : _GEN_12369; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12371 = 8'h53 == io_state_in_12 ? 8'h5f : _GEN_12370; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12372 = 8'h54 == io_state_in_12 ? 8'h75 : _GEN_12371; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12373 = 8'h55 == io_state_in_12 ? 8'h7b : _GEN_12372; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12374 = 8'h56 == io_state_in_12 ? 8'h69 : _GEN_12373; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12375 = 8'h57 == io_state_in_12 ? 8'h67 : _GEN_12374; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12376 = 8'h58 == io_state_in_12 ? 8'h3d : _GEN_12375; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12377 = 8'h59 == io_state_in_12 ? 8'h33 : _GEN_12376; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12378 = 8'h5a == io_state_in_12 ? 8'h21 : _GEN_12377; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12379 = 8'h5b == io_state_in_12 ? 8'h2f : _GEN_12378; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12380 = 8'h5c == io_state_in_12 ? 8'h5 : _GEN_12379; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12381 = 8'h5d == io_state_in_12 ? 8'hb : _GEN_12380; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12382 = 8'h5e == io_state_in_12 ? 8'h19 : _GEN_12381; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12383 = 8'h5f == io_state_in_12 ? 8'h17 : _GEN_12382; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12384 = 8'h60 == io_state_in_12 ? 8'h76 : _GEN_12383; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12385 = 8'h61 == io_state_in_12 ? 8'h78 : _GEN_12384; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12386 = 8'h62 == io_state_in_12 ? 8'h6a : _GEN_12385; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12387 = 8'h63 == io_state_in_12 ? 8'h64 : _GEN_12386; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12388 = 8'h64 == io_state_in_12 ? 8'h4e : _GEN_12387; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12389 = 8'h65 == io_state_in_12 ? 8'h40 : _GEN_12388; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12390 = 8'h66 == io_state_in_12 ? 8'h52 : _GEN_12389; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12391 = 8'h67 == io_state_in_12 ? 8'h5c : _GEN_12390; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12392 = 8'h68 == io_state_in_12 ? 8'h6 : _GEN_12391; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12393 = 8'h69 == io_state_in_12 ? 8'h8 : _GEN_12392; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12394 = 8'h6a == io_state_in_12 ? 8'h1a : _GEN_12393; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12395 = 8'h6b == io_state_in_12 ? 8'h14 : _GEN_12394; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12396 = 8'h6c == io_state_in_12 ? 8'h3e : _GEN_12395; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12397 = 8'h6d == io_state_in_12 ? 8'h30 : _GEN_12396; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12398 = 8'h6e == io_state_in_12 ? 8'h22 : _GEN_12397; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12399 = 8'h6f == io_state_in_12 ? 8'h2c : _GEN_12398; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12400 = 8'h70 == io_state_in_12 ? 8'h96 : _GEN_12399; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12401 = 8'h71 == io_state_in_12 ? 8'h98 : _GEN_12400; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12402 = 8'h72 == io_state_in_12 ? 8'h8a : _GEN_12401; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12403 = 8'h73 == io_state_in_12 ? 8'h84 : _GEN_12402; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12404 = 8'h74 == io_state_in_12 ? 8'hae : _GEN_12403; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12405 = 8'h75 == io_state_in_12 ? 8'ha0 : _GEN_12404; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12406 = 8'h76 == io_state_in_12 ? 8'hb2 : _GEN_12405; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12407 = 8'h77 == io_state_in_12 ? 8'hbc : _GEN_12406; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12408 = 8'h78 == io_state_in_12 ? 8'he6 : _GEN_12407; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12409 = 8'h79 == io_state_in_12 ? 8'he8 : _GEN_12408; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12410 = 8'h7a == io_state_in_12 ? 8'hfa : _GEN_12409; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12411 = 8'h7b == io_state_in_12 ? 8'hf4 : _GEN_12410; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12412 = 8'h7c == io_state_in_12 ? 8'hde : _GEN_12411; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12413 = 8'h7d == io_state_in_12 ? 8'hd0 : _GEN_12412; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12414 = 8'h7e == io_state_in_12 ? 8'hc2 : _GEN_12413; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12415 = 8'h7f == io_state_in_12 ? 8'hcc : _GEN_12414; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12416 = 8'h80 == io_state_in_12 ? 8'h41 : _GEN_12415; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12417 = 8'h81 == io_state_in_12 ? 8'h4f : _GEN_12416; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12418 = 8'h82 == io_state_in_12 ? 8'h5d : _GEN_12417; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12419 = 8'h83 == io_state_in_12 ? 8'h53 : _GEN_12418; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12420 = 8'h84 == io_state_in_12 ? 8'h79 : _GEN_12419; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12421 = 8'h85 == io_state_in_12 ? 8'h77 : _GEN_12420; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12422 = 8'h86 == io_state_in_12 ? 8'h65 : _GEN_12421; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12423 = 8'h87 == io_state_in_12 ? 8'h6b : _GEN_12422; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12424 = 8'h88 == io_state_in_12 ? 8'h31 : _GEN_12423; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12425 = 8'h89 == io_state_in_12 ? 8'h3f : _GEN_12424; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12426 = 8'h8a == io_state_in_12 ? 8'h2d : _GEN_12425; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12427 = 8'h8b == io_state_in_12 ? 8'h23 : _GEN_12426; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12428 = 8'h8c == io_state_in_12 ? 8'h9 : _GEN_12427; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12429 = 8'h8d == io_state_in_12 ? 8'h7 : _GEN_12428; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12430 = 8'h8e == io_state_in_12 ? 8'h15 : _GEN_12429; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12431 = 8'h8f == io_state_in_12 ? 8'h1b : _GEN_12430; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12432 = 8'h90 == io_state_in_12 ? 8'ha1 : _GEN_12431; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12433 = 8'h91 == io_state_in_12 ? 8'haf : _GEN_12432; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12434 = 8'h92 == io_state_in_12 ? 8'hbd : _GEN_12433; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12435 = 8'h93 == io_state_in_12 ? 8'hb3 : _GEN_12434; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12436 = 8'h94 == io_state_in_12 ? 8'h99 : _GEN_12435; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12437 = 8'h95 == io_state_in_12 ? 8'h97 : _GEN_12436; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12438 = 8'h96 == io_state_in_12 ? 8'h85 : _GEN_12437; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12439 = 8'h97 == io_state_in_12 ? 8'h8b : _GEN_12438; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12440 = 8'h98 == io_state_in_12 ? 8'hd1 : _GEN_12439; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12441 = 8'h99 == io_state_in_12 ? 8'hdf : _GEN_12440; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12442 = 8'h9a == io_state_in_12 ? 8'hcd : _GEN_12441; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12443 = 8'h9b == io_state_in_12 ? 8'hc3 : _GEN_12442; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12444 = 8'h9c == io_state_in_12 ? 8'he9 : _GEN_12443; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12445 = 8'h9d == io_state_in_12 ? 8'he7 : _GEN_12444; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12446 = 8'h9e == io_state_in_12 ? 8'hf5 : _GEN_12445; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12447 = 8'h9f == io_state_in_12 ? 8'hfb : _GEN_12446; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12448 = 8'ha0 == io_state_in_12 ? 8'h9a : _GEN_12447; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12449 = 8'ha1 == io_state_in_12 ? 8'h94 : _GEN_12448; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12450 = 8'ha2 == io_state_in_12 ? 8'h86 : _GEN_12449; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12451 = 8'ha3 == io_state_in_12 ? 8'h88 : _GEN_12450; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12452 = 8'ha4 == io_state_in_12 ? 8'ha2 : _GEN_12451; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12453 = 8'ha5 == io_state_in_12 ? 8'hac : _GEN_12452; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12454 = 8'ha6 == io_state_in_12 ? 8'hbe : _GEN_12453; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12455 = 8'ha7 == io_state_in_12 ? 8'hb0 : _GEN_12454; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12456 = 8'ha8 == io_state_in_12 ? 8'hea : _GEN_12455; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12457 = 8'ha9 == io_state_in_12 ? 8'he4 : _GEN_12456; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12458 = 8'haa == io_state_in_12 ? 8'hf6 : _GEN_12457; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12459 = 8'hab == io_state_in_12 ? 8'hf8 : _GEN_12458; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12460 = 8'hac == io_state_in_12 ? 8'hd2 : _GEN_12459; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12461 = 8'had == io_state_in_12 ? 8'hdc : _GEN_12460; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12462 = 8'hae == io_state_in_12 ? 8'hce : _GEN_12461; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12463 = 8'haf == io_state_in_12 ? 8'hc0 : _GEN_12462; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12464 = 8'hb0 == io_state_in_12 ? 8'h7a : _GEN_12463; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12465 = 8'hb1 == io_state_in_12 ? 8'h74 : _GEN_12464; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12466 = 8'hb2 == io_state_in_12 ? 8'h66 : _GEN_12465; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12467 = 8'hb3 == io_state_in_12 ? 8'h68 : _GEN_12466; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12468 = 8'hb4 == io_state_in_12 ? 8'h42 : _GEN_12467; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12469 = 8'hb5 == io_state_in_12 ? 8'h4c : _GEN_12468; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12470 = 8'hb6 == io_state_in_12 ? 8'h5e : _GEN_12469; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12471 = 8'hb7 == io_state_in_12 ? 8'h50 : _GEN_12470; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12472 = 8'hb8 == io_state_in_12 ? 8'ha : _GEN_12471; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12473 = 8'hb9 == io_state_in_12 ? 8'h4 : _GEN_12472; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12474 = 8'hba == io_state_in_12 ? 8'h16 : _GEN_12473; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12475 = 8'hbb == io_state_in_12 ? 8'h18 : _GEN_12474; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12476 = 8'hbc == io_state_in_12 ? 8'h32 : _GEN_12475; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12477 = 8'hbd == io_state_in_12 ? 8'h3c : _GEN_12476; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12478 = 8'hbe == io_state_in_12 ? 8'h2e : _GEN_12477; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12479 = 8'hbf == io_state_in_12 ? 8'h20 : _GEN_12478; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12480 = 8'hc0 == io_state_in_12 ? 8'hec : _GEN_12479; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12481 = 8'hc1 == io_state_in_12 ? 8'he2 : _GEN_12480; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12482 = 8'hc2 == io_state_in_12 ? 8'hf0 : _GEN_12481; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12483 = 8'hc3 == io_state_in_12 ? 8'hfe : _GEN_12482; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12484 = 8'hc4 == io_state_in_12 ? 8'hd4 : _GEN_12483; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12485 = 8'hc5 == io_state_in_12 ? 8'hda : _GEN_12484; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12486 = 8'hc6 == io_state_in_12 ? 8'hc8 : _GEN_12485; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12487 = 8'hc7 == io_state_in_12 ? 8'hc6 : _GEN_12486; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12488 = 8'hc8 == io_state_in_12 ? 8'h9c : _GEN_12487; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12489 = 8'hc9 == io_state_in_12 ? 8'h92 : _GEN_12488; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12490 = 8'hca == io_state_in_12 ? 8'h80 : _GEN_12489; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12491 = 8'hcb == io_state_in_12 ? 8'h8e : _GEN_12490; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12492 = 8'hcc == io_state_in_12 ? 8'ha4 : _GEN_12491; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12493 = 8'hcd == io_state_in_12 ? 8'haa : _GEN_12492; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12494 = 8'hce == io_state_in_12 ? 8'hb8 : _GEN_12493; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12495 = 8'hcf == io_state_in_12 ? 8'hb6 : _GEN_12494; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12496 = 8'hd0 == io_state_in_12 ? 8'hc : _GEN_12495; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12497 = 8'hd1 == io_state_in_12 ? 8'h2 : _GEN_12496; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12498 = 8'hd2 == io_state_in_12 ? 8'h10 : _GEN_12497; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12499 = 8'hd3 == io_state_in_12 ? 8'h1e : _GEN_12498; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12500 = 8'hd4 == io_state_in_12 ? 8'h34 : _GEN_12499; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12501 = 8'hd5 == io_state_in_12 ? 8'h3a : _GEN_12500; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12502 = 8'hd6 == io_state_in_12 ? 8'h28 : _GEN_12501; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12503 = 8'hd7 == io_state_in_12 ? 8'h26 : _GEN_12502; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12504 = 8'hd8 == io_state_in_12 ? 8'h7c : _GEN_12503; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12505 = 8'hd9 == io_state_in_12 ? 8'h72 : _GEN_12504; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12506 = 8'hda == io_state_in_12 ? 8'h60 : _GEN_12505; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12507 = 8'hdb == io_state_in_12 ? 8'h6e : _GEN_12506; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12508 = 8'hdc == io_state_in_12 ? 8'h44 : _GEN_12507; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12509 = 8'hdd == io_state_in_12 ? 8'h4a : _GEN_12508; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12510 = 8'hde == io_state_in_12 ? 8'h58 : _GEN_12509; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12511 = 8'hdf == io_state_in_12 ? 8'h56 : _GEN_12510; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12512 = 8'he0 == io_state_in_12 ? 8'h37 : _GEN_12511; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12513 = 8'he1 == io_state_in_12 ? 8'h39 : _GEN_12512; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12514 = 8'he2 == io_state_in_12 ? 8'h2b : _GEN_12513; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12515 = 8'he3 == io_state_in_12 ? 8'h25 : _GEN_12514; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12516 = 8'he4 == io_state_in_12 ? 8'hf : _GEN_12515; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12517 = 8'he5 == io_state_in_12 ? 8'h1 : _GEN_12516; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12518 = 8'he6 == io_state_in_12 ? 8'h13 : _GEN_12517; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12519 = 8'he7 == io_state_in_12 ? 8'h1d : _GEN_12518; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12520 = 8'he8 == io_state_in_12 ? 8'h47 : _GEN_12519; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12521 = 8'he9 == io_state_in_12 ? 8'h49 : _GEN_12520; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12522 = 8'hea == io_state_in_12 ? 8'h5b : _GEN_12521; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12523 = 8'heb == io_state_in_12 ? 8'h55 : _GEN_12522; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12524 = 8'hec == io_state_in_12 ? 8'h7f : _GEN_12523; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12525 = 8'hed == io_state_in_12 ? 8'h71 : _GEN_12524; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12526 = 8'hee == io_state_in_12 ? 8'h63 : _GEN_12525; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12527 = 8'hef == io_state_in_12 ? 8'h6d : _GEN_12526; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12528 = 8'hf0 == io_state_in_12 ? 8'hd7 : _GEN_12527; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12529 = 8'hf1 == io_state_in_12 ? 8'hd9 : _GEN_12528; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12530 = 8'hf2 == io_state_in_12 ? 8'hcb : _GEN_12529; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12531 = 8'hf3 == io_state_in_12 ? 8'hc5 : _GEN_12530; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12532 = 8'hf4 == io_state_in_12 ? 8'hef : _GEN_12531; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12533 = 8'hf5 == io_state_in_12 ? 8'he1 : _GEN_12532; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12534 = 8'hf6 == io_state_in_12 ? 8'hf3 : _GEN_12533; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12535 = 8'hf7 == io_state_in_12 ? 8'hfd : _GEN_12534; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12536 = 8'hf8 == io_state_in_12 ? 8'ha7 : _GEN_12535; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12537 = 8'hf9 == io_state_in_12 ? 8'ha9 : _GEN_12536; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12538 = 8'hfa == io_state_in_12 ? 8'hbb : _GEN_12537; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12539 = 8'hfb == io_state_in_12 ? 8'hb5 : _GEN_12538; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12540 = 8'hfc == io_state_in_12 ? 8'h9f : _GEN_12539; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12541 = 8'hfd == io_state_in_12 ? 8'h91 : _GEN_12540; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12542 = 8'hfe == io_state_in_12 ? 8'h83 : _GEN_12541; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12543 = 8'hff == io_state_in_12 ? 8'h8d : _GEN_12542; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12545 = 8'h1 == io_state_in_13 ? 8'hb : 8'h0; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12546 = 8'h2 == io_state_in_13 ? 8'h16 : _GEN_12545; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12547 = 8'h3 == io_state_in_13 ? 8'h1d : _GEN_12546; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12548 = 8'h4 == io_state_in_13 ? 8'h2c : _GEN_12547; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12549 = 8'h5 == io_state_in_13 ? 8'h27 : _GEN_12548; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12550 = 8'h6 == io_state_in_13 ? 8'h3a : _GEN_12549; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12551 = 8'h7 == io_state_in_13 ? 8'h31 : _GEN_12550; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12552 = 8'h8 == io_state_in_13 ? 8'h58 : _GEN_12551; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12553 = 8'h9 == io_state_in_13 ? 8'h53 : _GEN_12552; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12554 = 8'ha == io_state_in_13 ? 8'h4e : _GEN_12553; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12555 = 8'hb == io_state_in_13 ? 8'h45 : _GEN_12554; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12556 = 8'hc == io_state_in_13 ? 8'h74 : _GEN_12555; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12557 = 8'hd == io_state_in_13 ? 8'h7f : _GEN_12556; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12558 = 8'he == io_state_in_13 ? 8'h62 : _GEN_12557; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12559 = 8'hf == io_state_in_13 ? 8'h69 : _GEN_12558; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12560 = 8'h10 == io_state_in_13 ? 8'hb0 : _GEN_12559; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12561 = 8'h11 == io_state_in_13 ? 8'hbb : _GEN_12560; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12562 = 8'h12 == io_state_in_13 ? 8'ha6 : _GEN_12561; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12563 = 8'h13 == io_state_in_13 ? 8'had : _GEN_12562; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12564 = 8'h14 == io_state_in_13 ? 8'h9c : _GEN_12563; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12565 = 8'h15 == io_state_in_13 ? 8'h97 : _GEN_12564; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12566 = 8'h16 == io_state_in_13 ? 8'h8a : _GEN_12565; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12567 = 8'h17 == io_state_in_13 ? 8'h81 : _GEN_12566; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12568 = 8'h18 == io_state_in_13 ? 8'he8 : _GEN_12567; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12569 = 8'h19 == io_state_in_13 ? 8'he3 : _GEN_12568; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12570 = 8'h1a == io_state_in_13 ? 8'hfe : _GEN_12569; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12571 = 8'h1b == io_state_in_13 ? 8'hf5 : _GEN_12570; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12572 = 8'h1c == io_state_in_13 ? 8'hc4 : _GEN_12571; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12573 = 8'h1d == io_state_in_13 ? 8'hcf : _GEN_12572; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12574 = 8'h1e == io_state_in_13 ? 8'hd2 : _GEN_12573; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12575 = 8'h1f == io_state_in_13 ? 8'hd9 : _GEN_12574; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12576 = 8'h20 == io_state_in_13 ? 8'h7b : _GEN_12575; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12577 = 8'h21 == io_state_in_13 ? 8'h70 : _GEN_12576; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12578 = 8'h22 == io_state_in_13 ? 8'h6d : _GEN_12577; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12579 = 8'h23 == io_state_in_13 ? 8'h66 : _GEN_12578; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12580 = 8'h24 == io_state_in_13 ? 8'h57 : _GEN_12579; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12581 = 8'h25 == io_state_in_13 ? 8'h5c : _GEN_12580; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12582 = 8'h26 == io_state_in_13 ? 8'h41 : _GEN_12581; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12583 = 8'h27 == io_state_in_13 ? 8'h4a : _GEN_12582; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12584 = 8'h28 == io_state_in_13 ? 8'h23 : _GEN_12583; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12585 = 8'h29 == io_state_in_13 ? 8'h28 : _GEN_12584; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12586 = 8'h2a == io_state_in_13 ? 8'h35 : _GEN_12585; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12587 = 8'h2b == io_state_in_13 ? 8'h3e : _GEN_12586; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12588 = 8'h2c == io_state_in_13 ? 8'hf : _GEN_12587; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12589 = 8'h2d == io_state_in_13 ? 8'h4 : _GEN_12588; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12590 = 8'h2e == io_state_in_13 ? 8'h19 : _GEN_12589; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12591 = 8'h2f == io_state_in_13 ? 8'h12 : _GEN_12590; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12592 = 8'h30 == io_state_in_13 ? 8'hcb : _GEN_12591; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12593 = 8'h31 == io_state_in_13 ? 8'hc0 : _GEN_12592; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12594 = 8'h32 == io_state_in_13 ? 8'hdd : _GEN_12593; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12595 = 8'h33 == io_state_in_13 ? 8'hd6 : _GEN_12594; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12596 = 8'h34 == io_state_in_13 ? 8'he7 : _GEN_12595; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12597 = 8'h35 == io_state_in_13 ? 8'hec : _GEN_12596; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12598 = 8'h36 == io_state_in_13 ? 8'hf1 : _GEN_12597; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12599 = 8'h37 == io_state_in_13 ? 8'hfa : _GEN_12598; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12600 = 8'h38 == io_state_in_13 ? 8'h93 : _GEN_12599; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12601 = 8'h39 == io_state_in_13 ? 8'h98 : _GEN_12600; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12602 = 8'h3a == io_state_in_13 ? 8'h85 : _GEN_12601; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12603 = 8'h3b == io_state_in_13 ? 8'h8e : _GEN_12602; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12604 = 8'h3c == io_state_in_13 ? 8'hbf : _GEN_12603; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12605 = 8'h3d == io_state_in_13 ? 8'hb4 : _GEN_12604; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12606 = 8'h3e == io_state_in_13 ? 8'ha9 : _GEN_12605; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12607 = 8'h3f == io_state_in_13 ? 8'ha2 : _GEN_12606; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12608 = 8'h40 == io_state_in_13 ? 8'hf6 : _GEN_12607; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12609 = 8'h41 == io_state_in_13 ? 8'hfd : _GEN_12608; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12610 = 8'h42 == io_state_in_13 ? 8'he0 : _GEN_12609; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12611 = 8'h43 == io_state_in_13 ? 8'heb : _GEN_12610; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12612 = 8'h44 == io_state_in_13 ? 8'hda : _GEN_12611; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12613 = 8'h45 == io_state_in_13 ? 8'hd1 : _GEN_12612; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12614 = 8'h46 == io_state_in_13 ? 8'hcc : _GEN_12613; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12615 = 8'h47 == io_state_in_13 ? 8'hc7 : _GEN_12614; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12616 = 8'h48 == io_state_in_13 ? 8'hae : _GEN_12615; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12617 = 8'h49 == io_state_in_13 ? 8'ha5 : _GEN_12616; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12618 = 8'h4a == io_state_in_13 ? 8'hb8 : _GEN_12617; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12619 = 8'h4b == io_state_in_13 ? 8'hb3 : _GEN_12618; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12620 = 8'h4c == io_state_in_13 ? 8'h82 : _GEN_12619; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12621 = 8'h4d == io_state_in_13 ? 8'h89 : _GEN_12620; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12622 = 8'h4e == io_state_in_13 ? 8'h94 : _GEN_12621; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12623 = 8'h4f == io_state_in_13 ? 8'h9f : _GEN_12622; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12624 = 8'h50 == io_state_in_13 ? 8'h46 : _GEN_12623; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12625 = 8'h51 == io_state_in_13 ? 8'h4d : _GEN_12624; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12626 = 8'h52 == io_state_in_13 ? 8'h50 : _GEN_12625; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12627 = 8'h53 == io_state_in_13 ? 8'h5b : _GEN_12626; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12628 = 8'h54 == io_state_in_13 ? 8'h6a : _GEN_12627; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12629 = 8'h55 == io_state_in_13 ? 8'h61 : _GEN_12628; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12630 = 8'h56 == io_state_in_13 ? 8'h7c : _GEN_12629; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12631 = 8'h57 == io_state_in_13 ? 8'h77 : _GEN_12630; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12632 = 8'h58 == io_state_in_13 ? 8'h1e : _GEN_12631; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12633 = 8'h59 == io_state_in_13 ? 8'h15 : _GEN_12632; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12634 = 8'h5a == io_state_in_13 ? 8'h8 : _GEN_12633; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12635 = 8'h5b == io_state_in_13 ? 8'h3 : _GEN_12634; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12636 = 8'h5c == io_state_in_13 ? 8'h32 : _GEN_12635; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12637 = 8'h5d == io_state_in_13 ? 8'h39 : _GEN_12636; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12638 = 8'h5e == io_state_in_13 ? 8'h24 : _GEN_12637; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12639 = 8'h5f == io_state_in_13 ? 8'h2f : _GEN_12638; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12640 = 8'h60 == io_state_in_13 ? 8'h8d : _GEN_12639; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12641 = 8'h61 == io_state_in_13 ? 8'h86 : _GEN_12640; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12642 = 8'h62 == io_state_in_13 ? 8'h9b : _GEN_12641; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12643 = 8'h63 == io_state_in_13 ? 8'h90 : _GEN_12642; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12644 = 8'h64 == io_state_in_13 ? 8'ha1 : _GEN_12643; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12645 = 8'h65 == io_state_in_13 ? 8'haa : _GEN_12644; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12646 = 8'h66 == io_state_in_13 ? 8'hb7 : _GEN_12645; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12647 = 8'h67 == io_state_in_13 ? 8'hbc : _GEN_12646; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12648 = 8'h68 == io_state_in_13 ? 8'hd5 : _GEN_12647; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12649 = 8'h69 == io_state_in_13 ? 8'hde : _GEN_12648; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12650 = 8'h6a == io_state_in_13 ? 8'hc3 : _GEN_12649; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12651 = 8'h6b == io_state_in_13 ? 8'hc8 : _GEN_12650; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12652 = 8'h6c == io_state_in_13 ? 8'hf9 : _GEN_12651; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12653 = 8'h6d == io_state_in_13 ? 8'hf2 : _GEN_12652; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12654 = 8'h6e == io_state_in_13 ? 8'hef : _GEN_12653; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12655 = 8'h6f == io_state_in_13 ? 8'he4 : _GEN_12654; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12656 = 8'h70 == io_state_in_13 ? 8'h3d : _GEN_12655; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12657 = 8'h71 == io_state_in_13 ? 8'h36 : _GEN_12656; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12658 = 8'h72 == io_state_in_13 ? 8'h2b : _GEN_12657; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12659 = 8'h73 == io_state_in_13 ? 8'h20 : _GEN_12658; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12660 = 8'h74 == io_state_in_13 ? 8'h11 : _GEN_12659; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12661 = 8'h75 == io_state_in_13 ? 8'h1a : _GEN_12660; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12662 = 8'h76 == io_state_in_13 ? 8'h7 : _GEN_12661; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12663 = 8'h77 == io_state_in_13 ? 8'hc : _GEN_12662; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12664 = 8'h78 == io_state_in_13 ? 8'h65 : _GEN_12663; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12665 = 8'h79 == io_state_in_13 ? 8'h6e : _GEN_12664; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12666 = 8'h7a == io_state_in_13 ? 8'h73 : _GEN_12665; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12667 = 8'h7b == io_state_in_13 ? 8'h78 : _GEN_12666; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12668 = 8'h7c == io_state_in_13 ? 8'h49 : _GEN_12667; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12669 = 8'h7d == io_state_in_13 ? 8'h42 : _GEN_12668; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12670 = 8'h7e == io_state_in_13 ? 8'h5f : _GEN_12669; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12671 = 8'h7f == io_state_in_13 ? 8'h54 : _GEN_12670; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12672 = 8'h80 == io_state_in_13 ? 8'hf7 : _GEN_12671; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12673 = 8'h81 == io_state_in_13 ? 8'hfc : _GEN_12672; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12674 = 8'h82 == io_state_in_13 ? 8'he1 : _GEN_12673; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12675 = 8'h83 == io_state_in_13 ? 8'hea : _GEN_12674; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12676 = 8'h84 == io_state_in_13 ? 8'hdb : _GEN_12675; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12677 = 8'h85 == io_state_in_13 ? 8'hd0 : _GEN_12676; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12678 = 8'h86 == io_state_in_13 ? 8'hcd : _GEN_12677; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12679 = 8'h87 == io_state_in_13 ? 8'hc6 : _GEN_12678; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12680 = 8'h88 == io_state_in_13 ? 8'haf : _GEN_12679; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12681 = 8'h89 == io_state_in_13 ? 8'ha4 : _GEN_12680; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12682 = 8'h8a == io_state_in_13 ? 8'hb9 : _GEN_12681; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12683 = 8'h8b == io_state_in_13 ? 8'hb2 : _GEN_12682; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12684 = 8'h8c == io_state_in_13 ? 8'h83 : _GEN_12683; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12685 = 8'h8d == io_state_in_13 ? 8'h88 : _GEN_12684; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12686 = 8'h8e == io_state_in_13 ? 8'h95 : _GEN_12685; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12687 = 8'h8f == io_state_in_13 ? 8'h9e : _GEN_12686; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12688 = 8'h90 == io_state_in_13 ? 8'h47 : _GEN_12687; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12689 = 8'h91 == io_state_in_13 ? 8'h4c : _GEN_12688; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12690 = 8'h92 == io_state_in_13 ? 8'h51 : _GEN_12689; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12691 = 8'h93 == io_state_in_13 ? 8'h5a : _GEN_12690; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12692 = 8'h94 == io_state_in_13 ? 8'h6b : _GEN_12691; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12693 = 8'h95 == io_state_in_13 ? 8'h60 : _GEN_12692; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12694 = 8'h96 == io_state_in_13 ? 8'h7d : _GEN_12693; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12695 = 8'h97 == io_state_in_13 ? 8'h76 : _GEN_12694; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12696 = 8'h98 == io_state_in_13 ? 8'h1f : _GEN_12695; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12697 = 8'h99 == io_state_in_13 ? 8'h14 : _GEN_12696; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12698 = 8'h9a == io_state_in_13 ? 8'h9 : _GEN_12697; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12699 = 8'h9b == io_state_in_13 ? 8'h2 : _GEN_12698; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12700 = 8'h9c == io_state_in_13 ? 8'h33 : _GEN_12699; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12701 = 8'h9d == io_state_in_13 ? 8'h38 : _GEN_12700; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12702 = 8'h9e == io_state_in_13 ? 8'h25 : _GEN_12701; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12703 = 8'h9f == io_state_in_13 ? 8'h2e : _GEN_12702; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12704 = 8'ha0 == io_state_in_13 ? 8'h8c : _GEN_12703; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12705 = 8'ha1 == io_state_in_13 ? 8'h87 : _GEN_12704; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12706 = 8'ha2 == io_state_in_13 ? 8'h9a : _GEN_12705; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12707 = 8'ha3 == io_state_in_13 ? 8'h91 : _GEN_12706; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12708 = 8'ha4 == io_state_in_13 ? 8'ha0 : _GEN_12707; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12709 = 8'ha5 == io_state_in_13 ? 8'hab : _GEN_12708; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12710 = 8'ha6 == io_state_in_13 ? 8'hb6 : _GEN_12709; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12711 = 8'ha7 == io_state_in_13 ? 8'hbd : _GEN_12710; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12712 = 8'ha8 == io_state_in_13 ? 8'hd4 : _GEN_12711; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12713 = 8'ha9 == io_state_in_13 ? 8'hdf : _GEN_12712; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12714 = 8'haa == io_state_in_13 ? 8'hc2 : _GEN_12713; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12715 = 8'hab == io_state_in_13 ? 8'hc9 : _GEN_12714; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12716 = 8'hac == io_state_in_13 ? 8'hf8 : _GEN_12715; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12717 = 8'had == io_state_in_13 ? 8'hf3 : _GEN_12716; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12718 = 8'hae == io_state_in_13 ? 8'hee : _GEN_12717; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12719 = 8'haf == io_state_in_13 ? 8'he5 : _GEN_12718; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12720 = 8'hb0 == io_state_in_13 ? 8'h3c : _GEN_12719; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12721 = 8'hb1 == io_state_in_13 ? 8'h37 : _GEN_12720; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12722 = 8'hb2 == io_state_in_13 ? 8'h2a : _GEN_12721; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12723 = 8'hb3 == io_state_in_13 ? 8'h21 : _GEN_12722; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12724 = 8'hb4 == io_state_in_13 ? 8'h10 : _GEN_12723; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12725 = 8'hb5 == io_state_in_13 ? 8'h1b : _GEN_12724; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12726 = 8'hb6 == io_state_in_13 ? 8'h6 : _GEN_12725; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12727 = 8'hb7 == io_state_in_13 ? 8'hd : _GEN_12726; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12728 = 8'hb8 == io_state_in_13 ? 8'h64 : _GEN_12727; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12729 = 8'hb9 == io_state_in_13 ? 8'h6f : _GEN_12728; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12730 = 8'hba == io_state_in_13 ? 8'h72 : _GEN_12729; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12731 = 8'hbb == io_state_in_13 ? 8'h79 : _GEN_12730; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12732 = 8'hbc == io_state_in_13 ? 8'h48 : _GEN_12731; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12733 = 8'hbd == io_state_in_13 ? 8'h43 : _GEN_12732; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12734 = 8'hbe == io_state_in_13 ? 8'h5e : _GEN_12733; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12735 = 8'hbf == io_state_in_13 ? 8'h55 : _GEN_12734; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12736 = 8'hc0 == io_state_in_13 ? 8'h1 : _GEN_12735; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12737 = 8'hc1 == io_state_in_13 ? 8'ha : _GEN_12736; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12738 = 8'hc2 == io_state_in_13 ? 8'h17 : _GEN_12737; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12739 = 8'hc3 == io_state_in_13 ? 8'h1c : _GEN_12738; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12740 = 8'hc4 == io_state_in_13 ? 8'h2d : _GEN_12739; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12741 = 8'hc5 == io_state_in_13 ? 8'h26 : _GEN_12740; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12742 = 8'hc6 == io_state_in_13 ? 8'h3b : _GEN_12741; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12743 = 8'hc7 == io_state_in_13 ? 8'h30 : _GEN_12742; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12744 = 8'hc8 == io_state_in_13 ? 8'h59 : _GEN_12743; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12745 = 8'hc9 == io_state_in_13 ? 8'h52 : _GEN_12744; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12746 = 8'hca == io_state_in_13 ? 8'h4f : _GEN_12745; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12747 = 8'hcb == io_state_in_13 ? 8'h44 : _GEN_12746; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12748 = 8'hcc == io_state_in_13 ? 8'h75 : _GEN_12747; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12749 = 8'hcd == io_state_in_13 ? 8'h7e : _GEN_12748; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12750 = 8'hce == io_state_in_13 ? 8'h63 : _GEN_12749; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12751 = 8'hcf == io_state_in_13 ? 8'h68 : _GEN_12750; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12752 = 8'hd0 == io_state_in_13 ? 8'hb1 : _GEN_12751; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12753 = 8'hd1 == io_state_in_13 ? 8'hba : _GEN_12752; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12754 = 8'hd2 == io_state_in_13 ? 8'ha7 : _GEN_12753; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12755 = 8'hd3 == io_state_in_13 ? 8'hac : _GEN_12754; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12756 = 8'hd4 == io_state_in_13 ? 8'h9d : _GEN_12755; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12757 = 8'hd5 == io_state_in_13 ? 8'h96 : _GEN_12756; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12758 = 8'hd6 == io_state_in_13 ? 8'h8b : _GEN_12757; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12759 = 8'hd7 == io_state_in_13 ? 8'h80 : _GEN_12758; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12760 = 8'hd8 == io_state_in_13 ? 8'he9 : _GEN_12759; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12761 = 8'hd9 == io_state_in_13 ? 8'he2 : _GEN_12760; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12762 = 8'hda == io_state_in_13 ? 8'hff : _GEN_12761; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12763 = 8'hdb == io_state_in_13 ? 8'hf4 : _GEN_12762; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12764 = 8'hdc == io_state_in_13 ? 8'hc5 : _GEN_12763; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12765 = 8'hdd == io_state_in_13 ? 8'hce : _GEN_12764; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12766 = 8'hde == io_state_in_13 ? 8'hd3 : _GEN_12765; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12767 = 8'hdf == io_state_in_13 ? 8'hd8 : _GEN_12766; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12768 = 8'he0 == io_state_in_13 ? 8'h7a : _GEN_12767; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12769 = 8'he1 == io_state_in_13 ? 8'h71 : _GEN_12768; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12770 = 8'he2 == io_state_in_13 ? 8'h6c : _GEN_12769; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12771 = 8'he3 == io_state_in_13 ? 8'h67 : _GEN_12770; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12772 = 8'he4 == io_state_in_13 ? 8'h56 : _GEN_12771; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12773 = 8'he5 == io_state_in_13 ? 8'h5d : _GEN_12772; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12774 = 8'he6 == io_state_in_13 ? 8'h40 : _GEN_12773; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12775 = 8'he7 == io_state_in_13 ? 8'h4b : _GEN_12774; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12776 = 8'he8 == io_state_in_13 ? 8'h22 : _GEN_12775; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12777 = 8'he9 == io_state_in_13 ? 8'h29 : _GEN_12776; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12778 = 8'hea == io_state_in_13 ? 8'h34 : _GEN_12777; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12779 = 8'heb == io_state_in_13 ? 8'h3f : _GEN_12778; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12780 = 8'hec == io_state_in_13 ? 8'he : _GEN_12779; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12781 = 8'hed == io_state_in_13 ? 8'h5 : _GEN_12780; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12782 = 8'hee == io_state_in_13 ? 8'h18 : _GEN_12781; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12783 = 8'hef == io_state_in_13 ? 8'h13 : _GEN_12782; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12784 = 8'hf0 == io_state_in_13 ? 8'hca : _GEN_12783; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12785 = 8'hf1 == io_state_in_13 ? 8'hc1 : _GEN_12784; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12786 = 8'hf2 == io_state_in_13 ? 8'hdc : _GEN_12785; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12787 = 8'hf3 == io_state_in_13 ? 8'hd7 : _GEN_12786; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12788 = 8'hf4 == io_state_in_13 ? 8'he6 : _GEN_12787; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12789 = 8'hf5 == io_state_in_13 ? 8'hed : _GEN_12788; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12790 = 8'hf6 == io_state_in_13 ? 8'hf0 : _GEN_12789; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12791 = 8'hf7 == io_state_in_13 ? 8'hfb : _GEN_12790; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12792 = 8'hf8 == io_state_in_13 ? 8'h92 : _GEN_12791; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12793 = 8'hf9 == io_state_in_13 ? 8'h99 : _GEN_12792; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12794 = 8'hfa == io_state_in_13 ? 8'h84 : _GEN_12793; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12795 = 8'hfb == io_state_in_13 ? 8'h8f : _GEN_12794; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12796 = 8'hfc == io_state_in_13 ? 8'hbe : _GEN_12795; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12797 = 8'hfd == io_state_in_13 ? 8'hb5 : _GEN_12796; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12798 = 8'hfe == io_state_in_13 ? 8'ha8 : _GEN_12797; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _GEN_12799 = 8'hff == io_state_in_13 ? 8'ha3 : _GEN_12798; // @[InvMixColumns.scala 141:{43,43}]
  wire [7:0] _tmp_state_12_T = _GEN_12543 ^ _GEN_12799; // @[InvMixColumns.scala 141:43]
  wire [7:0] _GEN_12801 = 8'h1 == io_state_in_14 ? 8'hd : 8'h0; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12802 = 8'h2 == io_state_in_14 ? 8'h1a : _GEN_12801; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12803 = 8'h3 == io_state_in_14 ? 8'h17 : _GEN_12802; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12804 = 8'h4 == io_state_in_14 ? 8'h34 : _GEN_12803; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12805 = 8'h5 == io_state_in_14 ? 8'h39 : _GEN_12804; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12806 = 8'h6 == io_state_in_14 ? 8'h2e : _GEN_12805; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12807 = 8'h7 == io_state_in_14 ? 8'h23 : _GEN_12806; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12808 = 8'h8 == io_state_in_14 ? 8'h68 : _GEN_12807; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12809 = 8'h9 == io_state_in_14 ? 8'h65 : _GEN_12808; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12810 = 8'ha == io_state_in_14 ? 8'h72 : _GEN_12809; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12811 = 8'hb == io_state_in_14 ? 8'h7f : _GEN_12810; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12812 = 8'hc == io_state_in_14 ? 8'h5c : _GEN_12811; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12813 = 8'hd == io_state_in_14 ? 8'h51 : _GEN_12812; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12814 = 8'he == io_state_in_14 ? 8'h46 : _GEN_12813; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12815 = 8'hf == io_state_in_14 ? 8'h4b : _GEN_12814; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12816 = 8'h10 == io_state_in_14 ? 8'hd0 : _GEN_12815; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12817 = 8'h11 == io_state_in_14 ? 8'hdd : _GEN_12816; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12818 = 8'h12 == io_state_in_14 ? 8'hca : _GEN_12817; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12819 = 8'h13 == io_state_in_14 ? 8'hc7 : _GEN_12818; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12820 = 8'h14 == io_state_in_14 ? 8'he4 : _GEN_12819; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12821 = 8'h15 == io_state_in_14 ? 8'he9 : _GEN_12820; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12822 = 8'h16 == io_state_in_14 ? 8'hfe : _GEN_12821; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12823 = 8'h17 == io_state_in_14 ? 8'hf3 : _GEN_12822; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12824 = 8'h18 == io_state_in_14 ? 8'hb8 : _GEN_12823; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12825 = 8'h19 == io_state_in_14 ? 8'hb5 : _GEN_12824; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12826 = 8'h1a == io_state_in_14 ? 8'ha2 : _GEN_12825; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12827 = 8'h1b == io_state_in_14 ? 8'haf : _GEN_12826; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12828 = 8'h1c == io_state_in_14 ? 8'h8c : _GEN_12827; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12829 = 8'h1d == io_state_in_14 ? 8'h81 : _GEN_12828; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12830 = 8'h1e == io_state_in_14 ? 8'h96 : _GEN_12829; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12831 = 8'h1f == io_state_in_14 ? 8'h9b : _GEN_12830; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12832 = 8'h20 == io_state_in_14 ? 8'hbb : _GEN_12831; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12833 = 8'h21 == io_state_in_14 ? 8'hb6 : _GEN_12832; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12834 = 8'h22 == io_state_in_14 ? 8'ha1 : _GEN_12833; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12835 = 8'h23 == io_state_in_14 ? 8'hac : _GEN_12834; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12836 = 8'h24 == io_state_in_14 ? 8'h8f : _GEN_12835; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12837 = 8'h25 == io_state_in_14 ? 8'h82 : _GEN_12836; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12838 = 8'h26 == io_state_in_14 ? 8'h95 : _GEN_12837; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12839 = 8'h27 == io_state_in_14 ? 8'h98 : _GEN_12838; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12840 = 8'h28 == io_state_in_14 ? 8'hd3 : _GEN_12839; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12841 = 8'h29 == io_state_in_14 ? 8'hde : _GEN_12840; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12842 = 8'h2a == io_state_in_14 ? 8'hc9 : _GEN_12841; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12843 = 8'h2b == io_state_in_14 ? 8'hc4 : _GEN_12842; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12844 = 8'h2c == io_state_in_14 ? 8'he7 : _GEN_12843; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12845 = 8'h2d == io_state_in_14 ? 8'hea : _GEN_12844; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12846 = 8'h2e == io_state_in_14 ? 8'hfd : _GEN_12845; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12847 = 8'h2f == io_state_in_14 ? 8'hf0 : _GEN_12846; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12848 = 8'h30 == io_state_in_14 ? 8'h6b : _GEN_12847; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12849 = 8'h31 == io_state_in_14 ? 8'h66 : _GEN_12848; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12850 = 8'h32 == io_state_in_14 ? 8'h71 : _GEN_12849; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12851 = 8'h33 == io_state_in_14 ? 8'h7c : _GEN_12850; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12852 = 8'h34 == io_state_in_14 ? 8'h5f : _GEN_12851; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12853 = 8'h35 == io_state_in_14 ? 8'h52 : _GEN_12852; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12854 = 8'h36 == io_state_in_14 ? 8'h45 : _GEN_12853; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12855 = 8'h37 == io_state_in_14 ? 8'h48 : _GEN_12854; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12856 = 8'h38 == io_state_in_14 ? 8'h3 : _GEN_12855; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12857 = 8'h39 == io_state_in_14 ? 8'he : _GEN_12856; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12858 = 8'h3a == io_state_in_14 ? 8'h19 : _GEN_12857; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12859 = 8'h3b == io_state_in_14 ? 8'h14 : _GEN_12858; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12860 = 8'h3c == io_state_in_14 ? 8'h37 : _GEN_12859; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12861 = 8'h3d == io_state_in_14 ? 8'h3a : _GEN_12860; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12862 = 8'h3e == io_state_in_14 ? 8'h2d : _GEN_12861; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12863 = 8'h3f == io_state_in_14 ? 8'h20 : _GEN_12862; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12864 = 8'h40 == io_state_in_14 ? 8'h6d : _GEN_12863; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12865 = 8'h41 == io_state_in_14 ? 8'h60 : _GEN_12864; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12866 = 8'h42 == io_state_in_14 ? 8'h77 : _GEN_12865; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12867 = 8'h43 == io_state_in_14 ? 8'h7a : _GEN_12866; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12868 = 8'h44 == io_state_in_14 ? 8'h59 : _GEN_12867; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12869 = 8'h45 == io_state_in_14 ? 8'h54 : _GEN_12868; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12870 = 8'h46 == io_state_in_14 ? 8'h43 : _GEN_12869; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12871 = 8'h47 == io_state_in_14 ? 8'h4e : _GEN_12870; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12872 = 8'h48 == io_state_in_14 ? 8'h5 : _GEN_12871; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12873 = 8'h49 == io_state_in_14 ? 8'h8 : _GEN_12872; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12874 = 8'h4a == io_state_in_14 ? 8'h1f : _GEN_12873; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12875 = 8'h4b == io_state_in_14 ? 8'h12 : _GEN_12874; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12876 = 8'h4c == io_state_in_14 ? 8'h31 : _GEN_12875; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12877 = 8'h4d == io_state_in_14 ? 8'h3c : _GEN_12876; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12878 = 8'h4e == io_state_in_14 ? 8'h2b : _GEN_12877; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12879 = 8'h4f == io_state_in_14 ? 8'h26 : _GEN_12878; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12880 = 8'h50 == io_state_in_14 ? 8'hbd : _GEN_12879; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12881 = 8'h51 == io_state_in_14 ? 8'hb0 : _GEN_12880; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12882 = 8'h52 == io_state_in_14 ? 8'ha7 : _GEN_12881; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12883 = 8'h53 == io_state_in_14 ? 8'haa : _GEN_12882; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12884 = 8'h54 == io_state_in_14 ? 8'h89 : _GEN_12883; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12885 = 8'h55 == io_state_in_14 ? 8'h84 : _GEN_12884; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12886 = 8'h56 == io_state_in_14 ? 8'h93 : _GEN_12885; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12887 = 8'h57 == io_state_in_14 ? 8'h9e : _GEN_12886; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12888 = 8'h58 == io_state_in_14 ? 8'hd5 : _GEN_12887; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12889 = 8'h59 == io_state_in_14 ? 8'hd8 : _GEN_12888; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12890 = 8'h5a == io_state_in_14 ? 8'hcf : _GEN_12889; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12891 = 8'h5b == io_state_in_14 ? 8'hc2 : _GEN_12890; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12892 = 8'h5c == io_state_in_14 ? 8'he1 : _GEN_12891; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12893 = 8'h5d == io_state_in_14 ? 8'hec : _GEN_12892; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12894 = 8'h5e == io_state_in_14 ? 8'hfb : _GEN_12893; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12895 = 8'h5f == io_state_in_14 ? 8'hf6 : _GEN_12894; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12896 = 8'h60 == io_state_in_14 ? 8'hd6 : _GEN_12895; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12897 = 8'h61 == io_state_in_14 ? 8'hdb : _GEN_12896; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12898 = 8'h62 == io_state_in_14 ? 8'hcc : _GEN_12897; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12899 = 8'h63 == io_state_in_14 ? 8'hc1 : _GEN_12898; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12900 = 8'h64 == io_state_in_14 ? 8'he2 : _GEN_12899; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12901 = 8'h65 == io_state_in_14 ? 8'hef : _GEN_12900; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12902 = 8'h66 == io_state_in_14 ? 8'hf8 : _GEN_12901; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12903 = 8'h67 == io_state_in_14 ? 8'hf5 : _GEN_12902; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12904 = 8'h68 == io_state_in_14 ? 8'hbe : _GEN_12903; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12905 = 8'h69 == io_state_in_14 ? 8'hb3 : _GEN_12904; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12906 = 8'h6a == io_state_in_14 ? 8'ha4 : _GEN_12905; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12907 = 8'h6b == io_state_in_14 ? 8'ha9 : _GEN_12906; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12908 = 8'h6c == io_state_in_14 ? 8'h8a : _GEN_12907; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12909 = 8'h6d == io_state_in_14 ? 8'h87 : _GEN_12908; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12910 = 8'h6e == io_state_in_14 ? 8'h90 : _GEN_12909; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12911 = 8'h6f == io_state_in_14 ? 8'h9d : _GEN_12910; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12912 = 8'h70 == io_state_in_14 ? 8'h6 : _GEN_12911; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12913 = 8'h71 == io_state_in_14 ? 8'hb : _GEN_12912; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12914 = 8'h72 == io_state_in_14 ? 8'h1c : _GEN_12913; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12915 = 8'h73 == io_state_in_14 ? 8'h11 : _GEN_12914; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12916 = 8'h74 == io_state_in_14 ? 8'h32 : _GEN_12915; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12917 = 8'h75 == io_state_in_14 ? 8'h3f : _GEN_12916; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12918 = 8'h76 == io_state_in_14 ? 8'h28 : _GEN_12917; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12919 = 8'h77 == io_state_in_14 ? 8'h25 : _GEN_12918; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12920 = 8'h78 == io_state_in_14 ? 8'h6e : _GEN_12919; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12921 = 8'h79 == io_state_in_14 ? 8'h63 : _GEN_12920; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12922 = 8'h7a == io_state_in_14 ? 8'h74 : _GEN_12921; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12923 = 8'h7b == io_state_in_14 ? 8'h79 : _GEN_12922; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12924 = 8'h7c == io_state_in_14 ? 8'h5a : _GEN_12923; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12925 = 8'h7d == io_state_in_14 ? 8'h57 : _GEN_12924; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12926 = 8'h7e == io_state_in_14 ? 8'h40 : _GEN_12925; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12927 = 8'h7f == io_state_in_14 ? 8'h4d : _GEN_12926; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12928 = 8'h80 == io_state_in_14 ? 8'hda : _GEN_12927; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12929 = 8'h81 == io_state_in_14 ? 8'hd7 : _GEN_12928; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12930 = 8'h82 == io_state_in_14 ? 8'hc0 : _GEN_12929; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12931 = 8'h83 == io_state_in_14 ? 8'hcd : _GEN_12930; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12932 = 8'h84 == io_state_in_14 ? 8'hee : _GEN_12931; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12933 = 8'h85 == io_state_in_14 ? 8'he3 : _GEN_12932; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12934 = 8'h86 == io_state_in_14 ? 8'hf4 : _GEN_12933; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12935 = 8'h87 == io_state_in_14 ? 8'hf9 : _GEN_12934; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12936 = 8'h88 == io_state_in_14 ? 8'hb2 : _GEN_12935; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12937 = 8'h89 == io_state_in_14 ? 8'hbf : _GEN_12936; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12938 = 8'h8a == io_state_in_14 ? 8'ha8 : _GEN_12937; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12939 = 8'h8b == io_state_in_14 ? 8'ha5 : _GEN_12938; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12940 = 8'h8c == io_state_in_14 ? 8'h86 : _GEN_12939; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12941 = 8'h8d == io_state_in_14 ? 8'h8b : _GEN_12940; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12942 = 8'h8e == io_state_in_14 ? 8'h9c : _GEN_12941; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12943 = 8'h8f == io_state_in_14 ? 8'h91 : _GEN_12942; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12944 = 8'h90 == io_state_in_14 ? 8'ha : _GEN_12943; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12945 = 8'h91 == io_state_in_14 ? 8'h7 : _GEN_12944; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12946 = 8'h92 == io_state_in_14 ? 8'h10 : _GEN_12945; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12947 = 8'h93 == io_state_in_14 ? 8'h1d : _GEN_12946; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12948 = 8'h94 == io_state_in_14 ? 8'h3e : _GEN_12947; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12949 = 8'h95 == io_state_in_14 ? 8'h33 : _GEN_12948; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12950 = 8'h96 == io_state_in_14 ? 8'h24 : _GEN_12949; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12951 = 8'h97 == io_state_in_14 ? 8'h29 : _GEN_12950; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12952 = 8'h98 == io_state_in_14 ? 8'h62 : _GEN_12951; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12953 = 8'h99 == io_state_in_14 ? 8'h6f : _GEN_12952; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12954 = 8'h9a == io_state_in_14 ? 8'h78 : _GEN_12953; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12955 = 8'h9b == io_state_in_14 ? 8'h75 : _GEN_12954; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12956 = 8'h9c == io_state_in_14 ? 8'h56 : _GEN_12955; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12957 = 8'h9d == io_state_in_14 ? 8'h5b : _GEN_12956; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12958 = 8'h9e == io_state_in_14 ? 8'h4c : _GEN_12957; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12959 = 8'h9f == io_state_in_14 ? 8'h41 : _GEN_12958; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12960 = 8'ha0 == io_state_in_14 ? 8'h61 : _GEN_12959; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12961 = 8'ha1 == io_state_in_14 ? 8'h6c : _GEN_12960; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12962 = 8'ha2 == io_state_in_14 ? 8'h7b : _GEN_12961; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12963 = 8'ha3 == io_state_in_14 ? 8'h76 : _GEN_12962; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12964 = 8'ha4 == io_state_in_14 ? 8'h55 : _GEN_12963; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12965 = 8'ha5 == io_state_in_14 ? 8'h58 : _GEN_12964; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12966 = 8'ha6 == io_state_in_14 ? 8'h4f : _GEN_12965; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12967 = 8'ha7 == io_state_in_14 ? 8'h42 : _GEN_12966; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12968 = 8'ha8 == io_state_in_14 ? 8'h9 : _GEN_12967; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12969 = 8'ha9 == io_state_in_14 ? 8'h4 : _GEN_12968; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12970 = 8'haa == io_state_in_14 ? 8'h13 : _GEN_12969; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12971 = 8'hab == io_state_in_14 ? 8'h1e : _GEN_12970; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12972 = 8'hac == io_state_in_14 ? 8'h3d : _GEN_12971; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12973 = 8'had == io_state_in_14 ? 8'h30 : _GEN_12972; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12974 = 8'hae == io_state_in_14 ? 8'h27 : _GEN_12973; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12975 = 8'haf == io_state_in_14 ? 8'h2a : _GEN_12974; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12976 = 8'hb0 == io_state_in_14 ? 8'hb1 : _GEN_12975; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12977 = 8'hb1 == io_state_in_14 ? 8'hbc : _GEN_12976; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12978 = 8'hb2 == io_state_in_14 ? 8'hab : _GEN_12977; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12979 = 8'hb3 == io_state_in_14 ? 8'ha6 : _GEN_12978; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12980 = 8'hb4 == io_state_in_14 ? 8'h85 : _GEN_12979; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12981 = 8'hb5 == io_state_in_14 ? 8'h88 : _GEN_12980; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12982 = 8'hb6 == io_state_in_14 ? 8'h9f : _GEN_12981; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12983 = 8'hb7 == io_state_in_14 ? 8'h92 : _GEN_12982; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12984 = 8'hb8 == io_state_in_14 ? 8'hd9 : _GEN_12983; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12985 = 8'hb9 == io_state_in_14 ? 8'hd4 : _GEN_12984; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12986 = 8'hba == io_state_in_14 ? 8'hc3 : _GEN_12985; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12987 = 8'hbb == io_state_in_14 ? 8'hce : _GEN_12986; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12988 = 8'hbc == io_state_in_14 ? 8'hed : _GEN_12987; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12989 = 8'hbd == io_state_in_14 ? 8'he0 : _GEN_12988; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12990 = 8'hbe == io_state_in_14 ? 8'hf7 : _GEN_12989; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12991 = 8'hbf == io_state_in_14 ? 8'hfa : _GEN_12990; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12992 = 8'hc0 == io_state_in_14 ? 8'hb7 : _GEN_12991; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12993 = 8'hc1 == io_state_in_14 ? 8'hba : _GEN_12992; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12994 = 8'hc2 == io_state_in_14 ? 8'had : _GEN_12993; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12995 = 8'hc3 == io_state_in_14 ? 8'ha0 : _GEN_12994; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12996 = 8'hc4 == io_state_in_14 ? 8'h83 : _GEN_12995; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12997 = 8'hc5 == io_state_in_14 ? 8'h8e : _GEN_12996; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12998 = 8'hc6 == io_state_in_14 ? 8'h99 : _GEN_12997; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_12999 = 8'hc7 == io_state_in_14 ? 8'h94 : _GEN_12998; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13000 = 8'hc8 == io_state_in_14 ? 8'hdf : _GEN_12999; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13001 = 8'hc9 == io_state_in_14 ? 8'hd2 : _GEN_13000; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13002 = 8'hca == io_state_in_14 ? 8'hc5 : _GEN_13001; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13003 = 8'hcb == io_state_in_14 ? 8'hc8 : _GEN_13002; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13004 = 8'hcc == io_state_in_14 ? 8'heb : _GEN_13003; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13005 = 8'hcd == io_state_in_14 ? 8'he6 : _GEN_13004; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13006 = 8'hce == io_state_in_14 ? 8'hf1 : _GEN_13005; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13007 = 8'hcf == io_state_in_14 ? 8'hfc : _GEN_13006; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13008 = 8'hd0 == io_state_in_14 ? 8'h67 : _GEN_13007; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13009 = 8'hd1 == io_state_in_14 ? 8'h6a : _GEN_13008; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13010 = 8'hd2 == io_state_in_14 ? 8'h7d : _GEN_13009; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13011 = 8'hd3 == io_state_in_14 ? 8'h70 : _GEN_13010; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13012 = 8'hd4 == io_state_in_14 ? 8'h53 : _GEN_13011; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13013 = 8'hd5 == io_state_in_14 ? 8'h5e : _GEN_13012; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13014 = 8'hd6 == io_state_in_14 ? 8'h49 : _GEN_13013; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13015 = 8'hd7 == io_state_in_14 ? 8'h44 : _GEN_13014; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13016 = 8'hd8 == io_state_in_14 ? 8'hf : _GEN_13015; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13017 = 8'hd9 == io_state_in_14 ? 8'h2 : _GEN_13016; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13018 = 8'hda == io_state_in_14 ? 8'h15 : _GEN_13017; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13019 = 8'hdb == io_state_in_14 ? 8'h18 : _GEN_13018; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13020 = 8'hdc == io_state_in_14 ? 8'h3b : _GEN_13019; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13021 = 8'hdd == io_state_in_14 ? 8'h36 : _GEN_13020; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13022 = 8'hde == io_state_in_14 ? 8'h21 : _GEN_13021; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13023 = 8'hdf == io_state_in_14 ? 8'h2c : _GEN_13022; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13024 = 8'he0 == io_state_in_14 ? 8'hc : _GEN_13023; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13025 = 8'he1 == io_state_in_14 ? 8'h1 : _GEN_13024; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13026 = 8'he2 == io_state_in_14 ? 8'h16 : _GEN_13025; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13027 = 8'he3 == io_state_in_14 ? 8'h1b : _GEN_13026; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13028 = 8'he4 == io_state_in_14 ? 8'h38 : _GEN_13027; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13029 = 8'he5 == io_state_in_14 ? 8'h35 : _GEN_13028; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13030 = 8'he6 == io_state_in_14 ? 8'h22 : _GEN_13029; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13031 = 8'he7 == io_state_in_14 ? 8'h2f : _GEN_13030; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13032 = 8'he8 == io_state_in_14 ? 8'h64 : _GEN_13031; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13033 = 8'he9 == io_state_in_14 ? 8'h69 : _GEN_13032; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13034 = 8'hea == io_state_in_14 ? 8'h7e : _GEN_13033; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13035 = 8'heb == io_state_in_14 ? 8'h73 : _GEN_13034; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13036 = 8'hec == io_state_in_14 ? 8'h50 : _GEN_13035; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13037 = 8'hed == io_state_in_14 ? 8'h5d : _GEN_13036; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13038 = 8'hee == io_state_in_14 ? 8'h4a : _GEN_13037; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13039 = 8'hef == io_state_in_14 ? 8'h47 : _GEN_13038; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13040 = 8'hf0 == io_state_in_14 ? 8'hdc : _GEN_13039; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13041 = 8'hf1 == io_state_in_14 ? 8'hd1 : _GEN_13040; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13042 = 8'hf2 == io_state_in_14 ? 8'hc6 : _GEN_13041; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13043 = 8'hf3 == io_state_in_14 ? 8'hcb : _GEN_13042; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13044 = 8'hf4 == io_state_in_14 ? 8'he8 : _GEN_13043; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13045 = 8'hf5 == io_state_in_14 ? 8'he5 : _GEN_13044; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13046 = 8'hf6 == io_state_in_14 ? 8'hf2 : _GEN_13045; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13047 = 8'hf7 == io_state_in_14 ? 8'hff : _GEN_13046; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13048 = 8'hf8 == io_state_in_14 ? 8'hb4 : _GEN_13047; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13049 = 8'hf9 == io_state_in_14 ? 8'hb9 : _GEN_13048; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13050 = 8'hfa == io_state_in_14 ? 8'hae : _GEN_13049; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13051 = 8'hfb == io_state_in_14 ? 8'ha3 : _GEN_13050; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13052 = 8'hfc == io_state_in_14 ? 8'h80 : _GEN_13051; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13053 = 8'hfd == io_state_in_14 ? 8'h8d : _GEN_13052; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13054 = 8'hfe == io_state_in_14 ? 8'h9a : _GEN_13053; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _GEN_13055 = 8'hff == io_state_in_14 ? 8'h97 : _GEN_13054; // @[InvMixColumns.scala 141:{68,68}]
  wire [7:0] _tmp_state_12_T_1 = _tmp_state_12_T ^ _GEN_13055; // @[InvMixColumns.scala 141:68]
  wire [7:0] _GEN_13057 = 8'h1 == io_state_in_15 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13058 = 8'h2 == io_state_in_15 ? 8'h12 : _GEN_13057; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13059 = 8'h3 == io_state_in_15 ? 8'h1b : _GEN_13058; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13060 = 8'h4 == io_state_in_15 ? 8'h24 : _GEN_13059; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13061 = 8'h5 == io_state_in_15 ? 8'h2d : _GEN_13060; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13062 = 8'h6 == io_state_in_15 ? 8'h36 : _GEN_13061; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13063 = 8'h7 == io_state_in_15 ? 8'h3f : _GEN_13062; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13064 = 8'h8 == io_state_in_15 ? 8'h48 : _GEN_13063; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13065 = 8'h9 == io_state_in_15 ? 8'h41 : _GEN_13064; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13066 = 8'ha == io_state_in_15 ? 8'h5a : _GEN_13065; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13067 = 8'hb == io_state_in_15 ? 8'h53 : _GEN_13066; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13068 = 8'hc == io_state_in_15 ? 8'h6c : _GEN_13067; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13069 = 8'hd == io_state_in_15 ? 8'h65 : _GEN_13068; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13070 = 8'he == io_state_in_15 ? 8'h7e : _GEN_13069; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13071 = 8'hf == io_state_in_15 ? 8'h77 : _GEN_13070; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13072 = 8'h10 == io_state_in_15 ? 8'h90 : _GEN_13071; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13073 = 8'h11 == io_state_in_15 ? 8'h99 : _GEN_13072; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13074 = 8'h12 == io_state_in_15 ? 8'h82 : _GEN_13073; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13075 = 8'h13 == io_state_in_15 ? 8'h8b : _GEN_13074; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13076 = 8'h14 == io_state_in_15 ? 8'hb4 : _GEN_13075; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13077 = 8'h15 == io_state_in_15 ? 8'hbd : _GEN_13076; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13078 = 8'h16 == io_state_in_15 ? 8'ha6 : _GEN_13077; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13079 = 8'h17 == io_state_in_15 ? 8'haf : _GEN_13078; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13080 = 8'h18 == io_state_in_15 ? 8'hd8 : _GEN_13079; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13081 = 8'h19 == io_state_in_15 ? 8'hd1 : _GEN_13080; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13082 = 8'h1a == io_state_in_15 ? 8'hca : _GEN_13081; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13083 = 8'h1b == io_state_in_15 ? 8'hc3 : _GEN_13082; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13084 = 8'h1c == io_state_in_15 ? 8'hfc : _GEN_13083; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13085 = 8'h1d == io_state_in_15 ? 8'hf5 : _GEN_13084; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13086 = 8'h1e == io_state_in_15 ? 8'hee : _GEN_13085; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13087 = 8'h1f == io_state_in_15 ? 8'he7 : _GEN_13086; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13088 = 8'h20 == io_state_in_15 ? 8'h3b : _GEN_13087; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13089 = 8'h21 == io_state_in_15 ? 8'h32 : _GEN_13088; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13090 = 8'h22 == io_state_in_15 ? 8'h29 : _GEN_13089; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13091 = 8'h23 == io_state_in_15 ? 8'h20 : _GEN_13090; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13092 = 8'h24 == io_state_in_15 ? 8'h1f : _GEN_13091; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13093 = 8'h25 == io_state_in_15 ? 8'h16 : _GEN_13092; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13094 = 8'h26 == io_state_in_15 ? 8'hd : _GEN_13093; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13095 = 8'h27 == io_state_in_15 ? 8'h4 : _GEN_13094; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13096 = 8'h28 == io_state_in_15 ? 8'h73 : _GEN_13095; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13097 = 8'h29 == io_state_in_15 ? 8'h7a : _GEN_13096; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13098 = 8'h2a == io_state_in_15 ? 8'h61 : _GEN_13097; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13099 = 8'h2b == io_state_in_15 ? 8'h68 : _GEN_13098; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13100 = 8'h2c == io_state_in_15 ? 8'h57 : _GEN_13099; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13101 = 8'h2d == io_state_in_15 ? 8'h5e : _GEN_13100; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13102 = 8'h2e == io_state_in_15 ? 8'h45 : _GEN_13101; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13103 = 8'h2f == io_state_in_15 ? 8'h4c : _GEN_13102; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13104 = 8'h30 == io_state_in_15 ? 8'hab : _GEN_13103; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13105 = 8'h31 == io_state_in_15 ? 8'ha2 : _GEN_13104; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13106 = 8'h32 == io_state_in_15 ? 8'hb9 : _GEN_13105; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13107 = 8'h33 == io_state_in_15 ? 8'hb0 : _GEN_13106; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13108 = 8'h34 == io_state_in_15 ? 8'h8f : _GEN_13107; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13109 = 8'h35 == io_state_in_15 ? 8'h86 : _GEN_13108; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13110 = 8'h36 == io_state_in_15 ? 8'h9d : _GEN_13109; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13111 = 8'h37 == io_state_in_15 ? 8'h94 : _GEN_13110; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13112 = 8'h38 == io_state_in_15 ? 8'he3 : _GEN_13111; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13113 = 8'h39 == io_state_in_15 ? 8'hea : _GEN_13112; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13114 = 8'h3a == io_state_in_15 ? 8'hf1 : _GEN_13113; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13115 = 8'h3b == io_state_in_15 ? 8'hf8 : _GEN_13114; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13116 = 8'h3c == io_state_in_15 ? 8'hc7 : _GEN_13115; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13117 = 8'h3d == io_state_in_15 ? 8'hce : _GEN_13116; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13118 = 8'h3e == io_state_in_15 ? 8'hd5 : _GEN_13117; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13119 = 8'h3f == io_state_in_15 ? 8'hdc : _GEN_13118; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13120 = 8'h40 == io_state_in_15 ? 8'h76 : _GEN_13119; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13121 = 8'h41 == io_state_in_15 ? 8'h7f : _GEN_13120; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13122 = 8'h42 == io_state_in_15 ? 8'h64 : _GEN_13121; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13123 = 8'h43 == io_state_in_15 ? 8'h6d : _GEN_13122; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13124 = 8'h44 == io_state_in_15 ? 8'h52 : _GEN_13123; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13125 = 8'h45 == io_state_in_15 ? 8'h5b : _GEN_13124; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13126 = 8'h46 == io_state_in_15 ? 8'h40 : _GEN_13125; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13127 = 8'h47 == io_state_in_15 ? 8'h49 : _GEN_13126; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13128 = 8'h48 == io_state_in_15 ? 8'h3e : _GEN_13127; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13129 = 8'h49 == io_state_in_15 ? 8'h37 : _GEN_13128; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13130 = 8'h4a == io_state_in_15 ? 8'h2c : _GEN_13129; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13131 = 8'h4b == io_state_in_15 ? 8'h25 : _GEN_13130; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13132 = 8'h4c == io_state_in_15 ? 8'h1a : _GEN_13131; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13133 = 8'h4d == io_state_in_15 ? 8'h13 : _GEN_13132; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13134 = 8'h4e == io_state_in_15 ? 8'h8 : _GEN_13133; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13135 = 8'h4f == io_state_in_15 ? 8'h1 : _GEN_13134; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13136 = 8'h50 == io_state_in_15 ? 8'he6 : _GEN_13135; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13137 = 8'h51 == io_state_in_15 ? 8'hef : _GEN_13136; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13138 = 8'h52 == io_state_in_15 ? 8'hf4 : _GEN_13137; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13139 = 8'h53 == io_state_in_15 ? 8'hfd : _GEN_13138; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13140 = 8'h54 == io_state_in_15 ? 8'hc2 : _GEN_13139; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13141 = 8'h55 == io_state_in_15 ? 8'hcb : _GEN_13140; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13142 = 8'h56 == io_state_in_15 ? 8'hd0 : _GEN_13141; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13143 = 8'h57 == io_state_in_15 ? 8'hd9 : _GEN_13142; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13144 = 8'h58 == io_state_in_15 ? 8'hae : _GEN_13143; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13145 = 8'h59 == io_state_in_15 ? 8'ha7 : _GEN_13144; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13146 = 8'h5a == io_state_in_15 ? 8'hbc : _GEN_13145; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13147 = 8'h5b == io_state_in_15 ? 8'hb5 : _GEN_13146; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13148 = 8'h5c == io_state_in_15 ? 8'h8a : _GEN_13147; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13149 = 8'h5d == io_state_in_15 ? 8'h83 : _GEN_13148; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13150 = 8'h5e == io_state_in_15 ? 8'h98 : _GEN_13149; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13151 = 8'h5f == io_state_in_15 ? 8'h91 : _GEN_13150; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13152 = 8'h60 == io_state_in_15 ? 8'h4d : _GEN_13151; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13153 = 8'h61 == io_state_in_15 ? 8'h44 : _GEN_13152; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13154 = 8'h62 == io_state_in_15 ? 8'h5f : _GEN_13153; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13155 = 8'h63 == io_state_in_15 ? 8'h56 : _GEN_13154; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13156 = 8'h64 == io_state_in_15 ? 8'h69 : _GEN_13155; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13157 = 8'h65 == io_state_in_15 ? 8'h60 : _GEN_13156; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13158 = 8'h66 == io_state_in_15 ? 8'h7b : _GEN_13157; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13159 = 8'h67 == io_state_in_15 ? 8'h72 : _GEN_13158; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13160 = 8'h68 == io_state_in_15 ? 8'h5 : _GEN_13159; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13161 = 8'h69 == io_state_in_15 ? 8'hc : _GEN_13160; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13162 = 8'h6a == io_state_in_15 ? 8'h17 : _GEN_13161; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13163 = 8'h6b == io_state_in_15 ? 8'h1e : _GEN_13162; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13164 = 8'h6c == io_state_in_15 ? 8'h21 : _GEN_13163; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13165 = 8'h6d == io_state_in_15 ? 8'h28 : _GEN_13164; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13166 = 8'h6e == io_state_in_15 ? 8'h33 : _GEN_13165; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13167 = 8'h6f == io_state_in_15 ? 8'h3a : _GEN_13166; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13168 = 8'h70 == io_state_in_15 ? 8'hdd : _GEN_13167; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13169 = 8'h71 == io_state_in_15 ? 8'hd4 : _GEN_13168; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13170 = 8'h72 == io_state_in_15 ? 8'hcf : _GEN_13169; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13171 = 8'h73 == io_state_in_15 ? 8'hc6 : _GEN_13170; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13172 = 8'h74 == io_state_in_15 ? 8'hf9 : _GEN_13171; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13173 = 8'h75 == io_state_in_15 ? 8'hf0 : _GEN_13172; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13174 = 8'h76 == io_state_in_15 ? 8'heb : _GEN_13173; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13175 = 8'h77 == io_state_in_15 ? 8'he2 : _GEN_13174; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13176 = 8'h78 == io_state_in_15 ? 8'h95 : _GEN_13175; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13177 = 8'h79 == io_state_in_15 ? 8'h9c : _GEN_13176; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13178 = 8'h7a == io_state_in_15 ? 8'h87 : _GEN_13177; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13179 = 8'h7b == io_state_in_15 ? 8'h8e : _GEN_13178; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13180 = 8'h7c == io_state_in_15 ? 8'hb1 : _GEN_13179; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13181 = 8'h7d == io_state_in_15 ? 8'hb8 : _GEN_13180; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13182 = 8'h7e == io_state_in_15 ? 8'ha3 : _GEN_13181; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13183 = 8'h7f == io_state_in_15 ? 8'haa : _GEN_13182; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13184 = 8'h80 == io_state_in_15 ? 8'hec : _GEN_13183; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13185 = 8'h81 == io_state_in_15 ? 8'he5 : _GEN_13184; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13186 = 8'h82 == io_state_in_15 ? 8'hfe : _GEN_13185; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13187 = 8'h83 == io_state_in_15 ? 8'hf7 : _GEN_13186; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13188 = 8'h84 == io_state_in_15 ? 8'hc8 : _GEN_13187; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13189 = 8'h85 == io_state_in_15 ? 8'hc1 : _GEN_13188; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13190 = 8'h86 == io_state_in_15 ? 8'hda : _GEN_13189; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13191 = 8'h87 == io_state_in_15 ? 8'hd3 : _GEN_13190; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13192 = 8'h88 == io_state_in_15 ? 8'ha4 : _GEN_13191; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13193 = 8'h89 == io_state_in_15 ? 8'had : _GEN_13192; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13194 = 8'h8a == io_state_in_15 ? 8'hb6 : _GEN_13193; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13195 = 8'h8b == io_state_in_15 ? 8'hbf : _GEN_13194; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13196 = 8'h8c == io_state_in_15 ? 8'h80 : _GEN_13195; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13197 = 8'h8d == io_state_in_15 ? 8'h89 : _GEN_13196; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13198 = 8'h8e == io_state_in_15 ? 8'h92 : _GEN_13197; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13199 = 8'h8f == io_state_in_15 ? 8'h9b : _GEN_13198; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13200 = 8'h90 == io_state_in_15 ? 8'h7c : _GEN_13199; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13201 = 8'h91 == io_state_in_15 ? 8'h75 : _GEN_13200; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13202 = 8'h92 == io_state_in_15 ? 8'h6e : _GEN_13201; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13203 = 8'h93 == io_state_in_15 ? 8'h67 : _GEN_13202; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13204 = 8'h94 == io_state_in_15 ? 8'h58 : _GEN_13203; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13205 = 8'h95 == io_state_in_15 ? 8'h51 : _GEN_13204; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13206 = 8'h96 == io_state_in_15 ? 8'h4a : _GEN_13205; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13207 = 8'h97 == io_state_in_15 ? 8'h43 : _GEN_13206; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13208 = 8'h98 == io_state_in_15 ? 8'h34 : _GEN_13207; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13209 = 8'h99 == io_state_in_15 ? 8'h3d : _GEN_13208; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13210 = 8'h9a == io_state_in_15 ? 8'h26 : _GEN_13209; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13211 = 8'h9b == io_state_in_15 ? 8'h2f : _GEN_13210; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13212 = 8'h9c == io_state_in_15 ? 8'h10 : _GEN_13211; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13213 = 8'h9d == io_state_in_15 ? 8'h19 : _GEN_13212; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13214 = 8'h9e == io_state_in_15 ? 8'h2 : _GEN_13213; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13215 = 8'h9f == io_state_in_15 ? 8'hb : _GEN_13214; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13216 = 8'ha0 == io_state_in_15 ? 8'hd7 : _GEN_13215; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13217 = 8'ha1 == io_state_in_15 ? 8'hde : _GEN_13216; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13218 = 8'ha2 == io_state_in_15 ? 8'hc5 : _GEN_13217; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13219 = 8'ha3 == io_state_in_15 ? 8'hcc : _GEN_13218; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13220 = 8'ha4 == io_state_in_15 ? 8'hf3 : _GEN_13219; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13221 = 8'ha5 == io_state_in_15 ? 8'hfa : _GEN_13220; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13222 = 8'ha6 == io_state_in_15 ? 8'he1 : _GEN_13221; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13223 = 8'ha7 == io_state_in_15 ? 8'he8 : _GEN_13222; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13224 = 8'ha8 == io_state_in_15 ? 8'h9f : _GEN_13223; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13225 = 8'ha9 == io_state_in_15 ? 8'h96 : _GEN_13224; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13226 = 8'haa == io_state_in_15 ? 8'h8d : _GEN_13225; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13227 = 8'hab == io_state_in_15 ? 8'h84 : _GEN_13226; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13228 = 8'hac == io_state_in_15 ? 8'hbb : _GEN_13227; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13229 = 8'had == io_state_in_15 ? 8'hb2 : _GEN_13228; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13230 = 8'hae == io_state_in_15 ? 8'ha9 : _GEN_13229; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13231 = 8'haf == io_state_in_15 ? 8'ha0 : _GEN_13230; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13232 = 8'hb0 == io_state_in_15 ? 8'h47 : _GEN_13231; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13233 = 8'hb1 == io_state_in_15 ? 8'h4e : _GEN_13232; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13234 = 8'hb2 == io_state_in_15 ? 8'h55 : _GEN_13233; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13235 = 8'hb3 == io_state_in_15 ? 8'h5c : _GEN_13234; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13236 = 8'hb4 == io_state_in_15 ? 8'h63 : _GEN_13235; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13237 = 8'hb5 == io_state_in_15 ? 8'h6a : _GEN_13236; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13238 = 8'hb6 == io_state_in_15 ? 8'h71 : _GEN_13237; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13239 = 8'hb7 == io_state_in_15 ? 8'h78 : _GEN_13238; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13240 = 8'hb8 == io_state_in_15 ? 8'hf : _GEN_13239; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13241 = 8'hb9 == io_state_in_15 ? 8'h6 : _GEN_13240; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13242 = 8'hba == io_state_in_15 ? 8'h1d : _GEN_13241; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13243 = 8'hbb == io_state_in_15 ? 8'h14 : _GEN_13242; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13244 = 8'hbc == io_state_in_15 ? 8'h2b : _GEN_13243; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13245 = 8'hbd == io_state_in_15 ? 8'h22 : _GEN_13244; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13246 = 8'hbe == io_state_in_15 ? 8'h39 : _GEN_13245; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13247 = 8'hbf == io_state_in_15 ? 8'h30 : _GEN_13246; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13248 = 8'hc0 == io_state_in_15 ? 8'h9a : _GEN_13247; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13249 = 8'hc1 == io_state_in_15 ? 8'h93 : _GEN_13248; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13250 = 8'hc2 == io_state_in_15 ? 8'h88 : _GEN_13249; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13251 = 8'hc3 == io_state_in_15 ? 8'h81 : _GEN_13250; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13252 = 8'hc4 == io_state_in_15 ? 8'hbe : _GEN_13251; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13253 = 8'hc5 == io_state_in_15 ? 8'hb7 : _GEN_13252; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13254 = 8'hc6 == io_state_in_15 ? 8'hac : _GEN_13253; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13255 = 8'hc7 == io_state_in_15 ? 8'ha5 : _GEN_13254; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13256 = 8'hc8 == io_state_in_15 ? 8'hd2 : _GEN_13255; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13257 = 8'hc9 == io_state_in_15 ? 8'hdb : _GEN_13256; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13258 = 8'hca == io_state_in_15 ? 8'hc0 : _GEN_13257; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13259 = 8'hcb == io_state_in_15 ? 8'hc9 : _GEN_13258; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13260 = 8'hcc == io_state_in_15 ? 8'hf6 : _GEN_13259; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13261 = 8'hcd == io_state_in_15 ? 8'hff : _GEN_13260; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13262 = 8'hce == io_state_in_15 ? 8'he4 : _GEN_13261; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13263 = 8'hcf == io_state_in_15 ? 8'hed : _GEN_13262; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13264 = 8'hd0 == io_state_in_15 ? 8'ha : _GEN_13263; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13265 = 8'hd1 == io_state_in_15 ? 8'h3 : _GEN_13264; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13266 = 8'hd2 == io_state_in_15 ? 8'h18 : _GEN_13265; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13267 = 8'hd3 == io_state_in_15 ? 8'h11 : _GEN_13266; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13268 = 8'hd4 == io_state_in_15 ? 8'h2e : _GEN_13267; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13269 = 8'hd5 == io_state_in_15 ? 8'h27 : _GEN_13268; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13270 = 8'hd6 == io_state_in_15 ? 8'h3c : _GEN_13269; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13271 = 8'hd7 == io_state_in_15 ? 8'h35 : _GEN_13270; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13272 = 8'hd8 == io_state_in_15 ? 8'h42 : _GEN_13271; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13273 = 8'hd9 == io_state_in_15 ? 8'h4b : _GEN_13272; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13274 = 8'hda == io_state_in_15 ? 8'h50 : _GEN_13273; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13275 = 8'hdb == io_state_in_15 ? 8'h59 : _GEN_13274; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13276 = 8'hdc == io_state_in_15 ? 8'h66 : _GEN_13275; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13277 = 8'hdd == io_state_in_15 ? 8'h6f : _GEN_13276; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13278 = 8'hde == io_state_in_15 ? 8'h74 : _GEN_13277; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13279 = 8'hdf == io_state_in_15 ? 8'h7d : _GEN_13278; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13280 = 8'he0 == io_state_in_15 ? 8'ha1 : _GEN_13279; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13281 = 8'he1 == io_state_in_15 ? 8'ha8 : _GEN_13280; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13282 = 8'he2 == io_state_in_15 ? 8'hb3 : _GEN_13281; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13283 = 8'he3 == io_state_in_15 ? 8'hba : _GEN_13282; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13284 = 8'he4 == io_state_in_15 ? 8'h85 : _GEN_13283; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13285 = 8'he5 == io_state_in_15 ? 8'h8c : _GEN_13284; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13286 = 8'he6 == io_state_in_15 ? 8'h97 : _GEN_13285; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13287 = 8'he7 == io_state_in_15 ? 8'h9e : _GEN_13286; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13288 = 8'he8 == io_state_in_15 ? 8'he9 : _GEN_13287; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13289 = 8'he9 == io_state_in_15 ? 8'he0 : _GEN_13288; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13290 = 8'hea == io_state_in_15 ? 8'hfb : _GEN_13289; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13291 = 8'heb == io_state_in_15 ? 8'hf2 : _GEN_13290; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13292 = 8'hec == io_state_in_15 ? 8'hcd : _GEN_13291; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13293 = 8'hed == io_state_in_15 ? 8'hc4 : _GEN_13292; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13294 = 8'hee == io_state_in_15 ? 8'hdf : _GEN_13293; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13295 = 8'hef == io_state_in_15 ? 8'hd6 : _GEN_13294; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13296 = 8'hf0 == io_state_in_15 ? 8'h31 : _GEN_13295; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13297 = 8'hf1 == io_state_in_15 ? 8'h38 : _GEN_13296; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13298 = 8'hf2 == io_state_in_15 ? 8'h23 : _GEN_13297; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13299 = 8'hf3 == io_state_in_15 ? 8'h2a : _GEN_13298; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13300 = 8'hf4 == io_state_in_15 ? 8'h15 : _GEN_13299; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13301 = 8'hf5 == io_state_in_15 ? 8'h1c : _GEN_13300; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13302 = 8'hf6 == io_state_in_15 ? 8'h7 : _GEN_13301; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13303 = 8'hf7 == io_state_in_15 ? 8'he : _GEN_13302; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13304 = 8'hf8 == io_state_in_15 ? 8'h79 : _GEN_13303; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13305 = 8'hf9 == io_state_in_15 ? 8'h70 : _GEN_13304; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13306 = 8'hfa == io_state_in_15 ? 8'h6b : _GEN_13305; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13307 = 8'hfb == io_state_in_15 ? 8'h62 : _GEN_13306; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13308 = 8'hfc == io_state_in_15 ? 8'h5d : _GEN_13307; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13309 = 8'hfd == io_state_in_15 ? 8'h54 : _GEN_13308; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13310 = 8'hfe == io_state_in_15 ? 8'h4f : _GEN_13309; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13311 = 8'hff == io_state_in_15 ? 8'h46 : _GEN_13310; // @[InvMixColumns.scala 141:{93,93}]
  wire [7:0] _GEN_13313 = 8'h1 == io_state_in_12 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13314 = 8'h2 == io_state_in_12 ? 8'h12 : _GEN_13313; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13315 = 8'h3 == io_state_in_12 ? 8'h1b : _GEN_13314; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13316 = 8'h4 == io_state_in_12 ? 8'h24 : _GEN_13315; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13317 = 8'h5 == io_state_in_12 ? 8'h2d : _GEN_13316; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13318 = 8'h6 == io_state_in_12 ? 8'h36 : _GEN_13317; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13319 = 8'h7 == io_state_in_12 ? 8'h3f : _GEN_13318; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13320 = 8'h8 == io_state_in_12 ? 8'h48 : _GEN_13319; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13321 = 8'h9 == io_state_in_12 ? 8'h41 : _GEN_13320; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13322 = 8'ha == io_state_in_12 ? 8'h5a : _GEN_13321; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13323 = 8'hb == io_state_in_12 ? 8'h53 : _GEN_13322; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13324 = 8'hc == io_state_in_12 ? 8'h6c : _GEN_13323; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13325 = 8'hd == io_state_in_12 ? 8'h65 : _GEN_13324; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13326 = 8'he == io_state_in_12 ? 8'h7e : _GEN_13325; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13327 = 8'hf == io_state_in_12 ? 8'h77 : _GEN_13326; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13328 = 8'h10 == io_state_in_12 ? 8'h90 : _GEN_13327; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13329 = 8'h11 == io_state_in_12 ? 8'h99 : _GEN_13328; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13330 = 8'h12 == io_state_in_12 ? 8'h82 : _GEN_13329; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13331 = 8'h13 == io_state_in_12 ? 8'h8b : _GEN_13330; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13332 = 8'h14 == io_state_in_12 ? 8'hb4 : _GEN_13331; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13333 = 8'h15 == io_state_in_12 ? 8'hbd : _GEN_13332; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13334 = 8'h16 == io_state_in_12 ? 8'ha6 : _GEN_13333; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13335 = 8'h17 == io_state_in_12 ? 8'haf : _GEN_13334; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13336 = 8'h18 == io_state_in_12 ? 8'hd8 : _GEN_13335; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13337 = 8'h19 == io_state_in_12 ? 8'hd1 : _GEN_13336; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13338 = 8'h1a == io_state_in_12 ? 8'hca : _GEN_13337; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13339 = 8'h1b == io_state_in_12 ? 8'hc3 : _GEN_13338; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13340 = 8'h1c == io_state_in_12 ? 8'hfc : _GEN_13339; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13341 = 8'h1d == io_state_in_12 ? 8'hf5 : _GEN_13340; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13342 = 8'h1e == io_state_in_12 ? 8'hee : _GEN_13341; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13343 = 8'h1f == io_state_in_12 ? 8'he7 : _GEN_13342; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13344 = 8'h20 == io_state_in_12 ? 8'h3b : _GEN_13343; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13345 = 8'h21 == io_state_in_12 ? 8'h32 : _GEN_13344; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13346 = 8'h22 == io_state_in_12 ? 8'h29 : _GEN_13345; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13347 = 8'h23 == io_state_in_12 ? 8'h20 : _GEN_13346; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13348 = 8'h24 == io_state_in_12 ? 8'h1f : _GEN_13347; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13349 = 8'h25 == io_state_in_12 ? 8'h16 : _GEN_13348; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13350 = 8'h26 == io_state_in_12 ? 8'hd : _GEN_13349; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13351 = 8'h27 == io_state_in_12 ? 8'h4 : _GEN_13350; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13352 = 8'h28 == io_state_in_12 ? 8'h73 : _GEN_13351; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13353 = 8'h29 == io_state_in_12 ? 8'h7a : _GEN_13352; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13354 = 8'h2a == io_state_in_12 ? 8'h61 : _GEN_13353; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13355 = 8'h2b == io_state_in_12 ? 8'h68 : _GEN_13354; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13356 = 8'h2c == io_state_in_12 ? 8'h57 : _GEN_13355; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13357 = 8'h2d == io_state_in_12 ? 8'h5e : _GEN_13356; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13358 = 8'h2e == io_state_in_12 ? 8'h45 : _GEN_13357; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13359 = 8'h2f == io_state_in_12 ? 8'h4c : _GEN_13358; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13360 = 8'h30 == io_state_in_12 ? 8'hab : _GEN_13359; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13361 = 8'h31 == io_state_in_12 ? 8'ha2 : _GEN_13360; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13362 = 8'h32 == io_state_in_12 ? 8'hb9 : _GEN_13361; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13363 = 8'h33 == io_state_in_12 ? 8'hb0 : _GEN_13362; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13364 = 8'h34 == io_state_in_12 ? 8'h8f : _GEN_13363; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13365 = 8'h35 == io_state_in_12 ? 8'h86 : _GEN_13364; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13366 = 8'h36 == io_state_in_12 ? 8'h9d : _GEN_13365; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13367 = 8'h37 == io_state_in_12 ? 8'h94 : _GEN_13366; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13368 = 8'h38 == io_state_in_12 ? 8'he3 : _GEN_13367; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13369 = 8'h39 == io_state_in_12 ? 8'hea : _GEN_13368; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13370 = 8'h3a == io_state_in_12 ? 8'hf1 : _GEN_13369; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13371 = 8'h3b == io_state_in_12 ? 8'hf8 : _GEN_13370; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13372 = 8'h3c == io_state_in_12 ? 8'hc7 : _GEN_13371; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13373 = 8'h3d == io_state_in_12 ? 8'hce : _GEN_13372; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13374 = 8'h3e == io_state_in_12 ? 8'hd5 : _GEN_13373; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13375 = 8'h3f == io_state_in_12 ? 8'hdc : _GEN_13374; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13376 = 8'h40 == io_state_in_12 ? 8'h76 : _GEN_13375; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13377 = 8'h41 == io_state_in_12 ? 8'h7f : _GEN_13376; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13378 = 8'h42 == io_state_in_12 ? 8'h64 : _GEN_13377; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13379 = 8'h43 == io_state_in_12 ? 8'h6d : _GEN_13378; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13380 = 8'h44 == io_state_in_12 ? 8'h52 : _GEN_13379; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13381 = 8'h45 == io_state_in_12 ? 8'h5b : _GEN_13380; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13382 = 8'h46 == io_state_in_12 ? 8'h40 : _GEN_13381; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13383 = 8'h47 == io_state_in_12 ? 8'h49 : _GEN_13382; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13384 = 8'h48 == io_state_in_12 ? 8'h3e : _GEN_13383; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13385 = 8'h49 == io_state_in_12 ? 8'h37 : _GEN_13384; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13386 = 8'h4a == io_state_in_12 ? 8'h2c : _GEN_13385; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13387 = 8'h4b == io_state_in_12 ? 8'h25 : _GEN_13386; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13388 = 8'h4c == io_state_in_12 ? 8'h1a : _GEN_13387; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13389 = 8'h4d == io_state_in_12 ? 8'h13 : _GEN_13388; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13390 = 8'h4e == io_state_in_12 ? 8'h8 : _GEN_13389; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13391 = 8'h4f == io_state_in_12 ? 8'h1 : _GEN_13390; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13392 = 8'h50 == io_state_in_12 ? 8'he6 : _GEN_13391; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13393 = 8'h51 == io_state_in_12 ? 8'hef : _GEN_13392; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13394 = 8'h52 == io_state_in_12 ? 8'hf4 : _GEN_13393; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13395 = 8'h53 == io_state_in_12 ? 8'hfd : _GEN_13394; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13396 = 8'h54 == io_state_in_12 ? 8'hc2 : _GEN_13395; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13397 = 8'h55 == io_state_in_12 ? 8'hcb : _GEN_13396; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13398 = 8'h56 == io_state_in_12 ? 8'hd0 : _GEN_13397; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13399 = 8'h57 == io_state_in_12 ? 8'hd9 : _GEN_13398; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13400 = 8'h58 == io_state_in_12 ? 8'hae : _GEN_13399; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13401 = 8'h59 == io_state_in_12 ? 8'ha7 : _GEN_13400; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13402 = 8'h5a == io_state_in_12 ? 8'hbc : _GEN_13401; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13403 = 8'h5b == io_state_in_12 ? 8'hb5 : _GEN_13402; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13404 = 8'h5c == io_state_in_12 ? 8'h8a : _GEN_13403; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13405 = 8'h5d == io_state_in_12 ? 8'h83 : _GEN_13404; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13406 = 8'h5e == io_state_in_12 ? 8'h98 : _GEN_13405; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13407 = 8'h5f == io_state_in_12 ? 8'h91 : _GEN_13406; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13408 = 8'h60 == io_state_in_12 ? 8'h4d : _GEN_13407; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13409 = 8'h61 == io_state_in_12 ? 8'h44 : _GEN_13408; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13410 = 8'h62 == io_state_in_12 ? 8'h5f : _GEN_13409; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13411 = 8'h63 == io_state_in_12 ? 8'h56 : _GEN_13410; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13412 = 8'h64 == io_state_in_12 ? 8'h69 : _GEN_13411; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13413 = 8'h65 == io_state_in_12 ? 8'h60 : _GEN_13412; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13414 = 8'h66 == io_state_in_12 ? 8'h7b : _GEN_13413; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13415 = 8'h67 == io_state_in_12 ? 8'h72 : _GEN_13414; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13416 = 8'h68 == io_state_in_12 ? 8'h5 : _GEN_13415; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13417 = 8'h69 == io_state_in_12 ? 8'hc : _GEN_13416; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13418 = 8'h6a == io_state_in_12 ? 8'h17 : _GEN_13417; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13419 = 8'h6b == io_state_in_12 ? 8'h1e : _GEN_13418; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13420 = 8'h6c == io_state_in_12 ? 8'h21 : _GEN_13419; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13421 = 8'h6d == io_state_in_12 ? 8'h28 : _GEN_13420; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13422 = 8'h6e == io_state_in_12 ? 8'h33 : _GEN_13421; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13423 = 8'h6f == io_state_in_12 ? 8'h3a : _GEN_13422; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13424 = 8'h70 == io_state_in_12 ? 8'hdd : _GEN_13423; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13425 = 8'h71 == io_state_in_12 ? 8'hd4 : _GEN_13424; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13426 = 8'h72 == io_state_in_12 ? 8'hcf : _GEN_13425; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13427 = 8'h73 == io_state_in_12 ? 8'hc6 : _GEN_13426; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13428 = 8'h74 == io_state_in_12 ? 8'hf9 : _GEN_13427; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13429 = 8'h75 == io_state_in_12 ? 8'hf0 : _GEN_13428; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13430 = 8'h76 == io_state_in_12 ? 8'heb : _GEN_13429; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13431 = 8'h77 == io_state_in_12 ? 8'he2 : _GEN_13430; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13432 = 8'h78 == io_state_in_12 ? 8'h95 : _GEN_13431; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13433 = 8'h79 == io_state_in_12 ? 8'h9c : _GEN_13432; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13434 = 8'h7a == io_state_in_12 ? 8'h87 : _GEN_13433; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13435 = 8'h7b == io_state_in_12 ? 8'h8e : _GEN_13434; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13436 = 8'h7c == io_state_in_12 ? 8'hb1 : _GEN_13435; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13437 = 8'h7d == io_state_in_12 ? 8'hb8 : _GEN_13436; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13438 = 8'h7e == io_state_in_12 ? 8'ha3 : _GEN_13437; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13439 = 8'h7f == io_state_in_12 ? 8'haa : _GEN_13438; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13440 = 8'h80 == io_state_in_12 ? 8'hec : _GEN_13439; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13441 = 8'h81 == io_state_in_12 ? 8'he5 : _GEN_13440; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13442 = 8'h82 == io_state_in_12 ? 8'hfe : _GEN_13441; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13443 = 8'h83 == io_state_in_12 ? 8'hf7 : _GEN_13442; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13444 = 8'h84 == io_state_in_12 ? 8'hc8 : _GEN_13443; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13445 = 8'h85 == io_state_in_12 ? 8'hc1 : _GEN_13444; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13446 = 8'h86 == io_state_in_12 ? 8'hda : _GEN_13445; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13447 = 8'h87 == io_state_in_12 ? 8'hd3 : _GEN_13446; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13448 = 8'h88 == io_state_in_12 ? 8'ha4 : _GEN_13447; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13449 = 8'h89 == io_state_in_12 ? 8'had : _GEN_13448; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13450 = 8'h8a == io_state_in_12 ? 8'hb6 : _GEN_13449; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13451 = 8'h8b == io_state_in_12 ? 8'hbf : _GEN_13450; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13452 = 8'h8c == io_state_in_12 ? 8'h80 : _GEN_13451; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13453 = 8'h8d == io_state_in_12 ? 8'h89 : _GEN_13452; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13454 = 8'h8e == io_state_in_12 ? 8'h92 : _GEN_13453; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13455 = 8'h8f == io_state_in_12 ? 8'h9b : _GEN_13454; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13456 = 8'h90 == io_state_in_12 ? 8'h7c : _GEN_13455; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13457 = 8'h91 == io_state_in_12 ? 8'h75 : _GEN_13456; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13458 = 8'h92 == io_state_in_12 ? 8'h6e : _GEN_13457; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13459 = 8'h93 == io_state_in_12 ? 8'h67 : _GEN_13458; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13460 = 8'h94 == io_state_in_12 ? 8'h58 : _GEN_13459; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13461 = 8'h95 == io_state_in_12 ? 8'h51 : _GEN_13460; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13462 = 8'h96 == io_state_in_12 ? 8'h4a : _GEN_13461; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13463 = 8'h97 == io_state_in_12 ? 8'h43 : _GEN_13462; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13464 = 8'h98 == io_state_in_12 ? 8'h34 : _GEN_13463; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13465 = 8'h99 == io_state_in_12 ? 8'h3d : _GEN_13464; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13466 = 8'h9a == io_state_in_12 ? 8'h26 : _GEN_13465; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13467 = 8'h9b == io_state_in_12 ? 8'h2f : _GEN_13466; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13468 = 8'h9c == io_state_in_12 ? 8'h10 : _GEN_13467; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13469 = 8'h9d == io_state_in_12 ? 8'h19 : _GEN_13468; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13470 = 8'h9e == io_state_in_12 ? 8'h2 : _GEN_13469; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13471 = 8'h9f == io_state_in_12 ? 8'hb : _GEN_13470; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13472 = 8'ha0 == io_state_in_12 ? 8'hd7 : _GEN_13471; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13473 = 8'ha1 == io_state_in_12 ? 8'hde : _GEN_13472; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13474 = 8'ha2 == io_state_in_12 ? 8'hc5 : _GEN_13473; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13475 = 8'ha3 == io_state_in_12 ? 8'hcc : _GEN_13474; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13476 = 8'ha4 == io_state_in_12 ? 8'hf3 : _GEN_13475; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13477 = 8'ha5 == io_state_in_12 ? 8'hfa : _GEN_13476; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13478 = 8'ha6 == io_state_in_12 ? 8'he1 : _GEN_13477; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13479 = 8'ha7 == io_state_in_12 ? 8'he8 : _GEN_13478; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13480 = 8'ha8 == io_state_in_12 ? 8'h9f : _GEN_13479; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13481 = 8'ha9 == io_state_in_12 ? 8'h96 : _GEN_13480; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13482 = 8'haa == io_state_in_12 ? 8'h8d : _GEN_13481; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13483 = 8'hab == io_state_in_12 ? 8'h84 : _GEN_13482; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13484 = 8'hac == io_state_in_12 ? 8'hbb : _GEN_13483; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13485 = 8'had == io_state_in_12 ? 8'hb2 : _GEN_13484; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13486 = 8'hae == io_state_in_12 ? 8'ha9 : _GEN_13485; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13487 = 8'haf == io_state_in_12 ? 8'ha0 : _GEN_13486; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13488 = 8'hb0 == io_state_in_12 ? 8'h47 : _GEN_13487; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13489 = 8'hb1 == io_state_in_12 ? 8'h4e : _GEN_13488; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13490 = 8'hb2 == io_state_in_12 ? 8'h55 : _GEN_13489; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13491 = 8'hb3 == io_state_in_12 ? 8'h5c : _GEN_13490; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13492 = 8'hb4 == io_state_in_12 ? 8'h63 : _GEN_13491; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13493 = 8'hb5 == io_state_in_12 ? 8'h6a : _GEN_13492; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13494 = 8'hb6 == io_state_in_12 ? 8'h71 : _GEN_13493; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13495 = 8'hb7 == io_state_in_12 ? 8'h78 : _GEN_13494; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13496 = 8'hb8 == io_state_in_12 ? 8'hf : _GEN_13495; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13497 = 8'hb9 == io_state_in_12 ? 8'h6 : _GEN_13496; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13498 = 8'hba == io_state_in_12 ? 8'h1d : _GEN_13497; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13499 = 8'hbb == io_state_in_12 ? 8'h14 : _GEN_13498; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13500 = 8'hbc == io_state_in_12 ? 8'h2b : _GEN_13499; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13501 = 8'hbd == io_state_in_12 ? 8'h22 : _GEN_13500; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13502 = 8'hbe == io_state_in_12 ? 8'h39 : _GEN_13501; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13503 = 8'hbf == io_state_in_12 ? 8'h30 : _GEN_13502; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13504 = 8'hc0 == io_state_in_12 ? 8'h9a : _GEN_13503; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13505 = 8'hc1 == io_state_in_12 ? 8'h93 : _GEN_13504; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13506 = 8'hc2 == io_state_in_12 ? 8'h88 : _GEN_13505; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13507 = 8'hc3 == io_state_in_12 ? 8'h81 : _GEN_13506; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13508 = 8'hc4 == io_state_in_12 ? 8'hbe : _GEN_13507; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13509 = 8'hc5 == io_state_in_12 ? 8'hb7 : _GEN_13508; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13510 = 8'hc6 == io_state_in_12 ? 8'hac : _GEN_13509; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13511 = 8'hc7 == io_state_in_12 ? 8'ha5 : _GEN_13510; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13512 = 8'hc8 == io_state_in_12 ? 8'hd2 : _GEN_13511; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13513 = 8'hc9 == io_state_in_12 ? 8'hdb : _GEN_13512; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13514 = 8'hca == io_state_in_12 ? 8'hc0 : _GEN_13513; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13515 = 8'hcb == io_state_in_12 ? 8'hc9 : _GEN_13514; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13516 = 8'hcc == io_state_in_12 ? 8'hf6 : _GEN_13515; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13517 = 8'hcd == io_state_in_12 ? 8'hff : _GEN_13516; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13518 = 8'hce == io_state_in_12 ? 8'he4 : _GEN_13517; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13519 = 8'hcf == io_state_in_12 ? 8'hed : _GEN_13518; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13520 = 8'hd0 == io_state_in_12 ? 8'ha : _GEN_13519; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13521 = 8'hd1 == io_state_in_12 ? 8'h3 : _GEN_13520; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13522 = 8'hd2 == io_state_in_12 ? 8'h18 : _GEN_13521; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13523 = 8'hd3 == io_state_in_12 ? 8'h11 : _GEN_13522; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13524 = 8'hd4 == io_state_in_12 ? 8'h2e : _GEN_13523; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13525 = 8'hd5 == io_state_in_12 ? 8'h27 : _GEN_13524; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13526 = 8'hd6 == io_state_in_12 ? 8'h3c : _GEN_13525; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13527 = 8'hd7 == io_state_in_12 ? 8'h35 : _GEN_13526; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13528 = 8'hd8 == io_state_in_12 ? 8'h42 : _GEN_13527; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13529 = 8'hd9 == io_state_in_12 ? 8'h4b : _GEN_13528; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13530 = 8'hda == io_state_in_12 ? 8'h50 : _GEN_13529; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13531 = 8'hdb == io_state_in_12 ? 8'h59 : _GEN_13530; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13532 = 8'hdc == io_state_in_12 ? 8'h66 : _GEN_13531; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13533 = 8'hdd == io_state_in_12 ? 8'h6f : _GEN_13532; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13534 = 8'hde == io_state_in_12 ? 8'h74 : _GEN_13533; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13535 = 8'hdf == io_state_in_12 ? 8'h7d : _GEN_13534; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13536 = 8'he0 == io_state_in_12 ? 8'ha1 : _GEN_13535; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13537 = 8'he1 == io_state_in_12 ? 8'ha8 : _GEN_13536; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13538 = 8'he2 == io_state_in_12 ? 8'hb3 : _GEN_13537; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13539 = 8'he3 == io_state_in_12 ? 8'hba : _GEN_13538; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13540 = 8'he4 == io_state_in_12 ? 8'h85 : _GEN_13539; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13541 = 8'he5 == io_state_in_12 ? 8'h8c : _GEN_13540; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13542 = 8'he6 == io_state_in_12 ? 8'h97 : _GEN_13541; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13543 = 8'he7 == io_state_in_12 ? 8'h9e : _GEN_13542; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13544 = 8'he8 == io_state_in_12 ? 8'he9 : _GEN_13543; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13545 = 8'he9 == io_state_in_12 ? 8'he0 : _GEN_13544; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13546 = 8'hea == io_state_in_12 ? 8'hfb : _GEN_13545; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13547 = 8'heb == io_state_in_12 ? 8'hf2 : _GEN_13546; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13548 = 8'hec == io_state_in_12 ? 8'hcd : _GEN_13547; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13549 = 8'hed == io_state_in_12 ? 8'hc4 : _GEN_13548; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13550 = 8'hee == io_state_in_12 ? 8'hdf : _GEN_13549; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13551 = 8'hef == io_state_in_12 ? 8'hd6 : _GEN_13550; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13552 = 8'hf0 == io_state_in_12 ? 8'h31 : _GEN_13551; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13553 = 8'hf1 == io_state_in_12 ? 8'h38 : _GEN_13552; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13554 = 8'hf2 == io_state_in_12 ? 8'h23 : _GEN_13553; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13555 = 8'hf3 == io_state_in_12 ? 8'h2a : _GEN_13554; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13556 = 8'hf4 == io_state_in_12 ? 8'h15 : _GEN_13555; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13557 = 8'hf5 == io_state_in_12 ? 8'h1c : _GEN_13556; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13558 = 8'hf6 == io_state_in_12 ? 8'h7 : _GEN_13557; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13559 = 8'hf7 == io_state_in_12 ? 8'he : _GEN_13558; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13560 = 8'hf8 == io_state_in_12 ? 8'h79 : _GEN_13559; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13561 = 8'hf9 == io_state_in_12 ? 8'h70 : _GEN_13560; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13562 = 8'hfa == io_state_in_12 ? 8'h6b : _GEN_13561; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13563 = 8'hfb == io_state_in_12 ? 8'h62 : _GEN_13562; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13564 = 8'hfc == io_state_in_12 ? 8'h5d : _GEN_13563; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13565 = 8'hfd == io_state_in_12 ? 8'h54 : _GEN_13564; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13566 = 8'hfe == io_state_in_12 ? 8'h4f : _GEN_13565; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13567 = 8'hff == io_state_in_12 ? 8'h46 : _GEN_13566; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13569 = 8'h1 == io_state_in_13 ? 8'he : 8'h0; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13570 = 8'h2 == io_state_in_13 ? 8'h1c : _GEN_13569; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13571 = 8'h3 == io_state_in_13 ? 8'h12 : _GEN_13570; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13572 = 8'h4 == io_state_in_13 ? 8'h38 : _GEN_13571; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13573 = 8'h5 == io_state_in_13 ? 8'h36 : _GEN_13572; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13574 = 8'h6 == io_state_in_13 ? 8'h24 : _GEN_13573; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13575 = 8'h7 == io_state_in_13 ? 8'h2a : _GEN_13574; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13576 = 8'h8 == io_state_in_13 ? 8'h70 : _GEN_13575; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13577 = 8'h9 == io_state_in_13 ? 8'h7e : _GEN_13576; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13578 = 8'ha == io_state_in_13 ? 8'h6c : _GEN_13577; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13579 = 8'hb == io_state_in_13 ? 8'h62 : _GEN_13578; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13580 = 8'hc == io_state_in_13 ? 8'h48 : _GEN_13579; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13581 = 8'hd == io_state_in_13 ? 8'h46 : _GEN_13580; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13582 = 8'he == io_state_in_13 ? 8'h54 : _GEN_13581; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13583 = 8'hf == io_state_in_13 ? 8'h5a : _GEN_13582; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13584 = 8'h10 == io_state_in_13 ? 8'he0 : _GEN_13583; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13585 = 8'h11 == io_state_in_13 ? 8'hee : _GEN_13584; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13586 = 8'h12 == io_state_in_13 ? 8'hfc : _GEN_13585; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13587 = 8'h13 == io_state_in_13 ? 8'hf2 : _GEN_13586; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13588 = 8'h14 == io_state_in_13 ? 8'hd8 : _GEN_13587; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13589 = 8'h15 == io_state_in_13 ? 8'hd6 : _GEN_13588; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13590 = 8'h16 == io_state_in_13 ? 8'hc4 : _GEN_13589; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13591 = 8'h17 == io_state_in_13 ? 8'hca : _GEN_13590; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13592 = 8'h18 == io_state_in_13 ? 8'h90 : _GEN_13591; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13593 = 8'h19 == io_state_in_13 ? 8'h9e : _GEN_13592; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13594 = 8'h1a == io_state_in_13 ? 8'h8c : _GEN_13593; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13595 = 8'h1b == io_state_in_13 ? 8'h82 : _GEN_13594; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13596 = 8'h1c == io_state_in_13 ? 8'ha8 : _GEN_13595; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13597 = 8'h1d == io_state_in_13 ? 8'ha6 : _GEN_13596; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13598 = 8'h1e == io_state_in_13 ? 8'hb4 : _GEN_13597; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13599 = 8'h1f == io_state_in_13 ? 8'hba : _GEN_13598; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13600 = 8'h20 == io_state_in_13 ? 8'hdb : _GEN_13599; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13601 = 8'h21 == io_state_in_13 ? 8'hd5 : _GEN_13600; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13602 = 8'h22 == io_state_in_13 ? 8'hc7 : _GEN_13601; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13603 = 8'h23 == io_state_in_13 ? 8'hc9 : _GEN_13602; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13604 = 8'h24 == io_state_in_13 ? 8'he3 : _GEN_13603; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13605 = 8'h25 == io_state_in_13 ? 8'hed : _GEN_13604; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13606 = 8'h26 == io_state_in_13 ? 8'hff : _GEN_13605; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13607 = 8'h27 == io_state_in_13 ? 8'hf1 : _GEN_13606; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13608 = 8'h28 == io_state_in_13 ? 8'hab : _GEN_13607; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13609 = 8'h29 == io_state_in_13 ? 8'ha5 : _GEN_13608; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13610 = 8'h2a == io_state_in_13 ? 8'hb7 : _GEN_13609; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13611 = 8'h2b == io_state_in_13 ? 8'hb9 : _GEN_13610; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13612 = 8'h2c == io_state_in_13 ? 8'h93 : _GEN_13611; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13613 = 8'h2d == io_state_in_13 ? 8'h9d : _GEN_13612; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13614 = 8'h2e == io_state_in_13 ? 8'h8f : _GEN_13613; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13615 = 8'h2f == io_state_in_13 ? 8'h81 : _GEN_13614; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13616 = 8'h30 == io_state_in_13 ? 8'h3b : _GEN_13615; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13617 = 8'h31 == io_state_in_13 ? 8'h35 : _GEN_13616; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13618 = 8'h32 == io_state_in_13 ? 8'h27 : _GEN_13617; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13619 = 8'h33 == io_state_in_13 ? 8'h29 : _GEN_13618; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13620 = 8'h34 == io_state_in_13 ? 8'h3 : _GEN_13619; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13621 = 8'h35 == io_state_in_13 ? 8'hd : _GEN_13620; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13622 = 8'h36 == io_state_in_13 ? 8'h1f : _GEN_13621; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13623 = 8'h37 == io_state_in_13 ? 8'h11 : _GEN_13622; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13624 = 8'h38 == io_state_in_13 ? 8'h4b : _GEN_13623; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13625 = 8'h39 == io_state_in_13 ? 8'h45 : _GEN_13624; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13626 = 8'h3a == io_state_in_13 ? 8'h57 : _GEN_13625; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13627 = 8'h3b == io_state_in_13 ? 8'h59 : _GEN_13626; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13628 = 8'h3c == io_state_in_13 ? 8'h73 : _GEN_13627; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13629 = 8'h3d == io_state_in_13 ? 8'h7d : _GEN_13628; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13630 = 8'h3e == io_state_in_13 ? 8'h6f : _GEN_13629; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13631 = 8'h3f == io_state_in_13 ? 8'h61 : _GEN_13630; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13632 = 8'h40 == io_state_in_13 ? 8'had : _GEN_13631; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13633 = 8'h41 == io_state_in_13 ? 8'ha3 : _GEN_13632; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13634 = 8'h42 == io_state_in_13 ? 8'hb1 : _GEN_13633; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13635 = 8'h43 == io_state_in_13 ? 8'hbf : _GEN_13634; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13636 = 8'h44 == io_state_in_13 ? 8'h95 : _GEN_13635; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13637 = 8'h45 == io_state_in_13 ? 8'h9b : _GEN_13636; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13638 = 8'h46 == io_state_in_13 ? 8'h89 : _GEN_13637; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13639 = 8'h47 == io_state_in_13 ? 8'h87 : _GEN_13638; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13640 = 8'h48 == io_state_in_13 ? 8'hdd : _GEN_13639; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13641 = 8'h49 == io_state_in_13 ? 8'hd3 : _GEN_13640; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13642 = 8'h4a == io_state_in_13 ? 8'hc1 : _GEN_13641; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13643 = 8'h4b == io_state_in_13 ? 8'hcf : _GEN_13642; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13644 = 8'h4c == io_state_in_13 ? 8'he5 : _GEN_13643; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13645 = 8'h4d == io_state_in_13 ? 8'heb : _GEN_13644; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13646 = 8'h4e == io_state_in_13 ? 8'hf9 : _GEN_13645; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13647 = 8'h4f == io_state_in_13 ? 8'hf7 : _GEN_13646; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13648 = 8'h50 == io_state_in_13 ? 8'h4d : _GEN_13647; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13649 = 8'h51 == io_state_in_13 ? 8'h43 : _GEN_13648; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13650 = 8'h52 == io_state_in_13 ? 8'h51 : _GEN_13649; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13651 = 8'h53 == io_state_in_13 ? 8'h5f : _GEN_13650; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13652 = 8'h54 == io_state_in_13 ? 8'h75 : _GEN_13651; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13653 = 8'h55 == io_state_in_13 ? 8'h7b : _GEN_13652; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13654 = 8'h56 == io_state_in_13 ? 8'h69 : _GEN_13653; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13655 = 8'h57 == io_state_in_13 ? 8'h67 : _GEN_13654; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13656 = 8'h58 == io_state_in_13 ? 8'h3d : _GEN_13655; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13657 = 8'h59 == io_state_in_13 ? 8'h33 : _GEN_13656; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13658 = 8'h5a == io_state_in_13 ? 8'h21 : _GEN_13657; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13659 = 8'h5b == io_state_in_13 ? 8'h2f : _GEN_13658; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13660 = 8'h5c == io_state_in_13 ? 8'h5 : _GEN_13659; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13661 = 8'h5d == io_state_in_13 ? 8'hb : _GEN_13660; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13662 = 8'h5e == io_state_in_13 ? 8'h19 : _GEN_13661; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13663 = 8'h5f == io_state_in_13 ? 8'h17 : _GEN_13662; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13664 = 8'h60 == io_state_in_13 ? 8'h76 : _GEN_13663; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13665 = 8'h61 == io_state_in_13 ? 8'h78 : _GEN_13664; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13666 = 8'h62 == io_state_in_13 ? 8'h6a : _GEN_13665; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13667 = 8'h63 == io_state_in_13 ? 8'h64 : _GEN_13666; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13668 = 8'h64 == io_state_in_13 ? 8'h4e : _GEN_13667; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13669 = 8'h65 == io_state_in_13 ? 8'h40 : _GEN_13668; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13670 = 8'h66 == io_state_in_13 ? 8'h52 : _GEN_13669; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13671 = 8'h67 == io_state_in_13 ? 8'h5c : _GEN_13670; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13672 = 8'h68 == io_state_in_13 ? 8'h6 : _GEN_13671; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13673 = 8'h69 == io_state_in_13 ? 8'h8 : _GEN_13672; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13674 = 8'h6a == io_state_in_13 ? 8'h1a : _GEN_13673; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13675 = 8'h6b == io_state_in_13 ? 8'h14 : _GEN_13674; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13676 = 8'h6c == io_state_in_13 ? 8'h3e : _GEN_13675; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13677 = 8'h6d == io_state_in_13 ? 8'h30 : _GEN_13676; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13678 = 8'h6e == io_state_in_13 ? 8'h22 : _GEN_13677; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13679 = 8'h6f == io_state_in_13 ? 8'h2c : _GEN_13678; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13680 = 8'h70 == io_state_in_13 ? 8'h96 : _GEN_13679; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13681 = 8'h71 == io_state_in_13 ? 8'h98 : _GEN_13680; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13682 = 8'h72 == io_state_in_13 ? 8'h8a : _GEN_13681; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13683 = 8'h73 == io_state_in_13 ? 8'h84 : _GEN_13682; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13684 = 8'h74 == io_state_in_13 ? 8'hae : _GEN_13683; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13685 = 8'h75 == io_state_in_13 ? 8'ha0 : _GEN_13684; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13686 = 8'h76 == io_state_in_13 ? 8'hb2 : _GEN_13685; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13687 = 8'h77 == io_state_in_13 ? 8'hbc : _GEN_13686; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13688 = 8'h78 == io_state_in_13 ? 8'he6 : _GEN_13687; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13689 = 8'h79 == io_state_in_13 ? 8'he8 : _GEN_13688; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13690 = 8'h7a == io_state_in_13 ? 8'hfa : _GEN_13689; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13691 = 8'h7b == io_state_in_13 ? 8'hf4 : _GEN_13690; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13692 = 8'h7c == io_state_in_13 ? 8'hde : _GEN_13691; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13693 = 8'h7d == io_state_in_13 ? 8'hd0 : _GEN_13692; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13694 = 8'h7e == io_state_in_13 ? 8'hc2 : _GEN_13693; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13695 = 8'h7f == io_state_in_13 ? 8'hcc : _GEN_13694; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13696 = 8'h80 == io_state_in_13 ? 8'h41 : _GEN_13695; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13697 = 8'h81 == io_state_in_13 ? 8'h4f : _GEN_13696; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13698 = 8'h82 == io_state_in_13 ? 8'h5d : _GEN_13697; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13699 = 8'h83 == io_state_in_13 ? 8'h53 : _GEN_13698; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13700 = 8'h84 == io_state_in_13 ? 8'h79 : _GEN_13699; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13701 = 8'h85 == io_state_in_13 ? 8'h77 : _GEN_13700; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13702 = 8'h86 == io_state_in_13 ? 8'h65 : _GEN_13701; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13703 = 8'h87 == io_state_in_13 ? 8'h6b : _GEN_13702; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13704 = 8'h88 == io_state_in_13 ? 8'h31 : _GEN_13703; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13705 = 8'h89 == io_state_in_13 ? 8'h3f : _GEN_13704; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13706 = 8'h8a == io_state_in_13 ? 8'h2d : _GEN_13705; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13707 = 8'h8b == io_state_in_13 ? 8'h23 : _GEN_13706; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13708 = 8'h8c == io_state_in_13 ? 8'h9 : _GEN_13707; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13709 = 8'h8d == io_state_in_13 ? 8'h7 : _GEN_13708; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13710 = 8'h8e == io_state_in_13 ? 8'h15 : _GEN_13709; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13711 = 8'h8f == io_state_in_13 ? 8'h1b : _GEN_13710; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13712 = 8'h90 == io_state_in_13 ? 8'ha1 : _GEN_13711; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13713 = 8'h91 == io_state_in_13 ? 8'haf : _GEN_13712; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13714 = 8'h92 == io_state_in_13 ? 8'hbd : _GEN_13713; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13715 = 8'h93 == io_state_in_13 ? 8'hb3 : _GEN_13714; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13716 = 8'h94 == io_state_in_13 ? 8'h99 : _GEN_13715; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13717 = 8'h95 == io_state_in_13 ? 8'h97 : _GEN_13716; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13718 = 8'h96 == io_state_in_13 ? 8'h85 : _GEN_13717; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13719 = 8'h97 == io_state_in_13 ? 8'h8b : _GEN_13718; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13720 = 8'h98 == io_state_in_13 ? 8'hd1 : _GEN_13719; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13721 = 8'h99 == io_state_in_13 ? 8'hdf : _GEN_13720; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13722 = 8'h9a == io_state_in_13 ? 8'hcd : _GEN_13721; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13723 = 8'h9b == io_state_in_13 ? 8'hc3 : _GEN_13722; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13724 = 8'h9c == io_state_in_13 ? 8'he9 : _GEN_13723; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13725 = 8'h9d == io_state_in_13 ? 8'he7 : _GEN_13724; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13726 = 8'h9e == io_state_in_13 ? 8'hf5 : _GEN_13725; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13727 = 8'h9f == io_state_in_13 ? 8'hfb : _GEN_13726; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13728 = 8'ha0 == io_state_in_13 ? 8'h9a : _GEN_13727; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13729 = 8'ha1 == io_state_in_13 ? 8'h94 : _GEN_13728; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13730 = 8'ha2 == io_state_in_13 ? 8'h86 : _GEN_13729; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13731 = 8'ha3 == io_state_in_13 ? 8'h88 : _GEN_13730; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13732 = 8'ha4 == io_state_in_13 ? 8'ha2 : _GEN_13731; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13733 = 8'ha5 == io_state_in_13 ? 8'hac : _GEN_13732; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13734 = 8'ha6 == io_state_in_13 ? 8'hbe : _GEN_13733; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13735 = 8'ha7 == io_state_in_13 ? 8'hb0 : _GEN_13734; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13736 = 8'ha8 == io_state_in_13 ? 8'hea : _GEN_13735; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13737 = 8'ha9 == io_state_in_13 ? 8'he4 : _GEN_13736; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13738 = 8'haa == io_state_in_13 ? 8'hf6 : _GEN_13737; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13739 = 8'hab == io_state_in_13 ? 8'hf8 : _GEN_13738; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13740 = 8'hac == io_state_in_13 ? 8'hd2 : _GEN_13739; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13741 = 8'had == io_state_in_13 ? 8'hdc : _GEN_13740; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13742 = 8'hae == io_state_in_13 ? 8'hce : _GEN_13741; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13743 = 8'haf == io_state_in_13 ? 8'hc0 : _GEN_13742; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13744 = 8'hb0 == io_state_in_13 ? 8'h7a : _GEN_13743; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13745 = 8'hb1 == io_state_in_13 ? 8'h74 : _GEN_13744; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13746 = 8'hb2 == io_state_in_13 ? 8'h66 : _GEN_13745; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13747 = 8'hb3 == io_state_in_13 ? 8'h68 : _GEN_13746; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13748 = 8'hb4 == io_state_in_13 ? 8'h42 : _GEN_13747; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13749 = 8'hb5 == io_state_in_13 ? 8'h4c : _GEN_13748; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13750 = 8'hb6 == io_state_in_13 ? 8'h5e : _GEN_13749; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13751 = 8'hb7 == io_state_in_13 ? 8'h50 : _GEN_13750; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13752 = 8'hb8 == io_state_in_13 ? 8'ha : _GEN_13751; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13753 = 8'hb9 == io_state_in_13 ? 8'h4 : _GEN_13752; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13754 = 8'hba == io_state_in_13 ? 8'h16 : _GEN_13753; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13755 = 8'hbb == io_state_in_13 ? 8'h18 : _GEN_13754; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13756 = 8'hbc == io_state_in_13 ? 8'h32 : _GEN_13755; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13757 = 8'hbd == io_state_in_13 ? 8'h3c : _GEN_13756; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13758 = 8'hbe == io_state_in_13 ? 8'h2e : _GEN_13757; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13759 = 8'hbf == io_state_in_13 ? 8'h20 : _GEN_13758; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13760 = 8'hc0 == io_state_in_13 ? 8'hec : _GEN_13759; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13761 = 8'hc1 == io_state_in_13 ? 8'he2 : _GEN_13760; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13762 = 8'hc2 == io_state_in_13 ? 8'hf0 : _GEN_13761; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13763 = 8'hc3 == io_state_in_13 ? 8'hfe : _GEN_13762; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13764 = 8'hc4 == io_state_in_13 ? 8'hd4 : _GEN_13763; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13765 = 8'hc5 == io_state_in_13 ? 8'hda : _GEN_13764; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13766 = 8'hc6 == io_state_in_13 ? 8'hc8 : _GEN_13765; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13767 = 8'hc7 == io_state_in_13 ? 8'hc6 : _GEN_13766; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13768 = 8'hc8 == io_state_in_13 ? 8'h9c : _GEN_13767; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13769 = 8'hc9 == io_state_in_13 ? 8'h92 : _GEN_13768; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13770 = 8'hca == io_state_in_13 ? 8'h80 : _GEN_13769; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13771 = 8'hcb == io_state_in_13 ? 8'h8e : _GEN_13770; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13772 = 8'hcc == io_state_in_13 ? 8'ha4 : _GEN_13771; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13773 = 8'hcd == io_state_in_13 ? 8'haa : _GEN_13772; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13774 = 8'hce == io_state_in_13 ? 8'hb8 : _GEN_13773; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13775 = 8'hcf == io_state_in_13 ? 8'hb6 : _GEN_13774; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13776 = 8'hd0 == io_state_in_13 ? 8'hc : _GEN_13775; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13777 = 8'hd1 == io_state_in_13 ? 8'h2 : _GEN_13776; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13778 = 8'hd2 == io_state_in_13 ? 8'h10 : _GEN_13777; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13779 = 8'hd3 == io_state_in_13 ? 8'h1e : _GEN_13778; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13780 = 8'hd4 == io_state_in_13 ? 8'h34 : _GEN_13779; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13781 = 8'hd5 == io_state_in_13 ? 8'h3a : _GEN_13780; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13782 = 8'hd6 == io_state_in_13 ? 8'h28 : _GEN_13781; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13783 = 8'hd7 == io_state_in_13 ? 8'h26 : _GEN_13782; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13784 = 8'hd8 == io_state_in_13 ? 8'h7c : _GEN_13783; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13785 = 8'hd9 == io_state_in_13 ? 8'h72 : _GEN_13784; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13786 = 8'hda == io_state_in_13 ? 8'h60 : _GEN_13785; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13787 = 8'hdb == io_state_in_13 ? 8'h6e : _GEN_13786; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13788 = 8'hdc == io_state_in_13 ? 8'h44 : _GEN_13787; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13789 = 8'hdd == io_state_in_13 ? 8'h4a : _GEN_13788; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13790 = 8'hde == io_state_in_13 ? 8'h58 : _GEN_13789; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13791 = 8'hdf == io_state_in_13 ? 8'h56 : _GEN_13790; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13792 = 8'he0 == io_state_in_13 ? 8'h37 : _GEN_13791; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13793 = 8'he1 == io_state_in_13 ? 8'h39 : _GEN_13792; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13794 = 8'he2 == io_state_in_13 ? 8'h2b : _GEN_13793; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13795 = 8'he3 == io_state_in_13 ? 8'h25 : _GEN_13794; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13796 = 8'he4 == io_state_in_13 ? 8'hf : _GEN_13795; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13797 = 8'he5 == io_state_in_13 ? 8'h1 : _GEN_13796; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13798 = 8'he6 == io_state_in_13 ? 8'h13 : _GEN_13797; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13799 = 8'he7 == io_state_in_13 ? 8'h1d : _GEN_13798; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13800 = 8'he8 == io_state_in_13 ? 8'h47 : _GEN_13799; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13801 = 8'he9 == io_state_in_13 ? 8'h49 : _GEN_13800; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13802 = 8'hea == io_state_in_13 ? 8'h5b : _GEN_13801; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13803 = 8'heb == io_state_in_13 ? 8'h55 : _GEN_13802; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13804 = 8'hec == io_state_in_13 ? 8'h7f : _GEN_13803; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13805 = 8'hed == io_state_in_13 ? 8'h71 : _GEN_13804; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13806 = 8'hee == io_state_in_13 ? 8'h63 : _GEN_13805; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13807 = 8'hef == io_state_in_13 ? 8'h6d : _GEN_13806; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13808 = 8'hf0 == io_state_in_13 ? 8'hd7 : _GEN_13807; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13809 = 8'hf1 == io_state_in_13 ? 8'hd9 : _GEN_13808; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13810 = 8'hf2 == io_state_in_13 ? 8'hcb : _GEN_13809; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13811 = 8'hf3 == io_state_in_13 ? 8'hc5 : _GEN_13810; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13812 = 8'hf4 == io_state_in_13 ? 8'hef : _GEN_13811; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13813 = 8'hf5 == io_state_in_13 ? 8'he1 : _GEN_13812; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13814 = 8'hf6 == io_state_in_13 ? 8'hf3 : _GEN_13813; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13815 = 8'hf7 == io_state_in_13 ? 8'hfd : _GEN_13814; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13816 = 8'hf8 == io_state_in_13 ? 8'ha7 : _GEN_13815; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13817 = 8'hf9 == io_state_in_13 ? 8'ha9 : _GEN_13816; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13818 = 8'hfa == io_state_in_13 ? 8'hbb : _GEN_13817; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13819 = 8'hfb == io_state_in_13 ? 8'hb5 : _GEN_13818; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13820 = 8'hfc == io_state_in_13 ? 8'h9f : _GEN_13819; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13821 = 8'hfd == io_state_in_13 ? 8'h91 : _GEN_13820; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13822 = 8'hfe == io_state_in_13 ? 8'h83 : _GEN_13821; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _GEN_13823 = 8'hff == io_state_in_13 ? 8'h8d : _GEN_13822; // @[InvMixColumns.scala 142:{43,43}]
  wire [7:0] _tmp_state_13_T = _GEN_13567 ^ _GEN_13823; // @[InvMixColumns.scala 142:43]
  wire [7:0] _GEN_13825 = 8'h1 == io_state_in_14 ? 8'hb : 8'h0; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13826 = 8'h2 == io_state_in_14 ? 8'h16 : _GEN_13825; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13827 = 8'h3 == io_state_in_14 ? 8'h1d : _GEN_13826; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13828 = 8'h4 == io_state_in_14 ? 8'h2c : _GEN_13827; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13829 = 8'h5 == io_state_in_14 ? 8'h27 : _GEN_13828; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13830 = 8'h6 == io_state_in_14 ? 8'h3a : _GEN_13829; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13831 = 8'h7 == io_state_in_14 ? 8'h31 : _GEN_13830; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13832 = 8'h8 == io_state_in_14 ? 8'h58 : _GEN_13831; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13833 = 8'h9 == io_state_in_14 ? 8'h53 : _GEN_13832; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13834 = 8'ha == io_state_in_14 ? 8'h4e : _GEN_13833; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13835 = 8'hb == io_state_in_14 ? 8'h45 : _GEN_13834; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13836 = 8'hc == io_state_in_14 ? 8'h74 : _GEN_13835; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13837 = 8'hd == io_state_in_14 ? 8'h7f : _GEN_13836; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13838 = 8'he == io_state_in_14 ? 8'h62 : _GEN_13837; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13839 = 8'hf == io_state_in_14 ? 8'h69 : _GEN_13838; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13840 = 8'h10 == io_state_in_14 ? 8'hb0 : _GEN_13839; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13841 = 8'h11 == io_state_in_14 ? 8'hbb : _GEN_13840; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13842 = 8'h12 == io_state_in_14 ? 8'ha6 : _GEN_13841; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13843 = 8'h13 == io_state_in_14 ? 8'had : _GEN_13842; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13844 = 8'h14 == io_state_in_14 ? 8'h9c : _GEN_13843; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13845 = 8'h15 == io_state_in_14 ? 8'h97 : _GEN_13844; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13846 = 8'h16 == io_state_in_14 ? 8'h8a : _GEN_13845; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13847 = 8'h17 == io_state_in_14 ? 8'h81 : _GEN_13846; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13848 = 8'h18 == io_state_in_14 ? 8'he8 : _GEN_13847; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13849 = 8'h19 == io_state_in_14 ? 8'he3 : _GEN_13848; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13850 = 8'h1a == io_state_in_14 ? 8'hfe : _GEN_13849; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13851 = 8'h1b == io_state_in_14 ? 8'hf5 : _GEN_13850; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13852 = 8'h1c == io_state_in_14 ? 8'hc4 : _GEN_13851; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13853 = 8'h1d == io_state_in_14 ? 8'hcf : _GEN_13852; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13854 = 8'h1e == io_state_in_14 ? 8'hd2 : _GEN_13853; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13855 = 8'h1f == io_state_in_14 ? 8'hd9 : _GEN_13854; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13856 = 8'h20 == io_state_in_14 ? 8'h7b : _GEN_13855; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13857 = 8'h21 == io_state_in_14 ? 8'h70 : _GEN_13856; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13858 = 8'h22 == io_state_in_14 ? 8'h6d : _GEN_13857; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13859 = 8'h23 == io_state_in_14 ? 8'h66 : _GEN_13858; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13860 = 8'h24 == io_state_in_14 ? 8'h57 : _GEN_13859; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13861 = 8'h25 == io_state_in_14 ? 8'h5c : _GEN_13860; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13862 = 8'h26 == io_state_in_14 ? 8'h41 : _GEN_13861; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13863 = 8'h27 == io_state_in_14 ? 8'h4a : _GEN_13862; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13864 = 8'h28 == io_state_in_14 ? 8'h23 : _GEN_13863; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13865 = 8'h29 == io_state_in_14 ? 8'h28 : _GEN_13864; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13866 = 8'h2a == io_state_in_14 ? 8'h35 : _GEN_13865; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13867 = 8'h2b == io_state_in_14 ? 8'h3e : _GEN_13866; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13868 = 8'h2c == io_state_in_14 ? 8'hf : _GEN_13867; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13869 = 8'h2d == io_state_in_14 ? 8'h4 : _GEN_13868; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13870 = 8'h2e == io_state_in_14 ? 8'h19 : _GEN_13869; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13871 = 8'h2f == io_state_in_14 ? 8'h12 : _GEN_13870; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13872 = 8'h30 == io_state_in_14 ? 8'hcb : _GEN_13871; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13873 = 8'h31 == io_state_in_14 ? 8'hc0 : _GEN_13872; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13874 = 8'h32 == io_state_in_14 ? 8'hdd : _GEN_13873; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13875 = 8'h33 == io_state_in_14 ? 8'hd6 : _GEN_13874; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13876 = 8'h34 == io_state_in_14 ? 8'he7 : _GEN_13875; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13877 = 8'h35 == io_state_in_14 ? 8'hec : _GEN_13876; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13878 = 8'h36 == io_state_in_14 ? 8'hf1 : _GEN_13877; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13879 = 8'h37 == io_state_in_14 ? 8'hfa : _GEN_13878; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13880 = 8'h38 == io_state_in_14 ? 8'h93 : _GEN_13879; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13881 = 8'h39 == io_state_in_14 ? 8'h98 : _GEN_13880; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13882 = 8'h3a == io_state_in_14 ? 8'h85 : _GEN_13881; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13883 = 8'h3b == io_state_in_14 ? 8'h8e : _GEN_13882; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13884 = 8'h3c == io_state_in_14 ? 8'hbf : _GEN_13883; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13885 = 8'h3d == io_state_in_14 ? 8'hb4 : _GEN_13884; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13886 = 8'h3e == io_state_in_14 ? 8'ha9 : _GEN_13885; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13887 = 8'h3f == io_state_in_14 ? 8'ha2 : _GEN_13886; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13888 = 8'h40 == io_state_in_14 ? 8'hf6 : _GEN_13887; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13889 = 8'h41 == io_state_in_14 ? 8'hfd : _GEN_13888; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13890 = 8'h42 == io_state_in_14 ? 8'he0 : _GEN_13889; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13891 = 8'h43 == io_state_in_14 ? 8'heb : _GEN_13890; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13892 = 8'h44 == io_state_in_14 ? 8'hda : _GEN_13891; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13893 = 8'h45 == io_state_in_14 ? 8'hd1 : _GEN_13892; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13894 = 8'h46 == io_state_in_14 ? 8'hcc : _GEN_13893; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13895 = 8'h47 == io_state_in_14 ? 8'hc7 : _GEN_13894; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13896 = 8'h48 == io_state_in_14 ? 8'hae : _GEN_13895; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13897 = 8'h49 == io_state_in_14 ? 8'ha5 : _GEN_13896; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13898 = 8'h4a == io_state_in_14 ? 8'hb8 : _GEN_13897; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13899 = 8'h4b == io_state_in_14 ? 8'hb3 : _GEN_13898; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13900 = 8'h4c == io_state_in_14 ? 8'h82 : _GEN_13899; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13901 = 8'h4d == io_state_in_14 ? 8'h89 : _GEN_13900; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13902 = 8'h4e == io_state_in_14 ? 8'h94 : _GEN_13901; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13903 = 8'h4f == io_state_in_14 ? 8'h9f : _GEN_13902; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13904 = 8'h50 == io_state_in_14 ? 8'h46 : _GEN_13903; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13905 = 8'h51 == io_state_in_14 ? 8'h4d : _GEN_13904; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13906 = 8'h52 == io_state_in_14 ? 8'h50 : _GEN_13905; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13907 = 8'h53 == io_state_in_14 ? 8'h5b : _GEN_13906; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13908 = 8'h54 == io_state_in_14 ? 8'h6a : _GEN_13907; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13909 = 8'h55 == io_state_in_14 ? 8'h61 : _GEN_13908; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13910 = 8'h56 == io_state_in_14 ? 8'h7c : _GEN_13909; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13911 = 8'h57 == io_state_in_14 ? 8'h77 : _GEN_13910; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13912 = 8'h58 == io_state_in_14 ? 8'h1e : _GEN_13911; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13913 = 8'h59 == io_state_in_14 ? 8'h15 : _GEN_13912; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13914 = 8'h5a == io_state_in_14 ? 8'h8 : _GEN_13913; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13915 = 8'h5b == io_state_in_14 ? 8'h3 : _GEN_13914; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13916 = 8'h5c == io_state_in_14 ? 8'h32 : _GEN_13915; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13917 = 8'h5d == io_state_in_14 ? 8'h39 : _GEN_13916; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13918 = 8'h5e == io_state_in_14 ? 8'h24 : _GEN_13917; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13919 = 8'h5f == io_state_in_14 ? 8'h2f : _GEN_13918; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13920 = 8'h60 == io_state_in_14 ? 8'h8d : _GEN_13919; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13921 = 8'h61 == io_state_in_14 ? 8'h86 : _GEN_13920; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13922 = 8'h62 == io_state_in_14 ? 8'h9b : _GEN_13921; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13923 = 8'h63 == io_state_in_14 ? 8'h90 : _GEN_13922; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13924 = 8'h64 == io_state_in_14 ? 8'ha1 : _GEN_13923; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13925 = 8'h65 == io_state_in_14 ? 8'haa : _GEN_13924; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13926 = 8'h66 == io_state_in_14 ? 8'hb7 : _GEN_13925; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13927 = 8'h67 == io_state_in_14 ? 8'hbc : _GEN_13926; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13928 = 8'h68 == io_state_in_14 ? 8'hd5 : _GEN_13927; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13929 = 8'h69 == io_state_in_14 ? 8'hde : _GEN_13928; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13930 = 8'h6a == io_state_in_14 ? 8'hc3 : _GEN_13929; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13931 = 8'h6b == io_state_in_14 ? 8'hc8 : _GEN_13930; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13932 = 8'h6c == io_state_in_14 ? 8'hf9 : _GEN_13931; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13933 = 8'h6d == io_state_in_14 ? 8'hf2 : _GEN_13932; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13934 = 8'h6e == io_state_in_14 ? 8'hef : _GEN_13933; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13935 = 8'h6f == io_state_in_14 ? 8'he4 : _GEN_13934; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13936 = 8'h70 == io_state_in_14 ? 8'h3d : _GEN_13935; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13937 = 8'h71 == io_state_in_14 ? 8'h36 : _GEN_13936; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13938 = 8'h72 == io_state_in_14 ? 8'h2b : _GEN_13937; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13939 = 8'h73 == io_state_in_14 ? 8'h20 : _GEN_13938; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13940 = 8'h74 == io_state_in_14 ? 8'h11 : _GEN_13939; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13941 = 8'h75 == io_state_in_14 ? 8'h1a : _GEN_13940; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13942 = 8'h76 == io_state_in_14 ? 8'h7 : _GEN_13941; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13943 = 8'h77 == io_state_in_14 ? 8'hc : _GEN_13942; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13944 = 8'h78 == io_state_in_14 ? 8'h65 : _GEN_13943; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13945 = 8'h79 == io_state_in_14 ? 8'h6e : _GEN_13944; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13946 = 8'h7a == io_state_in_14 ? 8'h73 : _GEN_13945; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13947 = 8'h7b == io_state_in_14 ? 8'h78 : _GEN_13946; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13948 = 8'h7c == io_state_in_14 ? 8'h49 : _GEN_13947; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13949 = 8'h7d == io_state_in_14 ? 8'h42 : _GEN_13948; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13950 = 8'h7e == io_state_in_14 ? 8'h5f : _GEN_13949; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13951 = 8'h7f == io_state_in_14 ? 8'h54 : _GEN_13950; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13952 = 8'h80 == io_state_in_14 ? 8'hf7 : _GEN_13951; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13953 = 8'h81 == io_state_in_14 ? 8'hfc : _GEN_13952; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13954 = 8'h82 == io_state_in_14 ? 8'he1 : _GEN_13953; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13955 = 8'h83 == io_state_in_14 ? 8'hea : _GEN_13954; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13956 = 8'h84 == io_state_in_14 ? 8'hdb : _GEN_13955; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13957 = 8'h85 == io_state_in_14 ? 8'hd0 : _GEN_13956; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13958 = 8'h86 == io_state_in_14 ? 8'hcd : _GEN_13957; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13959 = 8'h87 == io_state_in_14 ? 8'hc6 : _GEN_13958; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13960 = 8'h88 == io_state_in_14 ? 8'haf : _GEN_13959; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13961 = 8'h89 == io_state_in_14 ? 8'ha4 : _GEN_13960; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13962 = 8'h8a == io_state_in_14 ? 8'hb9 : _GEN_13961; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13963 = 8'h8b == io_state_in_14 ? 8'hb2 : _GEN_13962; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13964 = 8'h8c == io_state_in_14 ? 8'h83 : _GEN_13963; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13965 = 8'h8d == io_state_in_14 ? 8'h88 : _GEN_13964; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13966 = 8'h8e == io_state_in_14 ? 8'h95 : _GEN_13965; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13967 = 8'h8f == io_state_in_14 ? 8'h9e : _GEN_13966; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13968 = 8'h90 == io_state_in_14 ? 8'h47 : _GEN_13967; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13969 = 8'h91 == io_state_in_14 ? 8'h4c : _GEN_13968; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13970 = 8'h92 == io_state_in_14 ? 8'h51 : _GEN_13969; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13971 = 8'h93 == io_state_in_14 ? 8'h5a : _GEN_13970; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13972 = 8'h94 == io_state_in_14 ? 8'h6b : _GEN_13971; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13973 = 8'h95 == io_state_in_14 ? 8'h60 : _GEN_13972; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13974 = 8'h96 == io_state_in_14 ? 8'h7d : _GEN_13973; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13975 = 8'h97 == io_state_in_14 ? 8'h76 : _GEN_13974; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13976 = 8'h98 == io_state_in_14 ? 8'h1f : _GEN_13975; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13977 = 8'h99 == io_state_in_14 ? 8'h14 : _GEN_13976; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13978 = 8'h9a == io_state_in_14 ? 8'h9 : _GEN_13977; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13979 = 8'h9b == io_state_in_14 ? 8'h2 : _GEN_13978; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13980 = 8'h9c == io_state_in_14 ? 8'h33 : _GEN_13979; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13981 = 8'h9d == io_state_in_14 ? 8'h38 : _GEN_13980; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13982 = 8'h9e == io_state_in_14 ? 8'h25 : _GEN_13981; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13983 = 8'h9f == io_state_in_14 ? 8'h2e : _GEN_13982; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13984 = 8'ha0 == io_state_in_14 ? 8'h8c : _GEN_13983; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13985 = 8'ha1 == io_state_in_14 ? 8'h87 : _GEN_13984; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13986 = 8'ha2 == io_state_in_14 ? 8'h9a : _GEN_13985; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13987 = 8'ha3 == io_state_in_14 ? 8'h91 : _GEN_13986; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13988 = 8'ha4 == io_state_in_14 ? 8'ha0 : _GEN_13987; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13989 = 8'ha5 == io_state_in_14 ? 8'hab : _GEN_13988; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13990 = 8'ha6 == io_state_in_14 ? 8'hb6 : _GEN_13989; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13991 = 8'ha7 == io_state_in_14 ? 8'hbd : _GEN_13990; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13992 = 8'ha8 == io_state_in_14 ? 8'hd4 : _GEN_13991; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13993 = 8'ha9 == io_state_in_14 ? 8'hdf : _GEN_13992; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13994 = 8'haa == io_state_in_14 ? 8'hc2 : _GEN_13993; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13995 = 8'hab == io_state_in_14 ? 8'hc9 : _GEN_13994; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13996 = 8'hac == io_state_in_14 ? 8'hf8 : _GEN_13995; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13997 = 8'had == io_state_in_14 ? 8'hf3 : _GEN_13996; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13998 = 8'hae == io_state_in_14 ? 8'hee : _GEN_13997; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_13999 = 8'haf == io_state_in_14 ? 8'he5 : _GEN_13998; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14000 = 8'hb0 == io_state_in_14 ? 8'h3c : _GEN_13999; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14001 = 8'hb1 == io_state_in_14 ? 8'h37 : _GEN_14000; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14002 = 8'hb2 == io_state_in_14 ? 8'h2a : _GEN_14001; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14003 = 8'hb3 == io_state_in_14 ? 8'h21 : _GEN_14002; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14004 = 8'hb4 == io_state_in_14 ? 8'h10 : _GEN_14003; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14005 = 8'hb5 == io_state_in_14 ? 8'h1b : _GEN_14004; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14006 = 8'hb6 == io_state_in_14 ? 8'h6 : _GEN_14005; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14007 = 8'hb7 == io_state_in_14 ? 8'hd : _GEN_14006; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14008 = 8'hb8 == io_state_in_14 ? 8'h64 : _GEN_14007; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14009 = 8'hb9 == io_state_in_14 ? 8'h6f : _GEN_14008; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14010 = 8'hba == io_state_in_14 ? 8'h72 : _GEN_14009; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14011 = 8'hbb == io_state_in_14 ? 8'h79 : _GEN_14010; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14012 = 8'hbc == io_state_in_14 ? 8'h48 : _GEN_14011; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14013 = 8'hbd == io_state_in_14 ? 8'h43 : _GEN_14012; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14014 = 8'hbe == io_state_in_14 ? 8'h5e : _GEN_14013; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14015 = 8'hbf == io_state_in_14 ? 8'h55 : _GEN_14014; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14016 = 8'hc0 == io_state_in_14 ? 8'h1 : _GEN_14015; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14017 = 8'hc1 == io_state_in_14 ? 8'ha : _GEN_14016; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14018 = 8'hc2 == io_state_in_14 ? 8'h17 : _GEN_14017; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14019 = 8'hc3 == io_state_in_14 ? 8'h1c : _GEN_14018; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14020 = 8'hc4 == io_state_in_14 ? 8'h2d : _GEN_14019; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14021 = 8'hc5 == io_state_in_14 ? 8'h26 : _GEN_14020; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14022 = 8'hc6 == io_state_in_14 ? 8'h3b : _GEN_14021; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14023 = 8'hc7 == io_state_in_14 ? 8'h30 : _GEN_14022; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14024 = 8'hc8 == io_state_in_14 ? 8'h59 : _GEN_14023; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14025 = 8'hc9 == io_state_in_14 ? 8'h52 : _GEN_14024; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14026 = 8'hca == io_state_in_14 ? 8'h4f : _GEN_14025; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14027 = 8'hcb == io_state_in_14 ? 8'h44 : _GEN_14026; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14028 = 8'hcc == io_state_in_14 ? 8'h75 : _GEN_14027; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14029 = 8'hcd == io_state_in_14 ? 8'h7e : _GEN_14028; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14030 = 8'hce == io_state_in_14 ? 8'h63 : _GEN_14029; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14031 = 8'hcf == io_state_in_14 ? 8'h68 : _GEN_14030; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14032 = 8'hd0 == io_state_in_14 ? 8'hb1 : _GEN_14031; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14033 = 8'hd1 == io_state_in_14 ? 8'hba : _GEN_14032; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14034 = 8'hd2 == io_state_in_14 ? 8'ha7 : _GEN_14033; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14035 = 8'hd3 == io_state_in_14 ? 8'hac : _GEN_14034; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14036 = 8'hd4 == io_state_in_14 ? 8'h9d : _GEN_14035; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14037 = 8'hd5 == io_state_in_14 ? 8'h96 : _GEN_14036; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14038 = 8'hd6 == io_state_in_14 ? 8'h8b : _GEN_14037; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14039 = 8'hd7 == io_state_in_14 ? 8'h80 : _GEN_14038; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14040 = 8'hd8 == io_state_in_14 ? 8'he9 : _GEN_14039; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14041 = 8'hd9 == io_state_in_14 ? 8'he2 : _GEN_14040; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14042 = 8'hda == io_state_in_14 ? 8'hff : _GEN_14041; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14043 = 8'hdb == io_state_in_14 ? 8'hf4 : _GEN_14042; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14044 = 8'hdc == io_state_in_14 ? 8'hc5 : _GEN_14043; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14045 = 8'hdd == io_state_in_14 ? 8'hce : _GEN_14044; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14046 = 8'hde == io_state_in_14 ? 8'hd3 : _GEN_14045; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14047 = 8'hdf == io_state_in_14 ? 8'hd8 : _GEN_14046; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14048 = 8'he0 == io_state_in_14 ? 8'h7a : _GEN_14047; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14049 = 8'he1 == io_state_in_14 ? 8'h71 : _GEN_14048; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14050 = 8'he2 == io_state_in_14 ? 8'h6c : _GEN_14049; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14051 = 8'he3 == io_state_in_14 ? 8'h67 : _GEN_14050; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14052 = 8'he4 == io_state_in_14 ? 8'h56 : _GEN_14051; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14053 = 8'he5 == io_state_in_14 ? 8'h5d : _GEN_14052; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14054 = 8'he6 == io_state_in_14 ? 8'h40 : _GEN_14053; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14055 = 8'he7 == io_state_in_14 ? 8'h4b : _GEN_14054; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14056 = 8'he8 == io_state_in_14 ? 8'h22 : _GEN_14055; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14057 = 8'he9 == io_state_in_14 ? 8'h29 : _GEN_14056; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14058 = 8'hea == io_state_in_14 ? 8'h34 : _GEN_14057; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14059 = 8'heb == io_state_in_14 ? 8'h3f : _GEN_14058; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14060 = 8'hec == io_state_in_14 ? 8'he : _GEN_14059; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14061 = 8'hed == io_state_in_14 ? 8'h5 : _GEN_14060; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14062 = 8'hee == io_state_in_14 ? 8'h18 : _GEN_14061; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14063 = 8'hef == io_state_in_14 ? 8'h13 : _GEN_14062; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14064 = 8'hf0 == io_state_in_14 ? 8'hca : _GEN_14063; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14065 = 8'hf1 == io_state_in_14 ? 8'hc1 : _GEN_14064; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14066 = 8'hf2 == io_state_in_14 ? 8'hdc : _GEN_14065; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14067 = 8'hf3 == io_state_in_14 ? 8'hd7 : _GEN_14066; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14068 = 8'hf4 == io_state_in_14 ? 8'he6 : _GEN_14067; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14069 = 8'hf5 == io_state_in_14 ? 8'hed : _GEN_14068; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14070 = 8'hf6 == io_state_in_14 ? 8'hf0 : _GEN_14069; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14071 = 8'hf7 == io_state_in_14 ? 8'hfb : _GEN_14070; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14072 = 8'hf8 == io_state_in_14 ? 8'h92 : _GEN_14071; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14073 = 8'hf9 == io_state_in_14 ? 8'h99 : _GEN_14072; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14074 = 8'hfa == io_state_in_14 ? 8'h84 : _GEN_14073; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14075 = 8'hfb == io_state_in_14 ? 8'h8f : _GEN_14074; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14076 = 8'hfc == io_state_in_14 ? 8'hbe : _GEN_14075; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14077 = 8'hfd == io_state_in_14 ? 8'hb5 : _GEN_14076; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14078 = 8'hfe == io_state_in_14 ? 8'ha8 : _GEN_14077; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _GEN_14079 = 8'hff == io_state_in_14 ? 8'ha3 : _GEN_14078; // @[InvMixColumns.scala 142:{68,68}]
  wire [7:0] _tmp_state_13_T_1 = _tmp_state_13_T ^ _GEN_14079; // @[InvMixColumns.scala 142:68]
  wire [7:0] _GEN_14081 = 8'h1 == io_state_in_15 ? 8'hd : 8'h0; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14082 = 8'h2 == io_state_in_15 ? 8'h1a : _GEN_14081; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14083 = 8'h3 == io_state_in_15 ? 8'h17 : _GEN_14082; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14084 = 8'h4 == io_state_in_15 ? 8'h34 : _GEN_14083; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14085 = 8'h5 == io_state_in_15 ? 8'h39 : _GEN_14084; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14086 = 8'h6 == io_state_in_15 ? 8'h2e : _GEN_14085; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14087 = 8'h7 == io_state_in_15 ? 8'h23 : _GEN_14086; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14088 = 8'h8 == io_state_in_15 ? 8'h68 : _GEN_14087; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14089 = 8'h9 == io_state_in_15 ? 8'h65 : _GEN_14088; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14090 = 8'ha == io_state_in_15 ? 8'h72 : _GEN_14089; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14091 = 8'hb == io_state_in_15 ? 8'h7f : _GEN_14090; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14092 = 8'hc == io_state_in_15 ? 8'h5c : _GEN_14091; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14093 = 8'hd == io_state_in_15 ? 8'h51 : _GEN_14092; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14094 = 8'he == io_state_in_15 ? 8'h46 : _GEN_14093; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14095 = 8'hf == io_state_in_15 ? 8'h4b : _GEN_14094; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14096 = 8'h10 == io_state_in_15 ? 8'hd0 : _GEN_14095; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14097 = 8'h11 == io_state_in_15 ? 8'hdd : _GEN_14096; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14098 = 8'h12 == io_state_in_15 ? 8'hca : _GEN_14097; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14099 = 8'h13 == io_state_in_15 ? 8'hc7 : _GEN_14098; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14100 = 8'h14 == io_state_in_15 ? 8'he4 : _GEN_14099; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14101 = 8'h15 == io_state_in_15 ? 8'he9 : _GEN_14100; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14102 = 8'h16 == io_state_in_15 ? 8'hfe : _GEN_14101; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14103 = 8'h17 == io_state_in_15 ? 8'hf3 : _GEN_14102; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14104 = 8'h18 == io_state_in_15 ? 8'hb8 : _GEN_14103; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14105 = 8'h19 == io_state_in_15 ? 8'hb5 : _GEN_14104; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14106 = 8'h1a == io_state_in_15 ? 8'ha2 : _GEN_14105; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14107 = 8'h1b == io_state_in_15 ? 8'haf : _GEN_14106; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14108 = 8'h1c == io_state_in_15 ? 8'h8c : _GEN_14107; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14109 = 8'h1d == io_state_in_15 ? 8'h81 : _GEN_14108; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14110 = 8'h1e == io_state_in_15 ? 8'h96 : _GEN_14109; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14111 = 8'h1f == io_state_in_15 ? 8'h9b : _GEN_14110; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14112 = 8'h20 == io_state_in_15 ? 8'hbb : _GEN_14111; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14113 = 8'h21 == io_state_in_15 ? 8'hb6 : _GEN_14112; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14114 = 8'h22 == io_state_in_15 ? 8'ha1 : _GEN_14113; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14115 = 8'h23 == io_state_in_15 ? 8'hac : _GEN_14114; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14116 = 8'h24 == io_state_in_15 ? 8'h8f : _GEN_14115; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14117 = 8'h25 == io_state_in_15 ? 8'h82 : _GEN_14116; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14118 = 8'h26 == io_state_in_15 ? 8'h95 : _GEN_14117; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14119 = 8'h27 == io_state_in_15 ? 8'h98 : _GEN_14118; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14120 = 8'h28 == io_state_in_15 ? 8'hd3 : _GEN_14119; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14121 = 8'h29 == io_state_in_15 ? 8'hde : _GEN_14120; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14122 = 8'h2a == io_state_in_15 ? 8'hc9 : _GEN_14121; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14123 = 8'h2b == io_state_in_15 ? 8'hc4 : _GEN_14122; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14124 = 8'h2c == io_state_in_15 ? 8'he7 : _GEN_14123; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14125 = 8'h2d == io_state_in_15 ? 8'hea : _GEN_14124; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14126 = 8'h2e == io_state_in_15 ? 8'hfd : _GEN_14125; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14127 = 8'h2f == io_state_in_15 ? 8'hf0 : _GEN_14126; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14128 = 8'h30 == io_state_in_15 ? 8'h6b : _GEN_14127; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14129 = 8'h31 == io_state_in_15 ? 8'h66 : _GEN_14128; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14130 = 8'h32 == io_state_in_15 ? 8'h71 : _GEN_14129; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14131 = 8'h33 == io_state_in_15 ? 8'h7c : _GEN_14130; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14132 = 8'h34 == io_state_in_15 ? 8'h5f : _GEN_14131; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14133 = 8'h35 == io_state_in_15 ? 8'h52 : _GEN_14132; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14134 = 8'h36 == io_state_in_15 ? 8'h45 : _GEN_14133; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14135 = 8'h37 == io_state_in_15 ? 8'h48 : _GEN_14134; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14136 = 8'h38 == io_state_in_15 ? 8'h3 : _GEN_14135; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14137 = 8'h39 == io_state_in_15 ? 8'he : _GEN_14136; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14138 = 8'h3a == io_state_in_15 ? 8'h19 : _GEN_14137; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14139 = 8'h3b == io_state_in_15 ? 8'h14 : _GEN_14138; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14140 = 8'h3c == io_state_in_15 ? 8'h37 : _GEN_14139; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14141 = 8'h3d == io_state_in_15 ? 8'h3a : _GEN_14140; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14142 = 8'h3e == io_state_in_15 ? 8'h2d : _GEN_14141; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14143 = 8'h3f == io_state_in_15 ? 8'h20 : _GEN_14142; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14144 = 8'h40 == io_state_in_15 ? 8'h6d : _GEN_14143; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14145 = 8'h41 == io_state_in_15 ? 8'h60 : _GEN_14144; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14146 = 8'h42 == io_state_in_15 ? 8'h77 : _GEN_14145; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14147 = 8'h43 == io_state_in_15 ? 8'h7a : _GEN_14146; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14148 = 8'h44 == io_state_in_15 ? 8'h59 : _GEN_14147; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14149 = 8'h45 == io_state_in_15 ? 8'h54 : _GEN_14148; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14150 = 8'h46 == io_state_in_15 ? 8'h43 : _GEN_14149; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14151 = 8'h47 == io_state_in_15 ? 8'h4e : _GEN_14150; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14152 = 8'h48 == io_state_in_15 ? 8'h5 : _GEN_14151; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14153 = 8'h49 == io_state_in_15 ? 8'h8 : _GEN_14152; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14154 = 8'h4a == io_state_in_15 ? 8'h1f : _GEN_14153; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14155 = 8'h4b == io_state_in_15 ? 8'h12 : _GEN_14154; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14156 = 8'h4c == io_state_in_15 ? 8'h31 : _GEN_14155; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14157 = 8'h4d == io_state_in_15 ? 8'h3c : _GEN_14156; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14158 = 8'h4e == io_state_in_15 ? 8'h2b : _GEN_14157; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14159 = 8'h4f == io_state_in_15 ? 8'h26 : _GEN_14158; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14160 = 8'h50 == io_state_in_15 ? 8'hbd : _GEN_14159; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14161 = 8'h51 == io_state_in_15 ? 8'hb0 : _GEN_14160; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14162 = 8'h52 == io_state_in_15 ? 8'ha7 : _GEN_14161; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14163 = 8'h53 == io_state_in_15 ? 8'haa : _GEN_14162; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14164 = 8'h54 == io_state_in_15 ? 8'h89 : _GEN_14163; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14165 = 8'h55 == io_state_in_15 ? 8'h84 : _GEN_14164; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14166 = 8'h56 == io_state_in_15 ? 8'h93 : _GEN_14165; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14167 = 8'h57 == io_state_in_15 ? 8'h9e : _GEN_14166; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14168 = 8'h58 == io_state_in_15 ? 8'hd5 : _GEN_14167; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14169 = 8'h59 == io_state_in_15 ? 8'hd8 : _GEN_14168; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14170 = 8'h5a == io_state_in_15 ? 8'hcf : _GEN_14169; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14171 = 8'h5b == io_state_in_15 ? 8'hc2 : _GEN_14170; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14172 = 8'h5c == io_state_in_15 ? 8'he1 : _GEN_14171; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14173 = 8'h5d == io_state_in_15 ? 8'hec : _GEN_14172; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14174 = 8'h5e == io_state_in_15 ? 8'hfb : _GEN_14173; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14175 = 8'h5f == io_state_in_15 ? 8'hf6 : _GEN_14174; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14176 = 8'h60 == io_state_in_15 ? 8'hd6 : _GEN_14175; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14177 = 8'h61 == io_state_in_15 ? 8'hdb : _GEN_14176; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14178 = 8'h62 == io_state_in_15 ? 8'hcc : _GEN_14177; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14179 = 8'h63 == io_state_in_15 ? 8'hc1 : _GEN_14178; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14180 = 8'h64 == io_state_in_15 ? 8'he2 : _GEN_14179; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14181 = 8'h65 == io_state_in_15 ? 8'hef : _GEN_14180; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14182 = 8'h66 == io_state_in_15 ? 8'hf8 : _GEN_14181; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14183 = 8'h67 == io_state_in_15 ? 8'hf5 : _GEN_14182; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14184 = 8'h68 == io_state_in_15 ? 8'hbe : _GEN_14183; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14185 = 8'h69 == io_state_in_15 ? 8'hb3 : _GEN_14184; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14186 = 8'h6a == io_state_in_15 ? 8'ha4 : _GEN_14185; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14187 = 8'h6b == io_state_in_15 ? 8'ha9 : _GEN_14186; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14188 = 8'h6c == io_state_in_15 ? 8'h8a : _GEN_14187; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14189 = 8'h6d == io_state_in_15 ? 8'h87 : _GEN_14188; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14190 = 8'h6e == io_state_in_15 ? 8'h90 : _GEN_14189; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14191 = 8'h6f == io_state_in_15 ? 8'h9d : _GEN_14190; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14192 = 8'h70 == io_state_in_15 ? 8'h6 : _GEN_14191; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14193 = 8'h71 == io_state_in_15 ? 8'hb : _GEN_14192; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14194 = 8'h72 == io_state_in_15 ? 8'h1c : _GEN_14193; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14195 = 8'h73 == io_state_in_15 ? 8'h11 : _GEN_14194; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14196 = 8'h74 == io_state_in_15 ? 8'h32 : _GEN_14195; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14197 = 8'h75 == io_state_in_15 ? 8'h3f : _GEN_14196; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14198 = 8'h76 == io_state_in_15 ? 8'h28 : _GEN_14197; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14199 = 8'h77 == io_state_in_15 ? 8'h25 : _GEN_14198; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14200 = 8'h78 == io_state_in_15 ? 8'h6e : _GEN_14199; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14201 = 8'h79 == io_state_in_15 ? 8'h63 : _GEN_14200; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14202 = 8'h7a == io_state_in_15 ? 8'h74 : _GEN_14201; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14203 = 8'h7b == io_state_in_15 ? 8'h79 : _GEN_14202; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14204 = 8'h7c == io_state_in_15 ? 8'h5a : _GEN_14203; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14205 = 8'h7d == io_state_in_15 ? 8'h57 : _GEN_14204; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14206 = 8'h7e == io_state_in_15 ? 8'h40 : _GEN_14205; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14207 = 8'h7f == io_state_in_15 ? 8'h4d : _GEN_14206; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14208 = 8'h80 == io_state_in_15 ? 8'hda : _GEN_14207; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14209 = 8'h81 == io_state_in_15 ? 8'hd7 : _GEN_14208; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14210 = 8'h82 == io_state_in_15 ? 8'hc0 : _GEN_14209; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14211 = 8'h83 == io_state_in_15 ? 8'hcd : _GEN_14210; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14212 = 8'h84 == io_state_in_15 ? 8'hee : _GEN_14211; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14213 = 8'h85 == io_state_in_15 ? 8'he3 : _GEN_14212; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14214 = 8'h86 == io_state_in_15 ? 8'hf4 : _GEN_14213; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14215 = 8'h87 == io_state_in_15 ? 8'hf9 : _GEN_14214; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14216 = 8'h88 == io_state_in_15 ? 8'hb2 : _GEN_14215; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14217 = 8'h89 == io_state_in_15 ? 8'hbf : _GEN_14216; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14218 = 8'h8a == io_state_in_15 ? 8'ha8 : _GEN_14217; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14219 = 8'h8b == io_state_in_15 ? 8'ha5 : _GEN_14218; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14220 = 8'h8c == io_state_in_15 ? 8'h86 : _GEN_14219; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14221 = 8'h8d == io_state_in_15 ? 8'h8b : _GEN_14220; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14222 = 8'h8e == io_state_in_15 ? 8'h9c : _GEN_14221; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14223 = 8'h8f == io_state_in_15 ? 8'h91 : _GEN_14222; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14224 = 8'h90 == io_state_in_15 ? 8'ha : _GEN_14223; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14225 = 8'h91 == io_state_in_15 ? 8'h7 : _GEN_14224; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14226 = 8'h92 == io_state_in_15 ? 8'h10 : _GEN_14225; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14227 = 8'h93 == io_state_in_15 ? 8'h1d : _GEN_14226; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14228 = 8'h94 == io_state_in_15 ? 8'h3e : _GEN_14227; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14229 = 8'h95 == io_state_in_15 ? 8'h33 : _GEN_14228; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14230 = 8'h96 == io_state_in_15 ? 8'h24 : _GEN_14229; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14231 = 8'h97 == io_state_in_15 ? 8'h29 : _GEN_14230; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14232 = 8'h98 == io_state_in_15 ? 8'h62 : _GEN_14231; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14233 = 8'h99 == io_state_in_15 ? 8'h6f : _GEN_14232; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14234 = 8'h9a == io_state_in_15 ? 8'h78 : _GEN_14233; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14235 = 8'h9b == io_state_in_15 ? 8'h75 : _GEN_14234; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14236 = 8'h9c == io_state_in_15 ? 8'h56 : _GEN_14235; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14237 = 8'h9d == io_state_in_15 ? 8'h5b : _GEN_14236; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14238 = 8'h9e == io_state_in_15 ? 8'h4c : _GEN_14237; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14239 = 8'h9f == io_state_in_15 ? 8'h41 : _GEN_14238; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14240 = 8'ha0 == io_state_in_15 ? 8'h61 : _GEN_14239; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14241 = 8'ha1 == io_state_in_15 ? 8'h6c : _GEN_14240; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14242 = 8'ha2 == io_state_in_15 ? 8'h7b : _GEN_14241; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14243 = 8'ha3 == io_state_in_15 ? 8'h76 : _GEN_14242; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14244 = 8'ha4 == io_state_in_15 ? 8'h55 : _GEN_14243; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14245 = 8'ha5 == io_state_in_15 ? 8'h58 : _GEN_14244; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14246 = 8'ha6 == io_state_in_15 ? 8'h4f : _GEN_14245; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14247 = 8'ha7 == io_state_in_15 ? 8'h42 : _GEN_14246; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14248 = 8'ha8 == io_state_in_15 ? 8'h9 : _GEN_14247; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14249 = 8'ha9 == io_state_in_15 ? 8'h4 : _GEN_14248; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14250 = 8'haa == io_state_in_15 ? 8'h13 : _GEN_14249; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14251 = 8'hab == io_state_in_15 ? 8'h1e : _GEN_14250; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14252 = 8'hac == io_state_in_15 ? 8'h3d : _GEN_14251; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14253 = 8'had == io_state_in_15 ? 8'h30 : _GEN_14252; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14254 = 8'hae == io_state_in_15 ? 8'h27 : _GEN_14253; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14255 = 8'haf == io_state_in_15 ? 8'h2a : _GEN_14254; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14256 = 8'hb0 == io_state_in_15 ? 8'hb1 : _GEN_14255; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14257 = 8'hb1 == io_state_in_15 ? 8'hbc : _GEN_14256; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14258 = 8'hb2 == io_state_in_15 ? 8'hab : _GEN_14257; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14259 = 8'hb3 == io_state_in_15 ? 8'ha6 : _GEN_14258; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14260 = 8'hb4 == io_state_in_15 ? 8'h85 : _GEN_14259; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14261 = 8'hb5 == io_state_in_15 ? 8'h88 : _GEN_14260; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14262 = 8'hb6 == io_state_in_15 ? 8'h9f : _GEN_14261; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14263 = 8'hb7 == io_state_in_15 ? 8'h92 : _GEN_14262; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14264 = 8'hb8 == io_state_in_15 ? 8'hd9 : _GEN_14263; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14265 = 8'hb9 == io_state_in_15 ? 8'hd4 : _GEN_14264; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14266 = 8'hba == io_state_in_15 ? 8'hc3 : _GEN_14265; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14267 = 8'hbb == io_state_in_15 ? 8'hce : _GEN_14266; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14268 = 8'hbc == io_state_in_15 ? 8'hed : _GEN_14267; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14269 = 8'hbd == io_state_in_15 ? 8'he0 : _GEN_14268; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14270 = 8'hbe == io_state_in_15 ? 8'hf7 : _GEN_14269; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14271 = 8'hbf == io_state_in_15 ? 8'hfa : _GEN_14270; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14272 = 8'hc0 == io_state_in_15 ? 8'hb7 : _GEN_14271; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14273 = 8'hc1 == io_state_in_15 ? 8'hba : _GEN_14272; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14274 = 8'hc2 == io_state_in_15 ? 8'had : _GEN_14273; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14275 = 8'hc3 == io_state_in_15 ? 8'ha0 : _GEN_14274; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14276 = 8'hc4 == io_state_in_15 ? 8'h83 : _GEN_14275; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14277 = 8'hc5 == io_state_in_15 ? 8'h8e : _GEN_14276; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14278 = 8'hc6 == io_state_in_15 ? 8'h99 : _GEN_14277; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14279 = 8'hc7 == io_state_in_15 ? 8'h94 : _GEN_14278; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14280 = 8'hc8 == io_state_in_15 ? 8'hdf : _GEN_14279; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14281 = 8'hc9 == io_state_in_15 ? 8'hd2 : _GEN_14280; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14282 = 8'hca == io_state_in_15 ? 8'hc5 : _GEN_14281; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14283 = 8'hcb == io_state_in_15 ? 8'hc8 : _GEN_14282; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14284 = 8'hcc == io_state_in_15 ? 8'heb : _GEN_14283; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14285 = 8'hcd == io_state_in_15 ? 8'he6 : _GEN_14284; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14286 = 8'hce == io_state_in_15 ? 8'hf1 : _GEN_14285; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14287 = 8'hcf == io_state_in_15 ? 8'hfc : _GEN_14286; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14288 = 8'hd0 == io_state_in_15 ? 8'h67 : _GEN_14287; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14289 = 8'hd1 == io_state_in_15 ? 8'h6a : _GEN_14288; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14290 = 8'hd2 == io_state_in_15 ? 8'h7d : _GEN_14289; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14291 = 8'hd3 == io_state_in_15 ? 8'h70 : _GEN_14290; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14292 = 8'hd4 == io_state_in_15 ? 8'h53 : _GEN_14291; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14293 = 8'hd5 == io_state_in_15 ? 8'h5e : _GEN_14292; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14294 = 8'hd6 == io_state_in_15 ? 8'h49 : _GEN_14293; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14295 = 8'hd7 == io_state_in_15 ? 8'h44 : _GEN_14294; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14296 = 8'hd8 == io_state_in_15 ? 8'hf : _GEN_14295; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14297 = 8'hd9 == io_state_in_15 ? 8'h2 : _GEN_14296; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14298 = 8'hda == io_state_in_15 ? 8'h15 : _GEN_14297; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14299 = 8'hdb == io_state_in_15 ? 8'h18 : _GEN_14298; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14300 = 8'hdc == io_state_in_15 ? 8'h3b : _GEN_14299; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14301 = 8'hdd == io_state_in_15 ? 8'h36 : _GEN_14300; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14302 = 8'hde == io_state_in_15 ? 8'h21 : _GEN_14301; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14303 = 8'hdf == io_state_in_15 ? 8'h2c : _GEN_14302; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14304 = 8'he0 == io_state_in_15 ? 8'hc : _GEN_14303; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14305 = 8'he1 == io_state_in_15 ? 8'h1 : _GEN_14304; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14306 = 8'he2 == io_state_in_15 ? 8'h16 : _GEN_14305; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14307 = 8'he3 == io_state_in_15 ? 8'h1b : _GEN_14306; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14308 = 8'he4 == io_state_in_15 ? 8'h38 : _GEN_14307; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14309 = 8'he5 == io_state_in_15 ? 8'h35 : _GEN_14308; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14310 = 8'he6 == io_state_in_15 ? 8'h22 : _GEN_14309; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14311 = 8'he7 == io_state_in_15 ? 8'h2f : _GEN_14310; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14312 = 8'he8 == io_state_in_15 ? 8'h64 : _GEN_14311; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14313 = 8'he9 == io_state_in_15 ? 8'h69 : _GEN_14312; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14314 = 8'hea == io_state_in_15 ? 8'h7e : _GEN_14313; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14315 = 8'heb == io_state_in_15 ? 8'h73 : _GEN_14314; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14316 = 8'hec == io_state_in_15 ? 8'h50 : _GEN_14315; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14317 = 8'hed == io_state_in_15 ? 8'h5d : _GEN_14316; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14318 = 8'hee == io_state_in_15 ? 8'h4a : _GEN_14317; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14319 = 8'hef == io_state_in_15 ? 8'h47 : _GEN_14318; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14320 = 8'hf0 == io_state_in_15 ? 8'hdc : _GEN_14319; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14321 = 8'hf1 == io_state_in_15 ? 8'hd1 : _GEN_14320; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14322 = 8'hf2 == io_state_in_15 ? 8'hc6 : _GEN_14321; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14323 = 8'hf3 == io_state_in_15 ? 8'hcb : _GEN_14322; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14324 = 8'hf4 == io_state_in_15 ? 8'he8 : _GEN_14323; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14325 = 8'hf5 == io_state_in_15 ? 8'he5 : _GEN_14324; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14326 = 8'hf6 == io_state_in_15 ? 8'hf2 : _GEN_14325; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14327 = 8'hf7 == io_state_in_15 ? 8'hff : _GEN_14326; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14328 = 8'hf8 == io_state_in_15 ? 8'hb4 : _GEN_14327; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14329 = 8'hf9 == io_state_in_15 ? 8'hb9 : _GEN_14328; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14330 = 8'hfa == io_state_in_15 ? 8'hae : _GEN_14329; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14331 = 8'hfb == io_state_in_15 ? 8'ha3 : _GEN_14330; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14332 = 8'hfc == io_state_in_15 ? 8'h80 : _GEN_14331; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14333 = 8'hfd == io_state_in_15 ? 8'h8d : _GEN_14332; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14334 = 8'hfe == io_state_in_15 ? 8'h9a : _GEN_14333; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14335 = 8'hff == io_state_in_15 ? 8'h97 : _GEN_14334; // @[InvMixColumns.scala 142:{93,93}]
  wire [7:0] _GEN_14337 = 8'h1 == io_state_in_12 ? 8'hd : 8'h0; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14338 = 8'h2 == io_state_in_12 ? 8'h1a : _GEN_14337; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14339 = 8'h3 == io_state_in_12 ? 8'h17 : _GEN_14338; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14340 = 8'h4 == io_state_in_12 ? 8'h34 : _GEN_14339; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14341 = 8'h5 == io_state_in_12 ? 8'h39 : _GEN_14340; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14342 = 8'h6 == io_state_in_12 ? 8'h2e : _GEN_14341; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14343 = 8'h7 == io_state_in_12 ? 8'h23 : _GEN_14342; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14344 = 8'h8 == io_state_in_12 ? 8'h68 : _GEN_14343; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14345 = 8'h9 == io_state_in_12 ? 8'h65 : _GEN_14344; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14346 = 8'ha == io_state_in_12 ? 8'h72 : _GEN_14345; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14347 = 8'hb == io_state_in_12 ? 8'h7f : _GEN_14346; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14348 = 8'hc == io_state_in_12 ? 8'h5c : _GEN_14347; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14349 = 8'hd == io_state_in_12 ? 8'h51 : _GEN_14348; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14350 = 8'he == io_state_in_12 ? 8'h46 : _GEN_14349; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14351 = 8'hf == io_state_in_12 ? 8'h4b : _GEN_14350; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14352 = 8'h10 == io_state_in_12 ? 8'hd0 : _GEN_14351; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14353 = 8'h11 == io_state_in_12 ? 8'hdd : _GEN_14352; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14354 = 8'h12 == io_state_in_12 ? 8'hca : _GEN_14353; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14355 = 8'h13 == io_state_in_12 ? 8'hc7 : _GEN_14354; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14356 = 8'h14 == io_state_in_12 ? 8'he4 : _GEN_14355; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14357 = 8'h15 == io_state_in_12 ? 8'he9 : _GEN_14356; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14358 = 8'h16 == io_state_in_12 ? 8'hfe : _GEN_14357; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14359 = 8'h17 == io_state_in_12 ? 8'hf3 : _GEN_14358; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14360 = 8'h18 == io_state_in_12 ? 8'hb8 : _GEN_14359; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14361 = 8'h19 == io_state_in_12 ? 8'hb5 : _GEN_14360; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14362 = 8'h1a == io_state_in_12 ? 8'ha2 : _GEN_14361; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14363 = 8'h1b == io_state_in_12 ? 8'haf : _GEN_14362; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14364 = 8'h1c == io_state_in_12 ? 8'h8c : _GEN_14363; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14365 = 8'h1d == io_state_in_12 ? 8'h81 : _GEN_14364; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14366 = 8'h1e == io_state_in_12 ? 8'h96 : _GEN_14365; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14367 = 8'h1f == io_state_in_12 ? 8'h9b : _GEN_14366; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14368 = 8'h20 == io_state_in_12 ? 8'hbb : _GEN_14367; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14369 = 8'h21 == io_state_in_12 ? 8'hb6 : _GEN_14368; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14370 = 8'h22 == io_state_in_12 ? 8'ha1 : _GEN_14369; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14371 = 8'h23 == io_state_in_12 ? 8'hac : _GEN_14370; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14372 = 8'h24 == io_state_in_12 ? 8'h8f : _GEN_14371; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14373 = 8'h25 == io_state_in_12 ? 8'h82 : _GEN_14372; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14374 = 8'h26 == io_state_in_12 ? 8'h95 : _GEN_14373; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14375 = 8'h27 == io_state_in_12 ? 8'h98 : _GEN_14374; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14376 = 8'h28 == io_state_in_12 ? 8'hd3 : _GEN_14375; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14377 = 8'h29 == io_state_in_12 ? 8'hde : _GEN_14376; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14378 = 8'h2a == io_state_in_12 ? 8'hc9 : _GEN_14377; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14379 = 8'h2b == io_state_in_12 ? 8'hc4 : _GEN_14378; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14380 = 8'h2c == io_state_in_12 ? 8'he7 : _GEN_14379; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14381 = 8'h2d == io_state_in_12 ? 8'hea : _GEN_14380; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14382 = 8'h2e == io_state_in_12 ? 8'hfd : _GEN_14381; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14383 = 8'h2f == io_state_in_12 ? 8'hf0 : _GEN_14382; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14384 = 8'h30 == io_state_in_12 ? 8'h6b : _GEN_14383; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14385 = 8'h31 == io_state_in_12 ? 8'h66 : _GEN_14384; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14386 = 8'h32 == io_state_in_12 ? 8'h71 : _GEN_14385; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14387 = 8'h33 == io_state_in_12 ? 8'h7c : _GEN_14386; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14388 = 8'h34 == io_state_in_12 ? 8'h5f : _GEN_14387; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14389 = 8'h35 == io_state_in_12 ? 8'h52 : _GEN_14388; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14390 = 8'h36 == io_state_in_12 ? 8'h45 : _GEN_14389; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14391 = 8'h37 == io_state_in_12 ? 8'h48 : _GEN_14390; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14392 = 8'h38 == io_state_in_12 ? 8'h3 : _GEN_14391; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14393 = 8'h39 == io_state_in_12 ? 8'he : _GEN_14392; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14394 = 8'h3a == io_state_in_12 ? 8'h19 : _GEN_14393; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14395 = 8'h3b == io_state_in_12 ? 8'h14 : _GEN_14394; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14396 = 8'h3c == io_state_in_12 ? 8'h37 : _GEN_14395; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14397 = 8'h3d == io_state_in_12 ? 8'h3a : _GEN_14396; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14398 = 8'h3e == io_state_in_12 ? 8'h2d : _GEN_14397; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14399 = 8'h3f == io_state_in_12 ? 8'h20 : _GEN_14398; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14400 = 8'h40 == io_state_in_12 ? 8'h6d : _GEN_14399; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14401 = 8'h41 == io_state_in_12 ? 8'h60 : _GEN_14400; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14402 = 8'h42 == io_state_in_12 ? 8'h77 : _GEN_14401; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14403 = 8'h43 == io_state_in_12 ? 8'h7a : _GEN_14402; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14404 = 8'h44 == io_state_in_12 ? 8'h59 : _GEN_14403; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14405 = 8'h45 == io_state_in_12 ? 8'h54 : _GEN_14404; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14406 = 8'h46 == io_state_in_12 ? 8'h43 : _GEN_14405; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14407 = 8'h47 == io_state_in_12 ? 8'h4e : _GEN_14406; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14408 = 8'h48 == io_state_in_12 ? 8'h5 : _GEN_14407; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14409 = 8'h49 == io_state_in_12 ? 8'h8 : _GEN_14408; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14410 = 8'h4a == io_state_in_12 ? 8'h1f : _GEN_14409; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14411 = 8'h4b == io_state_in_12 ? 8'h12 : _GEN_14410; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14412 = 8'h4c == io_state_in_12 ? 8'h31 : _GEN_14411; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14413 = 8'h4d == io_state_in_12 ? 8'h3c : _GEN_14412; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14414 = 8'h4e == io_state_in_12 ? 8'h2b : _GEN_14413; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14415 = 8'h4f == io_state_in_12 ? 8'h26 : _GEN_14414; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14416 = 8'h50 == io_state_in_12 ? 8'hbd : _GEN_14415; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14417 = 8'h51 == io_state_in_12 ? 8'hb0 : _GEN_14416; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14418 = 8'h52 == io_state_in_12 ? 8'ha7 : _GEN_14417; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14419 = 8'h53 == io_state_in_12 ? 8'haa : _GEN_14418; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14420 = 8'h54 == io_state_in_12 ? 8'h89 : _GEN_14419; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14421 = 8'h55 == io_state_in_12 ? 8'h84 : _GEN_14420; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14422 = 8'h56 == io_state_in_12 ? 8'h93 : _GEN_14421; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14423 = 8'h57 == io_state_in_12 ? 8'h9e : _GEN_14422; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14424 = 8'h58 == io_state_in_12 ? 8'hd5 : _GEN_14423; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14425 = 8'h59 == io_state_in_12 ? 8'hd8 : _GEN_14424; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14426 = 8'h5a == io_state_in_12 ? 8'hcf : _GEN_14425; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14427 = 8'h5b == io_state_in_12 ? 8'hc2 : _GEN_14426; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14428 = 8'h5c == io_state_in_12 ? 8'he1 : _GEN_14427; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14429 = 8'h5d == io_state_in_12 ? 8'hec : _GEN_14428; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14430 = 8'h5e == io_state_in_12 ? 8'hfb : _GEN_14429; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14431 = 8'h5f == io_state_in_12 ? 8'hf6 : _GEN_14430; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14432 = 8'h60 == io_state_in_12 ? 8'hd6 : _GEN_14431; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14433 = 8'h61 == io_state_in_12 ? 8'hdb : _GEN_14432; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14434 = 8'h62 == io_state_in_12 ? 8'hcc : _GEN_14433; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14435 = 8'h63 == io_state_in_12 ? 8'hc1 : _GEN_14434; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14436 = 8'h64 == io_state_in_12 ? 8'he2 : _GEN_14435; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14437 = 8'h65 == io_state_in_12 ? 8'hef : _GEN_14436; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14438 = 8'h66 == io_state_in_12 ? 8'hf8 : _GEN_14437; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14439 = 8'h67 == io_state_in_12 ? 8'hf5 : _GEN_14438; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14440 = 8'h68 == io_state_in_12 ? 8'hbe : _GEN_14439; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14441 = 8'h69 == io_state_in_12 ? 8'hb3 : _GEN_14440; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14442 = 8'h6a == io_state_in_12 ? 8'ha4 : _GEN_14441; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14443 = 8'h6b == io_state_in_12 ? 8'ha9 : _GEN_14442; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14444 = 8'h6c == io_state_in_12 ? 8'h8a : _GEN_14443; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14445 = 8'h6d == io_state_in_12 ? 8'h87 : _GEN_14444; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14446 = 8'h6e == io_state_in_12 ? 8'h90 : _GEN_14445; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14447 = 8'h6f == io_state_in_12 ? 8'h9d : _GEN_14446; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14448 = 8'h70 == io_state_in_12 ? 8'h6 : _GEN_14447; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14449 = 8'h71 == io_state_in_12 ? 8'hb : _GEN_14448; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14450 = 8'h72 == io_state_in_12 ? 8'h1c : _GEN_14449; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14451 = 8'h73 == io_state_in_12 ? 8'h11 : _GEN_14450; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14452 = 8'h74 == io_state_in_12 ? 8'h32 : _GEN_14451; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14453 = 8'h75 == io_state_in_12 ? 8'h3f : _GEN_14452; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14454 = 8'h76 == io_state_in_12 ? 8'h28 : _GEN_14453; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14455 = 8'h77 == io_state_in_12 ? 8'h25 : _GEN_14454; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14456 = 8'h78 == io_state_in_12 ? 8'h6e : _GEN_14455; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14457 = 8'h79 == io_state_in_12 ? 8'h63 : _GEN_14456; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14458 = 8'h7a == io_state_in_12 ? 8'h74 : _GEN_14457; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14459 = 8'h7b == io_state_in_12 ? 8'h79 : _GEN_14458; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14460 = 8'h7c == io_state_in_12 ? 8'h5a : _GEN_14459; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14461 = 8'h7d == io_state_in_12 ? 8'h57 : _GEN_14460; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14462 = 8'h7e == io_state_in_12 ? 8'h40 : _GEN_14461; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14463 = 8'h7f == io_state_in_12 ? 8'h4d : _GEN_14462; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14464 = 8'h80 == io_state_in_12 ? 8'hda : _GEN_14463; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14465 = 8'h81 == io_state_in_12 ? 8'hd7 : _GEN_14464; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14466 = 8'h82 == io_state_in_12 ? 8'hc0 : _GEN_14465; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14467 = 8'h83 == io_state_in_12 ? 8'hcd : _GEN_14466; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14468 = 8'h84 == io_state_in_12 ? 8'hee : _GEN_14467; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14469 = 8'h85 == io_state_in_12 ? 8'he3 : _GEN_14468; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14470 = 8'h86 == io_state_in_12 ? 8'hf4 : _GEN_14469; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14471 = 8'h87 == io_state_in_12 ? 8'hf9 : _GEN_14470; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14472 = 8'h88 == io_state_in_12 ? 8'hb2 : _GEN_14471; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14473 = 8'h89 == io_state_in_12 ? 8'hbf : _GEN_14472; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14474 = 8'h8a == io_state_in_12 ? 8'ha8 : _GEN_14473; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14475 = 8'h8b == io_state_in_12 ? 8'ha5 : _GEN_14474; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14476 = 8'h8c == io_state_in_12 ? 8'h86 : _GEN_14475; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14477 = 8'h8d == io_state_in_12 ? 8'h8b : _GEN_14476; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14478 = 8'h8e == io_state_in_12 ? 8'h9c : _GEN_14477; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14479 = 8'h8f == io_state_in_12 ? 8'h91 : _GEN_14478; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14480 = 8'h90 == io_state_in_12 ? 8'ha : _GEN_14479; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14481 = 8'h91 == io_state_in_12 ? 8'h7 : _GEN_14480; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14482 = 8'h92 == io_state_in_12 ? 8'h10 : _GEN_14481; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14483 = 8'h93 == io_state_in_12 ? 8'h1d : _GEN_14482; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14484 = 8'h94 == io_state_in_12 ? 8'h3e : _GEN_14483; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14485 = 8'h95 == io_state_in_12 ? 8'h33 : _GEN_14484; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14486 = 8'h96 == io_state_in_12 ? 8'h24 : _GEN_14485; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14487 = 8'h97 == io_state_in_12 ? 8'h29 : _GEN_14486; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14488 = 8'h98 == io_state_in_12 ? 8'h62 : _GEN_14487; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14489 = 8'h99 == io_state_in_12 ? 8'h6f : _GEN_14488; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14490 = 8'h9a == io_state_in_12 ? 8'h78 : _GEN_14489; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14491 = 8'h9b == io_state_in_12 ? 8'h75 : _GEN_14490; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14492 = 8'h9c == io_state_in_12 ? 8'h56 : _GEN_14491; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14493 = 8'h9d == io_state_in_12 ? 8'h5b : _GEN_14492; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14494 = 8'h9e == io_state_in_12 ? 8'h4c : _GEN_14493; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14495 = 8'h9f == io_state_in_12 ? 8'h41 : _GEN_14494; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14496 = 8'ha0 == io_state_in_12 ? 8'h61 : _GEN_14495; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14497 = 8'ha1 == io_state_in_12 ? 8'h6c : _GEN_14496; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14498 = 8'ha2 == io_state_in_12 ? 8'h7b : _GEN_14497; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14499 = 8'ha3 == io_state_in_12 ? 8'h76 : _GEN_14498; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14500 = 8'ha4 == io_state_in_12 ? 8'h55 : _GEN_14499; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14501 = 8'ha5 == io_state_in_12 ? 8'h58 : _GEN_14500; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14502 = 8'ha6 == io_state_in_12 ? 8'h4f : _GEN_14501; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14503 = 8'ha7 == io_state_in_12 ? 8'h42 : _GEN_14502; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14504 = 8'ha8 == io_state_in_12 ? 8'h9 : _GEN_14503; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14505 = 8'ha9 == io_state_in_12 ? 8'h4 : _GEN_14504; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14506 = 8'haa == io_state_in_12 ? 8'h13 : _GEN_14505; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14507 = 8'hab == io_state_in_12 ? 8'h1e : _GEN_14506; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14508 = 8'hac == io_state_in_12 ? 8'h3d : _GEN_14507; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14509 = 8'had == io_state_in_12 ? 8'h30 : _GEN_14508; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14510 = 8'hae == io_state_in_12 ? 8'h27 : _GEN_14509; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14511 = 8'haf == io_state_in_12 ? 8'h2a : _GEN_14510; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14512 = 8'hb0 == io_state_in_12 ? 8'hb1 : _GEN_14511; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14513 = 8'hb1 == io_state_in_12 ? 8'hbc : _GEN_14512; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14514 = 8'hb2 == io_state_in_12 ? 8'hab : _GEN_14513; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14515 = 8'hb3 == io_state_in_12 ? 8'ha6 : _GEN_14514; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14516 = 8'hb4 == io_state_in_12 ? 8'h85 : _GEN_14515; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14517 = 8'hb5 == io_state_in_12 ? 8'h88 : _GEN_14516; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14518 = 8'hb6 == io_state_in_12 ? 8'h9f : _GEN_14517; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14519 = 8'hb7 == io_state_in_12 ? 8'h92 : _GEN_14518; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14520 = 8'hb8 == io_state_in_12 ? 8'hd9 : _GEN_14519; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14521 = 8'hb9 == io_state_in_12 ? 8'hd4 : _GEN_14520; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14522 = 8'hba == io_state_in_12 ? 8'hc3 : _GEN_14521; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14523 = 8'hbb == io_state_in_12 ? 8'hce : _GEN_14522; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14524 = 8'hbc == io_state_in_12 ? 8'hed : _GEN_14523; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14525 = 8'hbd == io_state_in_12 ? 8'he0 : _GEN_14524; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14526 = 8'hbe == io_state_in_12 ? 8'hf7 : _GEN_14525; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14527 = 8'hbf == io_state_in_12 ? 8'hfa : _GEN_14526; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14528 = 8'hc0 == io_state_in_12 ? 8'hb7 : _GEN_14527; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14529 = 8'hc1 == io_state_in_12 ? 8'hba : _GEN_14528; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14530 = 8'hc2 == io_state_in_12 ? 8'had : _GEN_14529; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14531 = 8'hc3 == io_state_in_12 ? 8'ha0 : _GEN_14530; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14532 = 8'hc4 == io_state_in_12 ? 8'h83 : _GEN_14531; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14533 = 8'hc5 == io_state_in_12 ? 8'h8e : _GEN_14532; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14534 = 8'hc6 == io_state_in_12 ? 8'h99 : _GEN_14533; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14535 = 8'hc7 == io_state_in_12 ? 8'h94 : _GEN_14534; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14536 = 8'hc8 == io_state_in_12 ? 8'hdf : _GEN_14535; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14537 = 8'hc9 == io_state_in_12 ? 8'hd2 : _GEN_14536; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14538 = 8'hca == io_state_in_12 ? 8'hc5 : _GEN_14537; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14539 = 8'hcb == io_state_in_12 ? 8'hc8 : _GEN_14538; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14540 = 8'hcc == io_state_in_12 ? 8'heb : _GEN_14539; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14541 = 8'hcd == io_state_in_12 ? 8'he6 : _GEN_14540; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14542 = 8'hce == io_state_in_12 ? 8'hf1 : _GEN_14541; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14543 = 8'hcf == io_state_in_12 ? 8'hfc : _GEN_14542; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14544 = 8'hd0 == io_state_in_12 ? 8'h67 : _GEN_14543; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14545 = 8'hd1 == io_state_in_12 ? 8'h6a : _GEN_14544; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14546 = 8'hd2 == io_state_in_12 ? 8'h7d : _GEN_14545; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14547 = 8'hd3 == io_state_in_12 ? 8'h70 : _GEN_14546; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14548 = 8'hd4 == io_state_in_12 ? 8'h53 : _GEN_14547; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14549 = 8'hd5 == io_state_in_12 ? 8'h5e : _GEN_14548; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14550 = 8'hd6 == io_state_in_12 ? 8'h49 : _GEN_14549; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14551 = 8'hd7 == io_state_in_12 ? 8'h44 : _GEN_14550; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14552 = 8'hd8 == io_state_in_12 ? 8'hf : _GEN_14551; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14553 = 8'hd9 == io_state_in_12 ? 8'h2 : _GEN_14552; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14554 = 8'hda == io_state_in_12 ? 8'h15 : _GEN_14553; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14555 = 8'hdb == io_state_in_12 ? 8'h18 : _GEN_14554; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14556 = 8'hdc == io_state_in_12 ? 8'h3b : _GEN_14555; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14557 = 8'hdd == io_state_in_12 ? 8'h36 : _GEN_14556; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14558 = 8'hde == io_state_in_12 ? 8'h21 : _GEN_14557; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14559 = 8'hdf == io_state_in_12 ? 8'h2c : _GEN_14558; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14560 = 8'he0 == io_state_in_12 ? 8'hc : _GEN_14559; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14561 = 8'he1 == io_state_in_12 ? 8'h1 : _GEN_14560; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14562 = 8'he2 == io_state_in_12 ? 8'h16 : _GEN_14561; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14563 = 8'he3 == io_state_in_12 ? 8'h1b : _GEN_14562; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14564 = 8'he4 == io_state_in_12 ? 8'h38 : _GEN_14563; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14565 = 8'he5 == io_state_in_12 ? 8'h35 : _GEN_14564; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14566 = 8'he6 == io_state_in_12 ? 8'h22 : _GEN_14565; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14567 = 8'he7 == io_state_in_12 ? 8'h2f : _GEN_14566; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14568 = 8'he8 == io_state_in_12 ? 8'h64 : _GEN_14567; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14569 = 8'he9 == io_state_in_12 ? 8'h69 : _GEN_14568; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14570 = 8'hea == io_state_in_12 ? 8'h7e : _GEN_14569; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14571 = 8'heb == io_state_in_12 ? 8'h73 : _GEN_14570; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14572 = 8'hec == io_state_in_12 ? 8'h50 : _GEN_14571; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14573 = 8'hed == io_state_in_12 ? 8'h5d : _GEN_14572; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14574 = 8'hee == io_state_in_12 ? 8'h4a : _GEN_14573; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14575 = 8'hef == io_state_in_12 ? 8'h47 : _GEN_14574; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14576 = 8'hf0 == io_state_in_12 ? 8'hdc : _GEN_14575; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14577 = 8'hf1 == io_state_in_12 ? 8'hd1 : _GEN_14576; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14578 = 8'hf2 == io_state_in_12 ? 8'hc6 : _GEN_14577; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14579 = 8'hf3 == io_state_in_12 ? 8'hcb : _GEN_14578; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14580 = 8'hf4 == io_state_in_12 ? 8'he8 : _GEN_14579; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14581 = 8'hf5 == io_state_in_12 ? 8'he5 : _GEN_14580; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14582 = 8'hf6 == io_state_in_12 ? 8'hf2 : _GEN_14581; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14583 = 8'hf7 == io_state_in_12 ? 8'hff : _GEN_14582; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14584 = 8'hf8 == io_state_in_12 ? 8'hb4 : _GEN_14583; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14585 = 8'hf9 == io_state_in_12 ? 8'hb9 : _GEN_14584; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14586 = 8'hfa == io_state_in_12 ? 8'hae : _GEN_14585; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14587 = 8'hfb == io_state_in_12 ? 8'ha3 : _GEN_14586; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14588 = 8'hfc == io_state_in_12 ? 8'h80 : _GEN_14587; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14589 = 8'hfd == io_state_in_12 ? 8'h8d : _GEN_14588; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14590 = 8'hfe == io_state_in_12 ? 8'h9a : _GEN_14589; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14591 = 8'hff == io_state_in_12 ? 8'h97 : _GEN_14590; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14593 = 8'h1 == io_state_in_13 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14594 = 8'h2 == io_state_in_13 ? 8'h12 : _GEN_14593; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14595 = 8'h3 == io_state_in_13 ? 8'h1b : _GEN_14594; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14596 = 8'h4 == io_state_in_13 ? 8'h24 : _GEN_14595; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14597 = 8'h5 == io_state_in_13 ? 8'h2d : _GEN_14596; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14598 = 8'h6 == io_state_in_13 ? 8'h36 : _GEN_14597; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14599 = 8'h7 == io_state_in_13 ? 8'h3f : _GEN_14598; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14600 = 8'h8 == io_state_in_13 ? 8'h48 : _GEN_14599; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14601 = 8'h9 == io_state_in_13 ? 8'h41 : _GEN_14600; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14602 = 8'ha == io_state_in_13 ? 8'h5a : _GEN_14601; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14603 = 8'hb == io_state_in_13 ? 8'h53 : _GEN_14602; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14604 = 8'hc == io_state_in_13 ? 8'h6c : _GEN_14603; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14605 = 8'hd == io_state_in_13 ? 8'h65 : _GEN_14604; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14606 = 8'he == io_state_in_13 ? 8'h7e : _GEN_14605; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14607 = 8'hf == io_state_in_13 ? 8'h77 : _GEN_14606; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14608 = 8'h10 == io_state_in_13 ? 8'h90 : _GEN_14607; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14609 = 8'h11 == io_state_in_13 ? 8'h99 : _GEN_14608; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14610 = 8'h12 == io_state_in_13 ? 8'h82 : _GEN_14609; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14611 = 8'h13 == io_state_in_13 ? 8'h8b : _GEN_14610; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14612 = 8'h14 == io_state_in_13 ? 8'hb4 : _GEN_14611; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14613 = 8'h15 == io_state_in_13 ? 8'hbd : _GEN_14612; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14614 = 8'h16 == io_state_in_13 ? 8'ha6 : _GEN_14613; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14615 = 8'h17 == io_state_in_13 ? 8'haf : _GEN_14614; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14616 = 8'h18 == io_state_in_13 ? 8'hd8 : _GEN_14615; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14617 = 8'h19 == io_state_in_13 ? 8'hd1 : _GEN_14616; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14618 = 8'h1a == io_state_in_13 ? 8'hca : _GEN_14617; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14619 = 8'h1b == io_state_in_13 ? 8'hc3 : _GEN_14618; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14620 = 8'h1c == io_state_in_13 ? 8'hfc : _GEN_14619; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14621 = 8'h1d == io_state_in_13 ? 8'hf5 : _GEN_14620; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14622 = 8'h1e == io_state_in_13 ? 8'hee : _GEN_14621; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14623 = 8'h1f == io_state_in_13 ? 8'he7 : _GEN_14622; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14624 = 8'h20 == io_state_in_13 ? 8'h3b : _GEN_14623; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14625 = 8'h21 == io_state_in_13 ? 8'h32 : _GEN_14624; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14626 = 8'h22 == io_state_in_13 ? 8'h29 : _GEN_14625; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14627 = 8'h23 == io_state_in_13 ? 8'h20 : _GEN_14626; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14628 = 8'h24 == io_state_in_13 ? 8'h1f : _GEN_14627; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14629 = 8'h25 == io_state_in_13 ? 8'h16 : _GEN_14628; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14630 = 8'h26 == io_state_in_13 ? 8'hd : _GEN_14629; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14631 = 8'h27 == io_state_in_13 ? 8'h4 : _GEN_14630; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14632 = 8'h28 == io_state_in_13 ? 8'h73 : _GEN_14631; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14633 = 8'h29 == io_state_in_13 ? 8'h7a : _GEN_14632; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14634 = 8'h2a == io_state_in_13 ? 8'h61 : _GEN_14633; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14635 = 8'h2b == io_state_in_13 ? 8'h68 : _GEN_14634; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14636 = 8'h2c == io_state_in_13 ? 8'h57 : _GEN_14635; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14637 = 8'h2d == io_state_in_13 ? 8'h5e : _GEN_14636; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14638 = 8'h2e == io_state_in_13 ? 8'h45 : _GEN_14637; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14639 = 8'h2f == io_state_in_13 ? 8'h4c : _GEN_14638; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14640 = 8'h30 == io_state_in_13 ? 8'hab : _GEN_14639; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14641 = 8'h31 == io_state_in_13 ? 8'ha2 : _GEN_14640; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14642 = 8'h32 == io_state_in_13 ? 8'hb9 : _GEN_14641; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14643 = 8'h33 == io_state_in_13 ? 8'hb0 : _GEN_14642; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14644 = 8'h34 == io_state_in_13 ? 8'h8f : _GEN_14643; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14645 = 8'h35 == io_state_in_13 ? 8'h86 : _GEN_14644; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14646 = 8'h36 == io_state_in_13 ? 8'h9d : _GEN_14645; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14647 = 8'h37 == io_state_in_13 ? 8'h94 : _GEN_14646; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14648 = 8'h38 == io_state_in_13 ? 8'he3 : _GEN_14647; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14649 = 8'h39 == io_state_in_13 ? 8'hea : _GEN_14648; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14650 = 8'h3a == io_state_in_13 ? 8'hf1 : _GEN_14649; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14651 = 8'h3b == io_state_in_13 ? 8'hf8 : _GEN_14650; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14652 = 8'h3c == io_state_in_13 ? 8'hc7 : _GEN_14651; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14653 = 8'h3d == io_state_in_13 ? 8'hce : _GEN_14652; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14654 = 8'h3e == io_state_in_13 ? 8'hd5 : _GEN_14653; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14655 = 8'h3f == io_state_in_13 ? 8'hdc : _GEN_14654; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14656 = 8'h40 == io_state_in_13 ? 8'h76 : _GEN_14655; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14657 = 8'h41 == io_state_in_13 ? 8'h7f : _GEN_14656; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14658 = 8'h42 == io_state_in_13 ? 8'h64 : _GEN_14657; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14659 = 8'h43 == io_state_in_13 ? 8'h6d : _GEN_14658; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14660 = 8'h44 == io_state_in_13 ? 8'h52 : _GEN_14659; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14661 = 8'h45 == io_state_in_13 ? 8'h5b : _GEN_14660; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14662 = 8'h46 == io_state_in_13 ? 8'h40 : _GEN_14661; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14663 = 8'h47 == io_state_in_13 ? 8'h49 : _GEN_14662; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14664 = 8'h48 == io_state_in_13 ? 8'h3e : _GEN_14663; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14665 = 8'h49 == io_state_in_13 ? 8'h37 : _GEN_14664; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14666 = 8'h4a == io_state_in_13 ? 8'h2c : _GEN_14665; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14667 = 8'h4b == io_state_in_13 ? 8'h25 : _GEN_14666; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14668 = 8'h4c == io_state_in_13 ? 8'h1a : _GEN_14667; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14669 = 8'h4d == io_state_in_13 ? 8'h13 : _GEN_14668; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14670 = 8'h4e == io_state_in_13 ? 8'h8 : _GEN_14669; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14671 = 8'h4f == io_state_in_13 ? 8'h1 : _GEN_14670; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14672 = 8'h50 == io_state_in_13 ? 8'he6 : _GEN_14671; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14673 = 8'h51 == io_state_in_13 ? 8'hef : _GEN_14672; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14674 = 8'h52 == io_state_in_13 ? 8'hf4 : _GEN_14673; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14675 = 8'h53 == io_state_in_13 ? 8'hfd : _GEN_14674; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14676 = 8'h54 == io_state_in_13 ? 8'hc2 : _GEN_14675; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14677 = 8'h55 == io_state_in_13 ? 8'hcb : _GEN_14676; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14678 = 8'h56 == io_state_in_13 ? 8'hd0 : _GEN_14677; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14679 = 8'h57 == io_state_in_13 ? 8'hd9 : _GEN_14678; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14680 = 8'h58 == io_state_in_13 ? 8'hae : _GEN_14679; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14681 = 8'h59 == io_state_in_13 ? 8'ha7 : _GEN_14680; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14682 = 8'h5a == io_state_in_13 ? 8'hbc : _GEN_14681; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14683 = 8'h5b == io_state_in_13 ? 8'hb5 : _GEN_14682; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14684 = 8'h5c == io_state_in_13 ? 8'h8a : _GEN_14683; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14685 = 8'h5d == io_state_in_13 ? 8'h83 : _GEN_14684; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14686 = 8'h5e == io_state_in_13 ? 8'h98 : _GEN_14685; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14687 = 8'h5f == io_state_in_13 ? 8'h91 : _GEN_14686; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14688 = 8'h60 == io_state_in_13 ? 8'h4d : _GEN_14687; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14689 = 8'h61 == io_state_in_13 ? 8'h44 : _GEN_14688; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14690 = 8'h62 == io_state_in_13 ? 8'h5f : _GEN_14689; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14691 = 8'h63 == io_state_in_13 ? 8'h56 : _GEN_14690; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14692 = 8'h64 == io_state_in_13 ? 8'h69 : _GEN_14691; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14693 = 8'h65 == io_state_in_13 ? 8'h60 : _GEN_14692; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14694 = 8'h66 == io_state_in_13 ? 8'h7b : _GEN_14693; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14695 = 8'h67 == io_state_in_13 ? 8'h72 : _GEN_14694; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14696 = 8'h68 == io_state_in_13 ? 8'h5 : _GEN_14695; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14697 = 8'h69 == io_state_in_13 ? 8'hc : _GEN_14696; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14698 = 8'h6a == io_state_in_13 ? 8'h17 : _GEN_14697; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14699 = 8'h6b == io_state_in_13 ? 8'h1e : _GEN_14698; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14700 = 8'h6c == io_state_in_13 ? 8'h21 : _GEN_14699; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14701 = 8'h6d == io_state_in_13 ? 8'h28 : _GEN_14700; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14702 = 8'h6e == io_state_in_13 ? 8'h33 : _GEN_14701; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14703 = 8'h6f == io_state_in_13 ? 8'h3a : _GEN_14702; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14704 = 8'h70 == io_state_in_13 ? 8'hdd : _GEN_14703; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14705 = 8'h71 == io_state_in_13 ? 8'hd4 : _GEN_14704; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14706 = 8'h72 == io_state_in_13 ? 8'hcf : _GEN_14705; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14707 = 8'h73 == io_state_in_13 ? 8'hc6 : _GEN_14706; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14708 = 8'h74 == io_state_in_13 ? 8'hf9 : _GEN_14707; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14709 = 8'h75 == io_state_in_13 ? 8'hf0 : _GEN_14708; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14710 = 8'h76 == io_state_in_13 ? 8'heb : _GEN_14709; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14711 = 8'h77 == io_state_in_13 ? 8'he2 : _GEN_14710; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14712 = 8'h78 == io_state_in_13 ? 8'h95 : _GEN_14711; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14713 = 8'h79 == io_state_in_13 ? 8'h9c : _GEN_14712; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14714 = 8'h7a == io_state_in_13 ? 8'h87 : _GEN_14713; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14715 = 8'h7b == io_state_in_13 ? 8'h8e : _GEN_14714; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14716 = 8'h7c == io_state_in_13 ? 8'hb1 : _GEN_14715; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14717 = 8'h7d == io_state_in_13 ? 8'hb8 : _GEN_14716; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14718 = 8'h7e == io_state_in_13 ? 8'ha3 : _GEN_14717; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14719 = 8'h7f == io_state_in_13 ? 8'haa : _GEN_14718; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14720 = 8'h80 == io_state_in_13 ? 8'hec : _GEN_14719; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14721 = 8'h81 == io_state_in_13 ? 8'he5 : _GEN_14720; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14722 = 8'h82 == io_state_in_13 ? 8'hfe : _GEN_14721; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14723 = 8'h83 == io_state_in_13 ? 8'hf7 : _GEN_14722; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14724 = 8'h84 == io_state_in_13 ? 8'hc8 : _GEN_14723; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14725 = 8'h85 == io_state_in_13 ? 8'hc1 : _GEN_14724; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14726 = 8'h86 == io_state_in_13 ? 8'hda : _GEN_14725; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14727 = 8'h87 == io_state_in_13 ? 8'hd3 : _GEN_14726; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14728 = 8'h88 == io_state_in_13 ? 8'ha4 : _GEN_14727; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14729 = 8'h89 == io_state_in_13 ? 8'had : _GEN_14728; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14730 = 8'h8a == io_state_in_13 ? 8'hb6 : _GEN_14729; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14731 = 8'h8b == io_state_in_13 ? 8'hbf : _GEN_14730; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14732 = 8'h8c == io_state_in_13 ? 8'h80 : _GEN_14731; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14733 = 8'h8d == io_state_in_13 ? 8'h89 : _GEN_14732; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14734 = 8'h8e == io_state_in_13 ? 8'h92 : _GEN_14733; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14735 = 8'h8f == io_state_in_13 ? 8'h9b : _GEN_14734; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14736 = 8'h90 == io_state_in_13 ? 8'h7c : _GEN_14735; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14737 = 8'h91 == io_state_in_13 ? 8'h75 : _GEN_14736; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14738 = 8'h92 == io_state_in_13 ? 8'h6e : _GEN_14737; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14739 = 8'h93 == io_state_in_13 ? 8'h67 : _GEN_14738; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14740 = 8'h94 == io_state_in_13 ? 8'h58 : _GEN_14739; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14741 = 8'h95 == io_state_in_13 ? 8'h51 : _GEN_14740; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14742 = 8'h96 == io_state_in_13 ? 8'h4a : _GEN_14741; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14743 = 8'h97 == io_state_in_13 ? 8'h43 : _GEN_14742; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14744 = 8'h98 == io_state_in_13 ? 8'h34 : _GEN_14743; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14745 = 8'h99 == io_state_in_13 ? 8'h3d : _GEN_14744; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14746 = 8'h9a == io_state_in_13 ? 8'h26 : _GEN_14745; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14747 = 8'h9b == io_state_in_13 ? 8'h2f : _GEN_14746; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14748 = 8'h9c == io_state_in_13 ? 8'h10 : _GEN_14747; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14749 = 8'h9d == io_state_in_13 ? 8'h19 : _GEN_14748; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14750 = 8'h9e == io_state_in_13 ? 8'h2 : _GEN_14749; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14751 = 8'h9f == io_state_in_13 ? 8'hb : _GEN_14750; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14752 = 8'ha0 == io_state_in_13 ? 8'hd7 : _GEN_14751; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14753 = 8'ha1 == io_state_in_13 ? 8'hde : _GEN_14752; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14754 = 8'ha2 == io_state_in_13 ? 8'hc5 : _GEN_14753; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14755 = 8'ha3 == io_state_in_13 ? 8'hcc : _GEN_14754; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14756 = 8'ha4 == io_state_in_13 ? 8'hf3 : _GEN_14755; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14757 = 8'ha5 == io_state_in_13 ? 8'hfa : _GEN_14756; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14758 = 8'ha6 == io_state_in_13 ? 8'he1 : _GEN_14757; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14759 = 8'ha7 == io_state_in_13 ? 8'he8 : _GEN_14758; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14760 = 8'ha8 == io_state_in_13 ? 8'h9f : _GEN_14759; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14761 = 8'ha9 == io_state_in_13 ? 8'h96 : _GEN_14760; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14762 = 8'haa == io_state_in_13 ? 8'h8d : _GEN_14761; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14763 = 8'hab == io_state_in_13 ? 8'h84 : _GEN_14762; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14764 = 8'hac == io_state_in_13 ? 8'hbb : _GEN_14763; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14765 = 8'had == io_state_in_13 ? 8'hb2 : _GEN_14764; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14766 = 8'hae == io_state_in_13 ? 8'ha9 : _GEN_14765; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14767 = 8'haf == io_state_in_13 ? 8'ha0 : _GEN_14766; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14768 = 8'hb0 == io_state_in_13 ? 8'h47 : _GEN_14767; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14769 = 8'hb1 == io_state_in_13 ? 8'h4e : _GEN_14768; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14770 = 8'hb2 == io_state_in_13 ? 8'h55 : _GEN_14769; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14771 = 8'hb3 == io_state_in_13 ? 8'h5c : _GEN_14770; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14772 = 8'hb4 == io_state_in_13 ? 8'h63 : _GEN_14771; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14773 = 8'hb5 == io_state_in_13 ? 8'h6a : _GEN_14772; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14774 = 8'hb6 == io_state_in_13 ? 8'h71 : _GEN_14773; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14775 = 8'hb7 == io_state_in_13 ? 8'h78 : _GEN_14774; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14776 = 8'hb8 == io_state_in_13 ? 8'hf : _GEN_14775; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14777 = 8'hb9 == io_state_in_13 ? 8'h6 : _GEN_14776; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14778 = 8'hba == io_state_in_13 ? 8'h1d : _GEN_14777; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14779 = 8'hbb == io_state_in_13 ? 8'h14 : _GEN_14778; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14780 = 8'hbc == io_state_in_13 ? 8'h2b : _GEN_14779; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14781 = 8'hbd == io_state_in_13 ? 8'h22 : _GEN_14780; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14782 = 8'hbe == io_state_in_13 ? 8'h39 : _GEN_14781; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14783 = 8'hbf == io_state_in_13 ? 8'h30 : _GEN_14782; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14784 = 8'hc0 == io_state_in_13 ? 8'h9a : _GEN_14783; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14785 = 8'hc1 == io_state_in_13 ? 8'h93 : _GEN_14784; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14786 = 8'hc2 == io_state_in_13 ? 8'h88 : _GEN_14785; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14787 = 8'hc3 == io_state_in_13 ? 8'h81 : _GEN_14786; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14788 = 8'hc4 == io_state_in_13 ? 8'hbe : _GEN_14787; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14789 = 8'hc5 == io_state_in_13 ? 8'hb7 : _GEN_14788; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14790 = 8'hc6 == io_state_in_13 ? 8'hac : _GEN_14789; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14791 = 8'hc7 == io_state_in_13 ? 8'ha5 : _GEN_14790; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14792 = 8'hc8 == io_state_in_13 ? 8'hd2 : _GEN_14791; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14793 = 8'hc9 == io_state_in_13 ? 8'hdb : _GEN_14792; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14794 = 8'hca == io_state_in_13 ? 8'hc0 : _GEN_14793; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14795 = 8'hcb == io_state_in_13 ? 8'hc9 : _GEN_14794; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14796 = 8'hcc == io_state_in_13 ? 8'hf6 : _GEN_14795; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14797 = 8'hcd == io_state_in_13 ? 8'hff : _GEN_14796; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14798 = 8'hce == io_state_in_13 ? 8'he4 : _GEN_14797; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14799 = 8'hcf == io_state_in_13 ? 8'hed : _GEN_14798; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14800 = 8'hd0 == io_state_in_13 ? 8'ha : _GEN_14799; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14801 = 8'hd1 == io_state_in_13 ? 8'h3 : _GEN_14800; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14802 = 8'hd2 == io_state_in_13 ? 8'h18 : _GEN_14801; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14803 = 8'hd3 == io_state_in_13 ? 8'h11 : _GEN_14802; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14804 = 8'hd4 == io_state_in_13 ? 8'h2e : _GEN_14803; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14805 = 8'hd5 == io_state_in_13 ? 8'h27 : _GEN_14804; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14806 = 8'hd6 == io_state_in_13 ? 8'h3c : _GEN_14805; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14807 = 8'hd7 == io_state_in_13 ? 8'h35 : _GEN_14806; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14808 = 8'hd8 == io_state_in_13 ? 8'h42 : _GEN_14807; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14809 = 8'hd9 == io_state_in_13 ? 8'h4b : _GEN_14808; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14810 = 8'hda == io_state_in_13 ? 8'h50 : _GEN_14809; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14811 = 8'hdb == io_state_in_13 ? 8'h59 : _GEN_14810; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14812 = 8'hdc == io_state_in_13 ? 8'h66 : _GEN_14811; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14813 = 8'hdd == io_state_in_13 ? 8'h6f : _GEN_14812; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14814 = 8'hde == io_state_in_13 ? 8'h74 : _GEN_14813; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14815 = 8'hdf == io_state_in_13 ? 8'h7d : _GEN_14814; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14816 = 8'he0 == io_state_in_13 ? 8'ha1 : _GEN_14815; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14817 = 8'he1 == io_state_in_13 ? 8'ha8 : _GEN_14816; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14818 = 8'he2 == io_state_in_13 ? 8'hb3 : _GEN_14817; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14819 = 8'he3 == io_state_in_13 ? 8'hba : _GEN_14818; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14820 = 8'he4 == io_state_in_13 ? 8'h85 : _GEN_14819; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14821 = 8'he5 == io_state_in_13 ? 8'h8c : _GEN_14820; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14822 = 8'he6 == io_state_in_13 ? 8'h97 : _GEN_14821; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14823 = 8'he7 == io_state_in_13 ? 8'h9e : _GEN_14822; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14824 = 8'he8 == io_state_in_13 ? 8'he9 : _GEN_14823; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14825 = 8'he9 == io_state_in_13 ? 8'he0 : _GEN_14824; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14826 = 8'hea == io_state_in_13 ? 8'hfb : _GEN_14825; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14827 = 8'heb == io_state_in_13 ? 8'hf2 : _GEN_14826; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14828 = 8'hec == io_state_in_13 ? 8'hcd : _GEN_14827; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14829 = 8'hed == io_state_in_13 ? 8'hc4 : _GEN_14828; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14830 = 8'hee == io_state_in_13 ? 8'hdf : _GEN_14829; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14831 = 8'hef == io_state_in_13 ? 8'hd6 : _GEN_14830; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14832 = 8'hf0 == io_state_in_13 ? 8'h31 : _GEN_14831; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14833 = 8'hf1 == io_state_in_13 ? 8'h38 : _GEN_14832; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14834 = 8'hf2 == io_state_in_13 ? 8'h23 : _GEN_14833; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14835 = 8'hf3 == io_state_in_13 ? 8'h2a : _GEN_14834; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14836 = 8'hf4 == io_state_in_13 ? 8'h15 : _GEN_14835; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14837 = 8'hf5 == io_state_in_13 ? 8'h1c : _GEN_14836; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14838 = 8'hf6 == io_state_in_13 ? 8'h7 : _GEN_14837; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14839 = 8'hf7 == io_state_in_13 ? 8'he : _GEN_14838; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14840 = 8'hf8 == io_state_in_13 ? 8'h79 : _GEN_14839; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14841 = 8'hf9 == io_state_in_13 ? 8'h70 : _GEN_14840; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14842 = 8'hfa == io_state_in_13 ? 8'h6b : _GEN_14841; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14843 = 8'hfb == io_state_in_13 ? 8'h62 : _GEN_14842; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14844 = 8'hfc == io_state_in_13 ? 8'h5d : _GEN_14843; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14845 = 8'hfd == io_state_in_13 ? 8'h54 : _GEN_14844; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14846 = 8'hfe == io_state_in_13 ? 8'h4f : _GEN_14845; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_14847 = 8'hff == io_state_in_13 ? 8'h46 : _GEN_14846; // @[InvMixColumns.scala 143:{43,43}]
  wire [7:0] _tmp_state_14_T = _GEN_14591 ^ _GEN_14847; // @[InvMixColumns.scala 143:43]
  wire [7:0] _GEN_14849 = 8'h1 == io_state_in_14 ? 8'he : 8'h0; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14850 = 8'h2 == io_state_in_14 ? 8'h1c : _GEN_14849; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14851 = 8'h3 == io_state_in_14 ? 8'h12 : _GEN_14850; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14852 = 8'h4 == io_state_in_14 ? 8'h38 : _GEN_14851; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14853 = 8'h5 == io_state_in_14 ? 8'h36 : _GEN_14852; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14854 = 8'h6 == io_state_in_14 ? 8'h24 : _GEN_14853; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14855 = 8'h7 == io_state_in_14 ? 8'h2a : _GEN_14854; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14856 = 8'h8 == io_state_in_14 ? 8'h70 : _GEN_14855; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14857 = 8'h9 == io_state_in_14 ? 8'h7e : _GEN_14856; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14858 = 8'ha == io_state_in_14 ? 8'h6c : _GEN_14857; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14859 = 8'hb == io_state_in_14 ? 8'h62 : _GEN_14858; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14860 = 8'hc == io_state_in_14 ? 8'h48 : _GEN_14859; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14861 = 8'hd == io_state_in_14 ? 8'h46 : _GEN_14860; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14862 = 8'he == io_state_in_14 ? 8'h54 : _GEN_14861; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14863 = 8'hf == io_state_in_14 ? 8'h5a : _GEN_14862; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14864 = 8'h10 == io_state_in_14 ? 8'he0 : _GEN_14863; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14865 = 8'h11 == io_state_in_14 ? 8'hee : _GEN_14864; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14866 = 8'h12 == io_state_in_14 ? 8'hfc : _GEN_14865; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14867 = 8'h13 == io_state_in_14 ? 8'hf2 : _GEN_14866; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14868 = 8'h14 == io_state_in_14 ? 8'hd8 : _GEN_14867; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14869 = 8'h15 == io_state_in_14 ? 8'hd6 : _GEN_14868; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14870 = 8'h16 == io_state_in_14 ? 8'hc4 : _GEN_14869; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14871 = 8'h17 == io_state_in_14 ? 8'hca : _GEN_14870; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14872 = 8'h18 == io_state_in_14 ? 8'h90 : _GEN_14871; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14873 = 8'h19 == io_state_in_14 ? 8'h9e : _GEN_14872; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14874 = 8'h1a == io_state_in_14 ? 8'h8c : _GEN_14873; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14875 = 8'h1b == io_state_in_14 ? 8'h82 : _GEN_14874; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14876 = 8'h1c == io_state_in_14 ? 8'ha8 : _GEN_14875; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14877 = 8'h1d == io_state_in_14 ? 8'ha6 : _GEN_14876; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14878 = 8'h1e == io_state_in_14 ? 8'hb4 : _GEN_14877; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14879 = 8'h1f == io_state_in_14 ? 8'hba : _GEN_14878; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14880 = 8'h20 == io_state_in_14 ? 8'hdb : _GEN_14879; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14881 = 8'h21 == io_state_in_14 ? 8'hd5 : _GEN_14880; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14882 = 8'h22 == io_state_in_14 ? 8'hc7 : _GEN_14881; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14883 = 8'h23 == io_state_in_14 ? 8'hc9 : _GEN_14882; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14884 = 8'h24 == io_state_in_14 ? 8'he3 : _GEN_14883; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14885 = 8'h25 == io_state_in_14 ? 8'hed : _GEN_14884; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14886 = 8'h26 == io_state_in_14 ? 8'hff : _GEN_14885; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14887 = 8'h27 == io_state_in_14 ? 8'hf1 : _GEN_14886; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14888 = 8'h28 == io_state_in_14 ? 8'hab : _GEN_14887; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14889 = 8'h29 == io_state_in_14 ? 8'ha5 : _GEN_14888; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14890 = 8'h2a == io_state_in_14 ? 8'hb7 : _GEN_14889; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14891 = 8'h2b == io_state_in_14 ? 8'hb9 : _GEN_14890; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14892 = 8'h2c == io_state_in_14 ? 8'h93 : _GEN_14891; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14893 = 8'h2d == io_state_in_14 ? 8'h9d : _GEN_14892; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14894 = 8'h2e == io_state_in_14 ? 8'h8f : _GEN_14893; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14895 = 8'h2f == io_state_in_14 ? 8'h81 : _GEN_14894; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14896 = 8'h30 == io_state_in_14 ? 8'h3b : _GEN_14895; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14897 = 8'h31 == io_state_in_14 ? 8'h35 : _GEN_14896; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14898 = 8'h32 == io_state_in_14 ? 8'h27 : _GEN_14897; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14899 = 8'h33 == io_state_in_14 ? 8'h29 : _GEN_14898; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14900 = 8'h34 == io_state_in_14 ? 8'h3 : _GEN_14899; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14901 = 8'h35 == io_state_in_14 ? 8'hd : _GEN_14900; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14902 = 8'h36 == io_state_in_14 ? 8'h1f : _GEN_14901; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14903 = 8'h37 == io_state_in_14 ? 8'h11 : _GEN_14902; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14904 = 8'h38 == io_state_in_14 ? 8'h4b : _GEN_14903; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14905 = 8'h39 == io_state_in_14 ? 8'h45 : _GEN_14904; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14906 = 8'h3a == io_state_in_14 ? 8'h57 : _GEN_14905; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14907 = 8'h3b == io_state_in_14 ? 8'h59 : _GEN_14906; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14908 = 8'h3c == io_state_in_14 ? 8'h73 : _GEN_14907; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14909 = 8'h3d == io_state_in_14 ? 8'h7d : _GEN_14908; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14910 = 8'h3e == io_state_in_14 ? 8'h6f : _GEN_14909; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14911 = 8'h3f == io_state_in_14 ? 8'h61 : _GEN_14910; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14912 = 8'h40 == io_state_in_14 ? 8'had : _GEN_14911; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14913 = 8'h41 == io_state_in_14 ? 8'ha3 : _GEN_14912; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14914 = 8'h42 == io_state_in_14 ? 8'hb1 : _GEN_14913; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14915 = 8'h43 == io_state_in_14 ? 8'hbf : _GEN_14914; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14916 = 8'h44 == io_state_in_14 ? 8'h95 : _GEN_14915; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14917 = 8'h45 == io_state_in_14 ? 8'h9b : _GEN_14916; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14918 = 8'h46 == io_state_in_14 ? 8'h89 : _GEN_14917; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14919 = 8'h47 == io_state_in_14 ? 8'h87 : _GEN_14918; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14920 = 8'h48 == io_state_in_14 ? 8'hdd : _GEN_14919; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14921 = 8'h49 == io_state_in_14 ? 8'hd3 : _GEN_14920; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14922 = 8'h4a == io_state_in_14 ? 8'hc1 : _GEN_14921; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14923 = 8'h4b == io_state_in_14 ? 8'hcf : _GEN_14922; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14924 = 8'h4c == io_state_in_14 ? 8'he5 : _GEN_14923; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14925 = 8'h4d == io_state_in_14 ? 8'heb : _GEN_14924; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14926 = 8'h4e == io_state_in_14 ? 8'hf9 : _GEN_14925; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14927 = 8'h4f == io_state_in_14 ? 8'hf7 : _GEN_14926; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14928 = 8'h50 == io_state_in_14 ? 8'h4d : _GEN_14927; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14929 = 8'h51 == io_state_in_14 ? 8'h43 : _GEN_14928; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14930 = 8'h52 == io_state_in_14 ? 8'h51 : _GEN_14929; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14931 = 8'h53 == io_state_in_14 ? 8'h5f : _GEN_14930; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14932 = 8'h54 == io_state_in_14 ? 8'h75 : _GEN_14931; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14933 = 8'h55 == io_state_in_14 ? 8'h7b : _GEN_14932; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14934 = 8'h56 == io_state_in_14 ? 8'h69 : _GEN_14933; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14935 = 8'h57 == io_state_in_14 ? 8'h67 : _GEN_14934; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14936 = 8'h58 == io_state_in_14 ? 8'h3d : _GEN_14935; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14937 = 8'h59 == io_state_in_14 ? 8'h33 : _GEN_14936; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14938 = 8'h5a == io_state_in_14 ? 8'h21 : _GEN_14937; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14939 = 8'h5b == io_state_in_14 ? 8'h2f : _GEN_14938; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14940 = 8'h5c == io_state_in_14 ? 8'h5 : _GEN_14939; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14941 = 8'h5d == io_state_in_14 ? 8'hb : _GEN_14940; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14942 = 8'h5e == io_state_in_14 ? 8'h19 : _GEN_14941; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14943 = 8'h5f == io_state_in_14 ? 8'h17 : _GEN_14942; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14944 = 8'h60 == io_state_in_14 ? 8'h76 : _GEN_14943; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14945 = 8'h61 == io_state_in_14 ? 8'h78 : _GEN_14944; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14946 = 8'h62 == io_state_in_14 ? 8'h6a : _GEN_14945; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14947 = 8'h63 == io_state_in_14 ? 8'h64 : _GEN_14946; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14948 = 8'h64 == io_state_in_14 ? 8'h4e : _GEN_14947; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14949 = 8'h65 == io_state_in_14 ? 8'h40 : _GEN_14948; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14950 = 8'h66 == io_state_in_14 ? 8'h52 : _GEN_14949; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14951 = 8'h67 == io_state_in_14 ? 8'h5c : _GEN_14950; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14952 = 8'h68 == io_state_in_14 ? 8'h6 : _GEN_14951; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14953 = 8'h69 == io_state_in_14 ? 8'h8 : _GEN_14952; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14954 = 8'h6a == io_state_in_14 ? 8'h1a : _GEN_14953; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14955 = 8'h6b == io_state_in_14 ? 8'h14 : _GEN_14954; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14956 = 8'h6c == io_state_in_14 ? 8'h3e : _GEN_14955; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14957 = 8'h6d == io_state_in_14 ? 8'h30 : _GEN_14956; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14958 = 8'h6e == io_state_in_14 ? 8'h22 : _GEN_14957; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14959 = 8'h6f == io_state_in_14 ? 8'h2c : _GEN_14958; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14960 = 8'h70 == io_state_in_14 ? 8'h96 : _GEN_14959; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14961 = 8'h71 == io_state_in_14 ? 8'h98 : _GEN_14960; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14962 = 8'h72 == io_state_in_14 ? 8'h8a : _GEN_14961; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14963 = 8'h73 == io_state_in_14 ? 8'h84 : _GEN_14962; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14964 = 8'h74 == io_state_in_14 ? 8'hae : _GEN_14963; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14965 = 8'h75 == io_state_in_14 ? 8'ha0 : _GEN_14964; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14966 = 8'h76 == io_state_in_14 ? 8'hb2 : _GEN_14965; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14967 = 8'h77 == io_state_in_14 ? 8'hbc : _GEN_14966; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14968 = 8'h78 == io_state_in_14 ? 8'he6 : _GEN_14967; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14969 = 8'h79 == io_state_in_14 ? 8'he8 : _GEN_14968; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14970 = 8'h7a == io_state_in_14 ? 8'hfa : _GEN_14969; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14971 = 8'h7b == io_state_in_14 ? 8'hf4 : _GEN_14970; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14972 = 8'h7c == io_state_in_14 ? 8'hde : _GEN_14971; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14973 = 8'h7d == io_state_in_14 ? 8'hd0 : _GEN_14972; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14974 = 8'h7e == io_state_in_14 ? 8'hc2 : _GEN_14973; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14975 = 8'h7f == io_state_in_14 ? 8'hcc : _GEN_14974; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14976 = 8'h80 == io_state_in_14 ? 8'h41 : _GEN_14975; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14977 = 8'h81 == io_state_in_14 ? 8'h4f : _GEN_14976; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14978 = 8'h82 == io_state_in_14 ? 8'h5d : _GEN_14977; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14979 = 8'h83 == io_state_in_14 ? 8'h53 : _GEN_14978; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14980 = 8'h84 == io_state_in_14 ? 8'h79 : _GEN_14979; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14981 = 8'h85 == io_state_in_14 ? 8'h77 : _GEN_14980; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14982 = 8'h86 == io_state_in_14 ? 8'h65 : _GEN_14981; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14983 = 8'h87 == io_state_in_14 ? 8'h6b : _GEN_14982; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14984 = 8'h88 == io_state_in_14 ? 8'h31 : _GEN_14983; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14985 = 8'h89 == io_state_in_14 ? 8'h3f : _GEN_14984; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14986 = 8'h8a == io_state_in_14 ? 8'h2d : _GEN_14985; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14987 = 8'h8b == io_state_in_14 ? 8'h23 : _GEN_14986; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14988 = 8'h8c == io_state_in_14 ? 8'h9 : _GEN_14987; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14989 = 8'h8d == io_state_in_14 ? 8'h7 : _GEN_14988; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14990 = 8'h8e == io_state_in_14 ? 8'h15 : _GEN_14989; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14991 = 8'h8f == io_state_in_14 ? 8'h1b : _GEN_14990; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14992 = 8'h90 == io_state_in_14 ? 8'ha1 : _GEN_14991; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14993 = 8'h91 == io_state_in_14 ? 8'haf : _GEN_14992; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14994 = 8'h92 == io_state_in_14 ? 8'hbd : _GEN_14993; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14995 = 8'h93 == io_state_in_14 ? 8'hb3 : _GEN_14994; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14996 = 8'h94 == io_state_in_14 ? 8'h99 : _GEN_14995; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14997 = 8'h95 == io_state_in_14 ? 8'h97 : _GEN_14996; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14998 = 8'h96 == io_state_in_14 ? 8'h85 : _GEN_14997; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_14999 = 8'h97 == io_state_in_14 ? 8'h8b : _GEN_14998; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15000 = 8'h98 == io_state_in_14 ? 8'hd1 : _GEN_14999; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15001 = 8'h99 == io_state_in_14 ? 8'hdf : _GEN_15000; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15002 = 8'h9a == io_state_in_14 ? 8'hcd : _GEN_15001; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15003 = 8'h9b == io_state_in_14 ? 8'hc3 : _GEN_15002; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15004 = 8'h9c == io_state_in_14 ? 8'he9 : _GEN_15003; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15005 = 8'h9d == io_state_in_14 ? 8'he7 : _GEN_15004; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15006 = 8'h9e == io_state_in_14 ? 8'hf5 : _GEN_15005; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15007 = 8'h9f == io_state_in_14 ? 8'hfb : _GEN_15006; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15008 = 8'ha0 == io_state_in_14 ? 8'h9a : _GEN_15007; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15009 = 8'ha1 == io_state_in_14 ? 8'h94 : _GEN_15008; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15010 = 8'ha2 == io_state_in_14 ? 8'h86 : _GEN_15009; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15011 = 8'ha3 == io_state_in_14 ? 8'h88 : _GEN_15010; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15012 = 8'ha4 == io_state_in_14 ? 8'ha2 : _GEN_15011; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15013 = 8'ha5 == io_state_in_14 ? 8'hac : _GEN_15012; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15014 = 8'ha6 == io_state_in_14 ? 8'hbe : _GEN_15013; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15015 = 8'ha7 == io_state_in_14 ? 8'hb0 : _GEN_15014; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15016 = 8'ha8 == io_state_in_14 ? 8'hea : _GEN_15015; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15017 = 8'ha9 == io_state_in_14 ? 8'he4 : _GEN_15016; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15018 = 8'haa == io_state_in_14 ? 8'hf6 : _GEN_15017; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15019 = 8'hab == io_state_in_14 ? 8'hf8 : _GEN_15018; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15020 = 8'hac == io_state_in_14 ? 8'hd2 : _GEN_15019; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15021 = 8'had == io_state_in_14 ? 8'hdc : _GEN_15020; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15022 = 8'hae == io_state_in_14 ? 8'hce : _GEN_15021; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15023 = 8'haf == io_state_in_14 ? 8'hc0 : _GEN_15022; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15024 = 8'hb0 == io_state_in_14 ? 8'h7a : _GEN_15023; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15025 = 8'hb1 == io_state_in_14 ? 8'h74 : _GEN_15024; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15026 = 8'hb2 == io_state_in_14 ? 8'h66 : _GEN_15025; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15027 = 8'hb3 == io_state_in_14 ? 8'h68 : _GEN_15026; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15028 = 8'hb4 == io_state_in_14 ? 8'h42 : _GEN_15027; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15029 = 8'hb5 == io_state_in_14 ? 8'h4c : _GEN_15028; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15030 = 8'hb6 == io_state_in_14 ? 8'h5e : _GEN_15029; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15031 = 8'hb7 == io_state_in_14 ? 8'h50 : _GEN_15030; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15032 = 8'hb8 == io_state_in_14 ? 8'ha : _GEN_15031; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15033 = 8'hb9 == io_state_in_14 ? 8'h4 : _GEN_15032; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15034 = 8'hba == io_state_in_14 ? 8'h16 : _GEN_15033; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15035 = 8'hbb == io_state_in_14 ? 8'h18 : _GEN_15034; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15036 = 8'hbc == io_state_in_14 ? 8'h32 : _GEN_15035; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15037 = 8'hbd == io_state_in_14 ? 8'h3c : _GEN_15036; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15038 = 8'hbe == io_state_in_14 ? 8'h2e : _GEN_15037; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15039 = 8'hbf == io_state_in_14 ? 8'h20 : _GEN_15038; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15040 = 8'hc0 == io_state_in_14 ? 8'hec : _GEN_15039; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15041 = 8'hc1 == io_state_in_14 ? 8'he2 : _GEN_15040; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15042 = 8'hc2 == io_state_in_14 ? 8'hf0 : _GEN_15041; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15043 = 8'hc3 == io_state_in_14 ? 8'hfe : _GEN_15042; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15044 = 8'hc4 == io_state_in_14 ? 8'hd4 : _GEN_15043; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15045 = 8'hc5 == io_state_in_14 ? 8'hda : _GEN_15044; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15046 = 8'hc6 == io_state_in_14 ? 8'hc8 : _GEN_15045; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15047 = 8'hc7 == io_state_in_14 ? 8'hc6 : _GEN_15046; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15048 = 8'hc8 == io_state_in_14 ? 8'h9c : _GEN_15047; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15049 = 8'hc9 == io_state_in_14 ? 8'h92 : _GEN_15048; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15050 = 8'hca == io_state_in_14 ? 8'h80 : _GEN_15049; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15051 = 8'hcb == io_state_in_14 ? 8'h8e : _GEN_15050; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15052 = 8'hcc == io_state_in_14 ? 8'ha4 : _GEN_15051; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15053 = 8'hcd == io_state_in_14 ? 8'haa : _GEN_15052; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15054 = 8'hce == io_state_in_14 ? 8'hb8 : _GEN_15053; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15055 = 8'hcf == io_state_in_14 ? 8'hb6 : _GEN_15054; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15056 = 8'hd0 == io_state_in_14 ? 8'hc : _GEN_15055; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15057 = 8'hd1 == io_state_in_14 ? 8'h2 : _GEN_15056; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15058 = 8'hd2 == io_state_in_14 ? 8'h10 : _GEN_15057; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15059 = 8'hd3 == io_state_in_14 ? 8'h1e : _GEN_15058; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15060 = 8'hd4 == io_state_in_14 ? 8'h34 : _GEN_15059; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15061 = 8'hd5 == io_state_in_14 ? 8'h3a : _GEN_15060; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15062 = 8'hd6 == io_state_in_14 ? 8'h28 : _GEN_15061; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15063 = 8'hd7 == io_state_in_14 ? 8'h26 : _GEN_15062; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15064 = 8'hd8 == io_state_in_14 ? 8'h7c : _GEN_15063; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15065 = 8'hd9 == io_state_in_14 ? 8'h72 : _GEN_15064; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15066 = 8'hda == io_state_in_14 ? 8'h60 : _GEN_15065; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15067 = 8'hdb == io_state_in_14 ? 8'h6e : _GEN_15066; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15068 = 8'hdc == io_state_in_14 ? 8'h44 : _GEN_15067; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15069 = 8'hdd == io_state_in_14 ? 8'h4a : _GEN_15068; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15070 = 8'hde == io_state_in_14 ? 8'h58 : _GEN_15069; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15071 = 8'hdf == io_state_in_14 ? 8'h56 : _GEN_15070; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15072 = 8'he0 == io_state_in_14 ? 8'h37 : _GEN_15071; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15073 = 8'he1 == io_state_in_14 ? 8'h39 : _GEN_15072; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15074 = 8'he2 == io_state_in_14 ? 8'h2b : _GEN_15073; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15075 = 8'he3 == io_state_in_14 ? 8'h25 : _GEN_15074; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15076 = 8'he4 == io_state_in_14 ? 8'hf : _GEN_15075; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15077 = 8'he5 == io_state_in_14 ? 8'h1 : _GEN_15076; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15078 = 8'he6 == io_state_in_14 ? 8'h13 : _GEN_15077; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15079 = 8'he7 == io_state_in_14 ? 8'h1d : _GEN_15078; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15080 = 8'he8 == io_state_in_14 ? 8'h47 : _GEN_15079; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15081 = 8'he9 == io_state_in_14 ? 8'h49 : _GEN_15080; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15082 = 8'hea == io_state_in_14 ? 8'h5b : _GEN_15081; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15083 = 8'heb == io_state_in_14 ? 8'h55 : _GEN_15082; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15084 = 8'hec == io_state_in_14 ? 8'h7f : _GEN_15083; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15085 = 8'hed == io_state_in_14 ? 8'h71 : _GEN_15084; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15086 = 8'hee == io_state_in_14 ? 8'h63 : _GEN_15085; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15087 = 8'hef == io_state_in_14 ? 8'h6d : _GEN_15086; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15088 = 8'hf0 == io_state_in_14 ? 8'hd7 : _GEN_15087; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15089 = 8'hf1 == io_state_in_14 ? 8'hd9 : _GEN_15088; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15090 = 8'hf2 == io_state_in_14 ? 8'hcb : _GEN_15089; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15091 = 8'hf3 == io_state_in_14 ? 8'hc5 : _GEN_15090; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15092 = 8'hf4 == io_state_in_14 ? 8'hef : _GEN_15091; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15093 = 8'hf5 == io_state_in_14 ? 8'he1 : _GEN_15092; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15094 = 8'hf6 == io_state_in_14 ? 8'hf3 : _GEN_15093; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15095 = 8'hf7 == io_state_in_14 ? 8'hfd : _GEN_15094; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15096 = 8'hf8 == io_state_in_14 ? 8'ha7 : _GEN_15095; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15097 = 8'hf9 == io_state_in_14 ? 8'ha9 : _GEN_15096; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15098 = 8'hfa == io_state_in_14 ? 8'hbb : _GEN_15097; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15099 = 8'hfb == io_state_in_14 ? 8'hb5 : _GEN_15098; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15100 = 8'hfc == io_state_in_14 ? 8'h9f : _GEN_15099; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15101 = 8'hfd == io_state_in_14 ? 8'h91 : _GEN_15100; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15102 = 8'hfe == io_state_in_14 ? 8'h83 : _GEN_15101; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _GEN_15103 = 8'hff == io_state_in_14 ? 8'h8d : _GEN_15102; // @[InvMixColumns.scala 143:{68,68}]
  wire [7:0] _tmp_state_14_T_1 = _tmp_state_14_T ^ _GEN_15103; // @[InvMixColumns.scala 143:68]
  wire [7:0] _GEN_15105 = 8'h1 == io_state_in_15 ? 8'hb : 8'h0; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15106 = 8'h2 == io_state_in_15 ? 8'h16 : _GEN_15105; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15107 = 8'h3 == io_state_in_15 ? 8'h1d : _GEN_15106; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15108 = 8'h4 == io_state_in_15 ? 8'h2c : _GEN_15107; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15109 = 8'h5 == io_state_in_15 ? 8'h27 : _GEN_15108; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15110 = 8'h6 == io_state_in_15 ? 8'h3a : _GEN_15109; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15111 = 8'h7 == io_state_in_15 ? 8'h31 : _GEN_15110; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15112 = 8'h8 == io_state_in_15 ? 8'h58 : _GEN_15111; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15113 = 8'h9 == io_state_in_15 ? 8'h53 : _GEN_15112; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15114 = 8'ha == io_state_in_15 ? 8'h4e : _GEN_15113; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15115 = 8'hb == io_state_in_15 ? 8'h45 : _GEN_15114; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15116 = 8'hc == io_state_in_15 ? 8'h74 : _GEN_15115; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15117 = 8'hd == io_state_in_15 ? 8'h7f : _GEN_15116; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15118 = 8'he == io_state_in_15 ? 8'h62 : _GEN_15117; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15119 = 8'hf == io_state_in_15 ? 8'h69 : _GEN_15118; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15120 = 8'h10 == io_state_in_15 ? 8'hb0 : _GEN_15119; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15121 = 8'h11 == io_state_in_15 ? 8'hbb : _GEN_15120; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15122 = 8'h12 == io_state_in_15 ? 8'ha6 : _GEN_15121; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15123 = 8'h13 == io_state_in_15 ? 8'had : _GEN_15122; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15124 = 8'h14 == io_state_in_15 ? 8'h9c : _GEN_15123; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15125 = 8'h15 == io_state_in_15 ? 8'h97 : _GEN_15124; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15126 = 8'h16 == io_state_in_15 ? 8'h8a : _GEN_15125; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15127 = 8'h17 == io_state_in_15 ? 8'h81 : _GEN_15126; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15128 = 8'h18 == io_state_in_15 ? 8'he8 : _GEN_15127; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15129 = 8'h19 == io_state_in_15 ? 8'he3 : _GEN_15128; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15130 = 8'h1a == io_state_in_15 ? 8'hfe : _GEN_15129; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15131 = 8'h1b == io_state_in_15 ? 8'hf5 : _GEN_15130; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15132 = 8'h1c == io_state_in_15 ? 8'hc4 : _GEN_15131; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15133 = 8'h1d == io_state_in_15 ? 8'hcf : _GEN_15132; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15134 = 8'h1e == io_state_in_15 ? 8'hd2 : _GEN_15133; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15135 = 8'h1f == io_state_in_15 ? 8'hd9 : _GEN_15134; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15136 = 8'h20 == io_state_in_15 ? 8'h7b : _GEN_15135; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15137 = 8'h21 == io_state_in_15 ? 8'h70 : _GEN_15136; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15138 = 8'h22 == io_state_in_15 ? 8'h6d : _GEN_15137; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15139 = 8'h23 == io_state_in_15 ? 8'h66 : _GEN_15138; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15140 = 8'h24 == io_state_in_15 ? 8'h57 : _GEN_15139; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15141 = 8'h25 == io_state_in_15 ? 8'h5c : _GEN_15140; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15142 = 8'h26 == io_state_in_15 ? 8'h41 : _GEN_15141; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15143 = 8'h27 == io_state_in_15 ? 8'h4a : _GEN_15142; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15144 = 8'h28 == io_state_in_15 ? 8'h23 : _GEN_15143; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15145 = 8'h29 == io_state_in_15 ? 8'h28 : _GEN_15144; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15146 = 8'h2a == io_state_in_15 ? 8'h35 : _GEN_15145; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15147 = 8'h2b == io_state_in_15 ? 8'h3e : _GEN_15146; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15148 = 8'h2c == io_state_in_15 ? 8'hf : _GEN_15147; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15149 = 8'h2d == io_state_in_15 ? 8'h4 : _GEN_15148; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15150 = 8'h2e == io_state_in_15 ? 8'h19 : _GEN_15149; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15151 = 8'h2f == io_state_in_15 ? 8'h12 : _GEN_15150; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15152 = 8'h30 == io_state_in_15 ? 8'hcb : _GEN_15151; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15153 = 8'h31 == io_state_in_15 ? 8'hc0 : _GEN_15152; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15154 = 8'h32 == io_state_in_15 ? 8'hdd : _GEN_15153; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15155 = 8'h33 == io_state_in_15 ? 8'hd6 : _GEN_15154; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15156 = 8'h34 == io_state_in_15 ? 8'he7 : _GEN_15155; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15157 = 8'h35 == io_state_in_15 ? 8'hec : _GEN_15156; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15158 = 8'h36 == io_state_in_15 ? 8'hf1 : _GEN_15157; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15159 = 8'h37 == io_state_in_15 ? 8'hfa : _GEN_15158; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15160 = 8'h38 == io_state_in_15 ? 8'h93 : _GEN_15159; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15161 = 8'h39 == io_state_in_15 ? 8'h98 : _GEN_15160; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15162 = 8'h3a == io_state_in_15 ? 8'h85 : _GEN_15161; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15163 = 8'h3b == io_state_in_15 ? 8'h8e : _GEN_15162; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15164 = 8'h3c == io_state_in_15 ? 8'hbf : _GEN_15163; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15165 = 8'h3d == io_state_in_15 ? 8'hb4 : _GEN_15164; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15166 = 8'h3e == io_state_in_15 ? 8'ha9 : _GEN_15165; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15167 = 8'h3f == io_state_in_15 ? 8'ha2 : _GEN_15166; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15168 = 8'h40 == io_state_in_15 ? 8'hf6 : _GEN_15167; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15169 = 8'h41 == io_state_in_15 ? 8'hfd : _GEN_15168; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15170 = 8'h42 == io_state_in_15 ? 8'he0 : _GEN_15169; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15171 = 8'h43 == io_state_in_15 ? 8'heb : _GEN_15170; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15172 = 8'h44 == io_state_in_15 ? 8'hda : _GEN_15171; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15173 = 8'h45 == io_state_in_15 ? 8'hd1 : _GEN_15172; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15174 = 8'h46 == io_state_in_15 ? 8'hcc : _GEN_15173; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15175 = 8'h47 == io_state_in_15 ? 8'hc7 : _GEN_15174; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15176 = 8'h48 == io_state_in_15 ? 8'hae : _GEN_15175; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15177 = 8'h49 == io_state_in_15 ? 8'ha5 : _GEN_15176; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15178 = 8'h4a == io_state_in_15 ? 8'hb8 : _GEN_15177; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15179 = 8'h4b == io_state_in_15 ? 8'hb3 : _GEN_15178; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15180 = 8'h4c == io_state_in_15 ? 8'h82 : _GEN_15179; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15181 = 8'h4d == io_state_in_15 ? 8'h89 : _GEN_15180; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15182 = 8'h4e == io_state_in_15 ? 8'h94 : _GEN_15181; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15183 = 8'h4f == io_state_in_15 ? 8'h9f : _GEN_15182; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15184 = 8'h50 == io_state_in_15 ? 8'h46 : _GEN_15183; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15185 = 8'h51 == io_state_in_15 ? 8'h4d : _GEN_15184; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15186 = 8'h52 == io_state_in_15 ? 8'h50 : _GEN_15185; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15187 = 8'h53 == io_state_in_15 ? 8'h5b : _GEN_15186; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15188 = 8'h54 == io_state_in_15 ? 8'h6a : _GEN_15187; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15189 = 8'h55 == io_state_in_15 ? 8'h61 : _GEN_15188; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15190 = 8'h56 == io_state_in_15 ? 8'h7c : _GEN_15189; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15191 = 8'h57 == io_state_in_15 ? 8'h77 : _GEN_15190; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15192 = 8'h58 == io_state_in_15 ? 8'h1e : _GEN_15191; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15193 = 8'h59 == io_state_in_15 ? 8'h15 : _GEN_15192; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15194 = 8'h5a == io_state_in_15 ? 8'h8 : _GEN_15193; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15195 = 8'h5b == io_state_in_15 ? 8'h3 : _GEN_15194; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15196 = 8'h5c == io_state_in_15 ? 8'h32 : _GEN_15195; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15197 = 8'h5d == io_state_in_15 ? 8'h39 : _GEN_15196; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15198 = 8'h5e == io_state_in_15 ? 8'h24 : _GEN_15197; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15199 = 8'h5f == io_state_in_15 ? 8'h2f : _GEN_15198; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15200 = 8'h60 == io_state_in_15 ? 8'h8d : _GEN_15199; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15201 = 8'h61 == io_state_in_15 ? 8'h86 : _GEN_15200; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15202 = 8'h62 == io_state_in_15 ? 8'h9b : _GEN_15201; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15203 = 8'h63 == io_state_in_15 ? 8'h90 : _GEN_15202; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15204 = 8'h64 == io_state_in_15 ? 8'ha1 : _GEN_15203; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15205 = 8'h65 == io_state_in_15 ? 8'haa : _GEN_15204; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15206 = 8'h66 == io_state_in_15 ? 8'hb7 : _GEN_15205; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15207 = 8'h67 == io_state_in_15 ? 8'hbc : _GEN_15206; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15208 = 8'h68 == io_state_in_15 ? 8'hd5 : _GEN_15207; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15209 = 8'h69 == io_state_in_15 ? 8'hde : _GEN_15208; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15210 = 8'h6a == io_state_in_15 ? 8'hc3 : _GEN_15209; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15211 = 8'h6b == io_state_in_15 ? 8'hc8 : _GEN_15210; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15212 = 8'h6c == io_state_in_15 ? 8'hf9 : _GEN_15211; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15213 = 8'h6d == io_state_in_15 ? 8'hf2 : _GEN_15212; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15214 = 8'h6e == io_state_in_15 ? 8'hef : _GEN_15213; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15215 = 8'h6f == io_state_in_15 ? 8'he4 : _GEN_15214; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15216 = 8'h70 == io_state_in_15 ? 8'h3d : _GEN_15215; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15217 = 8'h71 == io_state_in_15 ? 8'h36 : _GEN_15216; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15218 = 8'h72 == io_state_in_15 ? 8'h2b : _GEN_15217; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15219 = 8'h73 == io_state_in_15 ? 8'h20 : _GEN_15218; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15220 = 8'h74 == io_state_in_15 ? 8'h11 : _GEN_15219; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15221 = 8'h75 == io_state_in_15 ? 8'h1a : _GEN_15220; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15222 = 8'h76 == io_state_in_15 ? 8'h7 : _GEN_15221; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15223 = 8'h77 == io_state_in_15 ? 8'hc : _GEN_15222; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15224 = 8'h78 == io_state_in_15 ? 8'h65 : _GEN_15223; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15225 = 8'h79 == io_state_in_15 ? 8'h6e : _GEN_15224; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15226 = 8'h7a == io_state_in_15 ? 8'h73 : _GEN_15225; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15227 = 8'h7b == io_state_in_15 ? 8'h78 : _GEN_15226; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15228 = 8'h7c == io_state_in_15 ? 8'h49 : _GEN_15227; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15229 = 8'h7d == io_state_in_15 ? 8'h42 : _GEN_15228; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15230 = 8'h7e == io_state_in_15 ? 8'h5f : _GEN_15229; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15231 = 8'h7f == io_state_in_15 ? 8'h54 : _GEN_15230; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15232 = 8'h80 == io_state_in_15 ? 8'hf7 : _GEN_15231; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15233 = 8'h81 == io_state_in_15 ? 8'hfc : _GEN_15232; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15234 = 8'h82 == io_state_in_15 ? 8'he1 : _GEN_15233; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15235 = 8'h83 == io_state_in_15 ? 8'hea : _GEN_15234; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15236 = 8'h84 == io_state_in_15 ? 8'hdb : _GEN_15235; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15237 = 8'h85 == io_state_in_15 ? 8'hd0 : _GEN_15236; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15238 = 8'h86 == io_state_in_15 ? 8'hcd : _GEN_15237; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15239 = 8'h87 == io_state_in_15 ? 8'hc6 : _GEN_15238; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15240 = 8'h88 == io_state_in_15 ? 8'haf : _GEN_15239; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15241 = 8'h89 == io_state_in_15 ? 8'ha4 : _GEN_15240; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15242 = 8'h8a == io_state_in_15 ? 8'hb9 : _GEN_15241; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15243 = 8'h8b == io_state_in_15 ? 8'hb2 : _GEN_15242; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15244 = 8'h8c == io_state_in_15 ? 8'h83 : _GEN_15243; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15245 = 8'h8d == io_state_in_15 ? 8'h88 : _GEN_15244; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15246 = 8'h8e == io_state_in_15 ? 8'h95 : _GEN_15245; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15247 = 8'h8f == io_state_in_15 ? 8'h9e : _GEN_15246; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15248 = 8'h90 == io_state_in_15 ? 8'h47 : _GEN_15247; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15249 = 8'h91 == io_state_in_15 ? 8'h4c : _GEN_15248; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15250 = 8'h92 == io_state_in_15 ? 8'h51 : _GEN_15249; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15251 = 8'h93 == io_state_in_15 ? 8'h5a : _GEN_15250; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15252 = 8'h94 == io_state_in_15 ? 8'h6b : _GEN_15251; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15253 = 8'h95 == io_state_in_15 ? 8'h60 : _GEN_15252; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15254 = 8'h96 == io_state_in_15 ? 8'h7d : _GEN_15253; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15255 = 8'h97 == io_state_in_15 ? 8'h76 : _GEN_15254; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15256 = 8'h98 == io_state_in_15 ? 8'h1f : _GEN_15255; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15257 = 8'h99 == io_state_in_15 ? 8'h14 : _GEN_15256; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15258 = 8'h9a == io_state_in_15 ? 8'h9 : _GEN_15257; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15259 = 8'h9b == io_state_in_15 ? 8'h2 : _GEN_15258; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15260 = 8'h9c == io_state_in_15 ? 8'h33 : _GEN_15259; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15261 = 8'h9d == io_state_in_15 ? 8'h38 : _GEN_15260; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15262 = 8'h9e == io_state_in_15 ? 8'h25 : _GEN_15261; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15263 = 8'h9f == io_state_in_15 ? 8'h2e : _GEN_15262; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15264 = 8'ha0 == io_state_in_15 ? 8'h8c : _GEN_15263; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15265 = 8'ha1 == io_state_in_15 ? 8'h87 : _GEN_15264; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15266 = 8'ha2 == io_state_in_15 ? 8'h9a : _GEN_15265; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15267 = 8'ha3 == io_state_in_15 ? 8'h91 : _GEN_15266; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15268 = 8'ha4 == io_state_in_15 ? 8'ha0 : _GEN_15267; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15269 = 8'ha5 == io_state_in_15 ? 8'hab : _GEN_15268; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15270 = 8'ha6 == io_state_in_15 ? 8'hb6 : _GEN_15269; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15271 = 8'ha7 == io_state_in_15 ? 8'hbd : _GEN_15270; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15272 = 8'ha8 == io_state_in_15 ? 8'hd4 : _GEN_15271; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15273 = 8'ha9 == io_state_in_15 ? 8'hdf : _GEN_15272; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15274 = 8'haa == io_state_in_15 ? 8'hc2 : _GEN_15273; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15275 = 8'hab == io_state_in_15 ? 8'hc9 : _GEN_15274; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15276 = 8'hac == io_state_in_15 ? 8'hf8 : _GEN_15275; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15277 = 8'had == io_state_in_15 ? 8'hf3 : _GEN_15276; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15278 = 8'hae == io_state_in_15 ? 8'hee : _GEN_15277; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15279 = 8'haf == io_state_in_15 ? 8'he5 : _GEN_15278; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15280 = 8'hb0 == io_state_in_15 ? 8'h3c : _GEN_15279; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15281 = 8'hb1 == io_state_in_15 ? 8'h37 : _GEN_15280; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15282 = 8'hb2 == io_state_in_15 ? 8'h2a : _GEN_15281; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15283 = 8'hb3 == io_state_in_15 ? 8'h21 : _GEN_15282; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15284 = 8'hb4 == io_state_in_15 ? 8'h10 : _GEN_15283; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15285 = 8'hb5 == io_state_in_15 ? 8'h1b : _GEN_15284; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15286 = 8'hb6 == io_state_in_15 ? 8'h6 : _GEN_15285; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15287 = 8'hb7 == io_state_in_15 ? 8'hd : _GEN_15286; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15288 = 8'hb8 == io_state_in_15 ? 8'h64 : _GEN_15287; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15289 = 8'hb9 == io_state_in_15 ? 8'h6f : _GEN_15288; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15290 = 8'hba == io_state_in_15 ? 8'h72 : _GEN_15289; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15291 = 8'hbb == io_state_in_15 ? 8'h79 : _GEN_15290; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15292 = 8'hbc == io_state_in_15 ? 8'h48 : _GEN_15291; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15293 = 8'hbd == io_state_in_15 ? 8'h43 : _GEN_15292; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15294 = 8'hbe == io_state_in_15 ? 8'h5e : _GEN_15293; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15295 = 8'hbf == io_state_in_15 ? 8'h55 : _GEN_15294; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15296 = 8'hc0 == io_state_in_15 ? 8'h1 : _GEN_15295; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15297 = 8'hc1 == io_state_in_15 ? 8'ha : _GEN_15296; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15298 = 8'hc2 == io_state_in_15 ? 8'h17 : _GEN_15297; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15299 = 8'hc3 == io_state_in_15 ? 8'h1c : _GEN_15298; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15300 = 8'hc4 == io_state_in_15 ? 8'h2d : _GEN_15299; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15301 = 8'hc5 == io_state_in_15 ? 8'h26 : _GEN_15300; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15302 = 8'hc6 == io_state_in_15 ? 8'h3b : _GEN_15301; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15303 = 8'hc7 == io_state_in_15 ? 8'h30 : _GEN_15302; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15304 = 8'hc8 == io_state_in_15 ? 8'h59 : _GEN_15303; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15305 = 8'hc9 == io_state_in_15 ? 8'h52 : _GEN_15304; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15306 = 8'hca == io_state_in_15 ? 8'h4f : _GEN_15305; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15307 = 8'hcb == io_state_in_15 ? 8'h44 : _GEN_15306; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15308 = 8'hcc == io_state_in_15 ? 8'h75 : _GEN_15307; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15309 = 8'hcd == io_state_in_15 ? 8'h7e : _GEN_15308; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15310 = 8'hce == io_state_in_15 ? 8'h63 : _GEN_15309; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15311 = 8'hcf == io_state_in_15 ? 8'h68 : _GEN_15310; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15312 = 8'hd0 == io_state_in_15 ? 8'hb1 : _GEN_15311; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15313 = 8'hd1 == io_state_in_15 ? 8'hba : _GEN_15312; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15314 = 8'hd2 == io_state_in_15 ? 8'ha7 : _GEN_15313; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15315 = 8'hd3 == io_state_in_15 ? 8'hac : _GEN_15314; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15316 = 8'hd4 == io_state_in_15 ? 8'h9d : _GEN_15315; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15317 = 8'hd5 == io_state_in_15 ? 8'h96 : _GEN_15316; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15318 = 8'hd6 == io_state_in_15 ? 8'h8b : _GEN_15317; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15319 = 8'hd7 == io_state_in_15 ? 8'h80 : _GEN_15318; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15320 = 8'hd8 == io_state_in_15 ? 8'he9 : _GEN_15319; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15321 = 8'hd9 == io_state_in_15 ? 8'he2 : _GEN_15320; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15322 = 8'hda == io_state_in_15 ? 8'hff : _GEN_15321; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15323 = 8'hdb == io_state_in_15 ? 8'hf4 : _GEN_15322; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15324 = 8'hdc == io_state_in_15 ? 8'hc5 : _GEN_15323; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15325 = 8'hdd == io_state_in_15 ? 8'hce : _GEN_15324; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15326 = 8'hde == io_state_in_15 ? 8'hd3 : _GEN_15325; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15327 = 8'hdf == io_state_in_15 ? 8'hd8 : _GEN_15326; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15328 = 8'he0 == io_state_in_15 ? 8'h7a : _GEN_15327; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15329 = 8'he1 == io_state_in_15 ? 8'h71 : _GEN_15328; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15330 = 8'he2 == io_state_in_15 ? 8'h6c : _GEN_15329; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15331 = 8'he3 == io_state_in_15 ? 8'h67 : _GEN_15330; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15332 = 8'he4 == io_state_in_15 ? 8'h56 : _GEN_15331; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15333 = 8'he5 == io_state_in_15 ? 8'h5d : _GEN_15332; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15334 = 8'he6 == io_state_in_15 ? 8'h40 : _GEN_15333; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15335 = 8'he7 == io_state_in_15 ? 8'h4b : _GEN_15334; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15336 = 8'he8 == io_state_in_15 ? 8'h22 : _GEN_15335; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15337 = 8'he9 == io_state_in_15 ? 8'h29 : _GEN_15336; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15338 = 8'hea == io_state_in_15 ? 8'h34 : _GEN_15337; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15339 = 8'heb == io_state_in_15 ? 8'h3f : _GEN_15338; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15340 = 8'hec == io_state_in_15 ? 8'he : _GEN_15339; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15341 = 8'hed == io_state_in_15 ? 8'h5 : _GEN_15340; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15342 = 8'hee == io_state_in_15 ? 8'h18 : _GEN_15341; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15343 = 8'hef == io_state_in_15 ? 8'h13 : _GEN_15342; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15344 = 8'hf0 == io_state_in_15 ? 8'hca : _GEN_15343; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15345 = 8'hf1 == io_state_in_15 ? 8'hc1 : _GEN_15344; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15346 = 8'hf2 == io_state_in_15 ? 8'hdc : _GEN_15345; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15347 = 8'hf3 == io_state_in_15 ? 8'hd7 : _GEN_15346; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15348 = 8'hf4 == io_state_in_15 ? 8'he6 : _GEN_15347; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15349 = 8'hf5 == io_state_in_15 ? 8'hed : _GEN_15348; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15350 = 8'hf6 == io_state_in_15 ? 8'hf0 : _GEN_15349; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15351 = 8'hf7 == io_state_in_15 ? 8'hfb : _GEN_15350; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15352 = 8'hf8 == io_state_in_15 ? 8'h92 : _GEN_15351; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15353 = 8'hf9 == io_state_in_15 ? 8'h99 : _GEN_15352; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15354 = 8'hfa == io_state_in_15 ? 8'h84 : _GEN_15353; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15355 = 8'hfb == io_state_in_15 ? 8'h8f : _GEN_15354; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15356 = 8'hfc == io_state_in_15 ? 8'hbe : _GEN_15355; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15357 = 8'hfd == io_state_in_15 ? 8'hb5 : _GEN_15356; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15358 = 8'hfe == io_state_in_15 ? 8'ha8 : _GEN_15357; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15359 = 8'hff == io_state_in_15 ? 8'ha3 : _GEN_15358; // @[InvMixColumns.scala 143:{93,93}]
  wire [7:0] _GEN_15361 = 8'h1 == io_state_in_12 ? 8'hb : 8'h0; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15362 = 8'h2 == io_state_in_12 ? 8'h16 : _GEN_15361; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15363 = 8'h3 == io_state_in_12 ? 8'h1d : _GEN_15362; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15364 = 8'h4 == io_state_in_12 ? 8'h2c : _GEN_15363; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15365 = 8'h5 == io_state_in_12 ? 8'h27 : _GEN_15364; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15366 = 8'h6 == io_state_in_12 ? 8'h3a : _GEN_15365; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15367 = 8'h7 == io_state_in_12 ? 8'h31 : _GEN_15366; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15368 = 8'h8 == io_state_in_12 ? 8'h58 : _GEN_15367; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15369 = 8'h9 == io_state_in_12 ? 8'h53 : _GEN_15368; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15370 = 8'ha == io_state_in_12 ? 8'h4e : _GEN_15369; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15371 = 8'hb == io_state_in_12 ? 8'h45 : _GEN_15370; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15372 = 8'hc == io_state_in_12 ? 8'h74 : _GEN_15371; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15373 = 8'hd == io_state_in_12 ? 8'h7f : _GEN_15372; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15374 = 8'he == io_state_in_12 ? 8'h62 : _GEN_15373; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15375 = 8'hf == io_state_in_12 ? 8'h69 : _GEN_15374; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15376 = 8'h10 == io_state_in_12 ? 8'hb0 : _GEN_15375; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15377 = 8'h11 == io_state_in_12 ? 8'hbb : _GEN_15376; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15378 = 8'h12 == io_state_in_12 ? 8'ha6 : _GEN_15377; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15379 = 8'h13 == io_state_in_12 ? 8'had : _GEN_15378; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15380 = 8'h14 == io_state_in_12 ? 8'h9c : _GEN_15379; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15381 = 8'h15 == io_state_in_12 ? 8'h97 : _GEN_15380; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15382 = 8'h16 == io_state_in_12 ? 8'h8a : _GEN_15381; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15383 = 8'h17 == io_state_in_12 ? 8'h81 : _GEN_15382; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15384 = 8'h18 == io_state_in_12 ? 8'he8 : _GEN_15383; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15385 = 8'h19 == io_state_in_12 ? 8'he3 : _GEN_15384; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15386 = 8'h1a == io_state_in_12 ? 8'hfe : _GEN_15385; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15387 = 8'h1b == io_state_in_12 ? 8'hf5 : _GEN_15386; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15388 = 8'h1c == io_state_in_12 ? 8'hc4 : _GEN_15387; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15389 = 8'h1d == io_state_in_12 ? 8'hcf : _GEN_15388; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15390 = 8'h1e == io_state_in_12 ? 8'hd2 : _GEN_15389; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15391 = 8'h1f == io_state_in_12 ? 8'hd9 : _GEN_15390; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15392 = 8'h20 == io_state_in_12 ? 8'h7b : _GEN_15391; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15393 = 8'h21 == io_state_in_12 ? 8'h70 : _GEN_15392; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15394 = 8'h22 == io_state_in_12 ? 8'h6d : _GEN_15393; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15395 = 8'h23 == io_state_in_12 ? 8'h66 : _GEN_15394; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15396 = 8'h24 == io_state_in_12 ? 8'h57 : _GEN_15395; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15397 = 8'h25 == io_state_in_12 ? 8'h5c : _GEN_15396; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15398 = 8'h26 == io_state_in_12 ? 8'h41 : _GEN_15397; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15399 = 8'h27 == io_state_in_12 ? 8'h4a : _GEN_15398; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15400 = 8'h28 == io_state_in_12 ? 8'h23 : _GEN_15399; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15401 = 8'h29 == io_state_in_12 ? 8'h28 : _GEN_15400; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15402 = 8'h2a == io_state_in_12 ? 8'h35 : _GEN_15401; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15403 = 8'h2b == io_state_in_12 ? 8'h3e : _GEN_15402; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15404 = 8'h2c == io_state_in_12 ? 8'hf : _GEN_15403; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15405 = 8'h2d == io_state_in_12 ? 8'h4 : _GEN_15404; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15406 = 8'h2e == io_state_in_12 ? 8'h19 : _GEN_15405; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15407 = 8'h2f == io_state_in_12 ? 8'h12 : _GEN_15406; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15408 = 8'h30 == io_state_in_12 ? 8'hcb : _GEN_15407; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15409 = 8'h31 == io_state_in_12 ? 8'hc0 : _GEN_15408; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15410 = 8'h32 == io_state_in_12 ? 8'hdd : _GEN_15409; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15411 = 8'h33 == io_state_in_12 ? 8'hd6 : _GEN_15410; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15412 = 8'h34 == io_state_in_12 ? 8'he7 : _GEN_15411; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15413 = 8'h35 == io_state_in_12 ? 8'hec : _GEN_15412; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15414 = 8'h36 == io_state_in_12 ? 8'hf1 : _GEN_15413; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15415 = 8'h37 == io_state_in_12 ? 8'hfa : _GEN_15414; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15416 = 8'h38 == io_state_in_12 ? 8'h93 : _GEN_15415; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15417 = 8'h39 == io_state_in_12 ? 8'h98 : _GEN_15416; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15418 = 8'h3a == io_state_in_12 ? 8'h85 : _GEN_15417; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15419 = 8'h3b == io_state_in_12 ? 8'h8e : _GEN_15418; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15420 = 8'h3c == io_state_in_12 ? 8'hbf : _GEN_15419; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15421 = 8'h3d == io_state_in_12 ? 8'hb4 : _GEN_15420; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15422 = 8'h3e == io_state_in_12 ? 8'ha9 : _GEN_15421; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15423 = 8'h3f == io_state_in_12 ? 8'ha2 : _GEN_15422; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15424 = 8'h40 == io_state_in_12 ? 8'hf6 : _GEN_15423; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15425 = 8'h41 == io_state_in_12 ? 8'hfd : _GEN_15424; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15426 = 8'h42 == io_state_in_12 ? 8'he0 : _GEN_15425; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15427 = 8'h43 == io_state_in_12 ? 8'heb : _GEN_15426; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15428 = 8'h44 == io_state_in_12 ? 8'hda : _GEN_15427; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15429 = 8'h45 == io_state_in_12 ? 8'hd1 : _GEN_15428; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15430 = 8'h46 == io_state_in_12 ? 8'hcc : _GEN_15429; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15431 = 8'h47 == io_state_in_12 ? 8'hc7 : _GEN_15430; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15432 = 8'h48 == io_state_in_12 ? 8'hae : _GEN_15431; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15433 = 8'h49 == io_state_in_12 ? 8'ha5 : _GEN_15432; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15434 = 8'h4a == io_state_in_12 ? 8'hb8 : _GEN_15433; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15435 = 8'h4b == io_state_in_12 ? 8'hb3 : _GEN_15434; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15436 = 8'h4c == io_state_in_12 ? 8'h82 : _GEN_15435; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15437 = 8'h4d == io_state_in_12 ? 8'h89 : _GEN_15436; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15438 = 8'h4e == io_state_in_12 ? 8'h94 : _GEN_15437; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15439 = 8'h4f == io_state_in_12 ? 8'h9f : _GEN_15438; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15440 = 8'h50 == io_state_in_12 ? 8'h46 : _GEN_15439; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15441 = 8'h51 == io_state_in_12 ? 8'h4d : _GEN_15440; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15442 = 8'h52 == io_state_in_12 ? 8'h50 : _GEN_15441; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15443 = 8'h53 == io_state_in_12 ? 8'h5b : _GEN_15442; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15444 = 8'h54 == io_state_in_12 ? 8'h6a : _GEN_15443; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15445 = 8'h55 == io_state_in_12 ? 8'h61 : _GEN_15444; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15446 = 8'h56 == io_state_in_12 ? 8'h7c : _GEN_15445; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15447 = 8'h57 == io_state_in_12 ? 8'h77 : _GEN_15446; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15448 = 8'h58 == io_state_in_12 ? 8'h1e : _GEN_15447; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15449 = 8'h59 == io_state_in_12 ? 8'h15 : _GEN_15448; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15450 = 8'h5a == io_state_in_12 ? 8'h8 : _GEN_15449; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15451 = 8'h5b == io_state_in_12 ? 8'h3 : _GEN_15450; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15452 = 8'h5c == io_state_in_12 ? 8'h32 : _GEN_15451; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15453 = 8'h5d == io_state_in_12 ? 8'h39 : _GEN_15452; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15454 = 8'h5e == io_state_in_12 ? 8'h24 : _GEN_15453; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15455 = 8'h5f == io_state_in_12 ? 8'h2f : _GEN_15454; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15456 = 8'h60 == io_state_in_12 ? 8'h8d : _GEN_15455; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15457 = 8'h61 == io_state_in_12 ? 8'h86 : _GEN_15456; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15458 = 8'h62 == io_state_in_12 ? 8'h9b : _GEN_15457; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15459 = 8'h63 == io_state_in_12 ? 8'h90 : _GEN_15458; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15460 = 8'h64 == io_state_in_12 ? 8'ha1 : _GEN_15459; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15461 = 8'h65 == io_state_in_12 ? 8'haa : _GEN_15460; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15462 = 8'h66 == io_state_in_12 ? 8'hb7 : _GEN_15461; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15463 = 8'h67 == io_state_in_12 ? 8'hbc : _GEN_15462; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15464 = 8'h68 == io_state_in_12 ? 8'hd5 : _GEN_15463; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15465 = 8'h69 == io_state_in_12 ? 8'hde : _GEN_15464; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15466 = 8'h6a == io_state_in_12 ? 8'hc3 : _GEN_15465; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15467 = 8'h6b == io_state_in_12 ? 8'hc8 : _GEN_15466; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15468 = 8'h6c == io_state_in_12 ? 8'hf9 : _GEN_15467; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15469 = 8'h6d == io_state_in_12 ? 8'hf2 : _GEN_15468; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15470 = 8'h6e == io_state_in_12 ? 8'hef : _GEN_15469; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15471 = 8'h6f == io_state_in_12 ? 8'he4 : _GEN_15470; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15472 = 8'h70 == io_state_in_12 ? 8'h3d : _GEN_15471; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15473 = 8'h71 == io_state_in_12 ? 8'h36 : _GEN_15472; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15474 = 8'h72 == io_state_in_12 ? 8'h2b : _GEN_15473; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15475 = 8'h73 == io_state_in_12 ? 8'h20 : _GEN_15474; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15476 = 8'h74 == io_state_in_12 ? 8'h11 : _GEN_15475; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15477 = 8'h75 == io_state_in_12 ? 8'h1a : _GEN_15476; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15478 = 8'h76 == io_state_in_12 ? 8'h7 : _GEN_15477; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15479 = 8'h77 == io_state_in_12 ? 8'hc : _GEN_15478; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15480 = 8'h78 == io_state_in_12 ? 8'h65 : _GEN_15479; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15481 = 8'h79 == io_state_in_12 ? 8'h6e : _GEN_15480; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15482 = 8'h7a == io_state_in_12 ? 8'h73 : _GEN_15481; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15483 = 8'h7b == io_state_in_12 ? 8'h78 : _GEN_15482; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15484 = 8'h7c == io_state_in_12 ? 8'h49 : _GEN_15483; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15485 = 8'h7d == io_state_in_12 ? 8'h42 : _GEN_15484; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15486 = 8'h7e == io_state_in_12 ? 8'h5f : _GEN_15485; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15487 = 8'h7f == io_state_in_12 ? 8'h54 : _GEN_15486; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15488 = 8'h80 == io_state_in_12 ? 8'hf7 : _GEN_15487; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15489 = 8'h81 == io_state_in_12 ? 8'hfc : _GEN_15488; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15490 = 8'h82 == io_state_in_12 ? 8'he1 : _GEN_15489; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15491 = 8'h83 == io_state_in_12 ? 8'hea : _GEN_15490; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15492 = 8'h84 == io_state_in_12 ? 8'hdb : _GEN_15491; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15493 = 8'h85 == io_state_in_12 ? 8'hd0 : _GEN_15492; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15494 = 8'h86 == io_state_in_12 ? 8'hcd : _GEN_15493; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15495 = 8'h87 == io_state_in_12 ? 8'hc6 : _GEN_15494; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15496 = 8'h88 == io_state_in_12 ? 8'haf : _GEN_15495; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15497 = 8'h89 == io_state_in_12 ? 8'ha4 : _GEN_15496; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15498 = 8'h8a == io_state_in_12 ? 8'hb9 : _GEN_15497; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15499 = 8'h8b == io_state_in_12 ? 8'hb2 : _GEN_15498; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15500 = 8'h8c == io_state_in_12 ? 8'h83 : _GEN_15499; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15501 = 8'h8d == io_state_in_12 ? 8'h88 : _GEN_15500; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15502 = 8'h8e == io_state_in_12 ? 8'h95 : _GEN_15501; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15503 = 8'h8f == io_state_in_12 ? 8'h9e : _GEN_15502; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15504 = 8'h90 == io_state_in_12 ? 8'h47 : _GEN_15503; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15505 = 8'h91 == io_state_in_12 ? 8'h4c : _GEN_15504; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15506 = 8'h92 == io_state_in_12 ? 8'h51 : _GEN_15505; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15507 = 8'h93 == io_state_in_12 ? 8'h5a : _GEN_15506; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15508 = 8'h94 == io_state_in_12 ? 8'h6b : _GEN_15507; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15509 = 8'h95 == io_state_in_12 ? 8'h60 : _GEN_15508; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15510 = 8'h96 == io_state_in_12 ? 8'h7d : _GEN_15509; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15511 = 8'h97 == io_state_in_12 ? 8'h76 : _GEN_15510; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15512 = 8'h98 == io_state_in_12 ? 8'h1f : _GEN_15511; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15513 = 8'h99 == io_state_in_12 ? 8'h14 : _GEN_15512; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15514 = 8'h9a == io_state_in_12 ? 8'h9 : _GEN_15513; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15515 = 8'h9b == io_state_in_12 ? 8'h2 : _GEN_15514; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15516 = 8'h9c == io_state_in_12 ? 8'h33 : _GEN_15515; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15517 = 8'h9d == io_state_in_12 ? 8'h38 : _GEN_15516; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15518 = 8'h9e == io_state_in_12 ? 8'h25 : _GEN_15517; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15519 = 8'h9f == io_state_in_12 ? 8'h2e : _GEN_15518; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15520 = 8'ha0 == io_state_in_12 ? 8'h8c : _GEN_15519; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15521 = 8'ha1 == io_state_in_12 ? 8'h87 : _GEN_15520; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15522 = 8'ha2 == io_state_in_12 ? 8'h9a : _GEN_15521; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15523 = 8'ha3 == io_state_in_12 ? 8'h91 : _GEN_15522; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15524 = 8'ha4 == io_state_in_12 ? 8'ha0 : _GEN_15523; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15525 = 8'ha5 == io_state_in_12 ? 8'hab : _GEN_15524; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15526 = 8'ha6 == io_state_in_12 ? 8'hb6 : _GEN_15525; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15527 = 8'ha7 == io_state_in_12 ? 8'hbd : _GEN_15526; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15528 = 8'ha8 == io_state_in_12 ? 8'hd4 : _GEN_15527; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15529 = 8'ha9 == io_state_in_12 ? 8'hdf : _GEN_15528; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15530 = 8'haa == io_state_in_12 ? 8'hc2 : _GEN_15529; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15531 = 8'hab == io_state_in_12 ? 8'hc9 : _GEN_15530; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15532 = 8'hac == io_state_in_12 ? 8'hf8 : _GEN_15531; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15533 = 8'had == io_state_in_12 ? 8'hf3 : _GEN_15532; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15534 = 8'hae == io_state_in_12 ? 8'hee : _GEN_15533; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15535 = 8'haf == io_state_in_12 ? 8'he5 : _GEN_15534; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15536 = 8'hb0 == io_state_in_12 ? 8'h3c : _GEN_15535; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15537 = 8'hb1 == io_state_in_12 ? 8'h37 : _GEN_15536; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15538 = 8'hb2 == io_state_in_12 ? 8'h2a : _GEN_15537; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15539 = 8'hb3 == io_state_in_12 ? 8'h21 : _GEN_15538; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15540 = 8'hb4 == io_state_in_12 ? 8'h10 : _GEN_15539; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15541 = 8'hb5 == io_state_in_12 ? 8'h1b : _GEN_15540; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15542 = 8'hb6 == io_state_in_12 ? 8'h6 : _GEN_15541; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15543 = 8'hb7 == io_state_in_12 ? 8'hd : _GEN_15542; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15544 = 8'hb8 == io_state_in_12 ? 8'h64 : _GEN_15543; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15545 = 8'hb9 == io_state_in_12 ? 8'h6f : _GEN_15544; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15546 = 8'hba == io_state_in_12 ? 8'h72 : _GEN_15545; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15547 = 8'hbb == io_state_in_12 ? 8'h79 : _GEN_15546; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15548 = 8'hbc == io_state_in_12 ? 8'h48 : _GEN_15547; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15549 = 8'hbd == io_state_in_12 ? 8'h43 : _GEN_15548; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15550 = 8'hbe == io_state_in_12 ? 8'h5e : _GEN_15549; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15551 = 8'hbf == io_state_in_12 ? 8'h55 : _GEN_15550; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15552 = 8'hc0 == io_state_in_12 ? 8'h1 : _GEN_15551; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15553 = 8'hc1 == io_state_in_12 ? 8'ha : _GEN_15552; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15554 = 8'hc2 == io_state_in_12 ? 8'h17 : _GEN_15553; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15555 = 8'hc3 == io_state_in_12 ? 8'h1c : _GEN_15554; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15556 = 8'hc4 == io_state_in_12 ? 8'h2d : _GEN_15555; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15557 = 8'hc5 == io_state_in_12 ? 8'h26 : _GEN_15556; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15558 = 8'hc6 == io_state_in_12 ? 8'h3b : _GEN_15557; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15559 = 8'hc7 == io_state_in_12 ? 8'h30 : _GEN_15558; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15560 = 8'hc8 == io_state_in_12 ? 8'h59 : _GEN_15559; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15561 = 8'hc9 == io_state_in_12 ? 8'h52 : _GEN_15560; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15562 = 8'hca == io_state_in_12 ? 8'h4f : _GEN_15561; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15563 = 8'hcb == io_state_in_12 ? 8'h44 : _GEN_15562; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15564 = 8'hcc == io_state_in_12 ? 8'h75 : _GEN_15563; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15565 = 8'hcd == io_state_in_12 ? 8'h7e : _GEN_15564; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15566 = 8'hce == io_state_in_12 ? 8'h63 : _GEN_15565; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15567 = 8'hcf == io_state_in_12 ? 8'h68 : _GEN_15566; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15568 = 8'hd0 == io_state_in_12 ? 8'hb1 : _GEN_15567; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15569 = 8'hd1 == io_state_in_12 ? 8'hba : _GEN_15568; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15570 = 8'hd2 == io_state_in_12 ? 8'ha7 : _GEN_15569; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15571 = 8'hd3 == io_state_in_12 ? 8'hac : _GEN_15570; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15572 = 8'hd4 == io_state_in_12 ? 8'h9d : _GEN_15571; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15573 = 8'hd5 == io_state_in_12 ? 8'h96 : _GEN_15572; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15574 = 8'hd6 == io_state_in_12 ? 8'h8b : _GEN_15573; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15575 = 8'hd7 == io_state_in_12 ? 8'h80 : _GEN_15574; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15576 = 8'hd8 == io_state_in_12 ? 8'he9 : _GEN_15575; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15577 = 8'hd9 == io_state_in_12 ? 8'he2 : _GEN_15576; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15578 = 8'hda == io_state_in_12 ? 8'hff : _GEN_15577; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15579 = 8'hdb == io_state_in_12 ? 8'hf4 : _GEN_15578; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15580 = 8'hdc == io_state_in_12 ? 8'hc5 : _GEN_15579; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15581 = 8'hdd == io_state_in_12 ? 8'hce : _GEN_15580; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15582 = 8'hde == io_state_in_12 ? 8'hd3 : _GEN_15581; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15583 = 8'hdf == io_state_in_12 ? 8'hd8 : _GEN_15582; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15584 = 8'he0 == io_state_in_12 ? 8'h7a : _GEN_15583; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15585 = 8'he1 == io_state_in_12 ? 8'h71 : _GEN_15584; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15586 = 8'he2 == io_state_in_12 ? 8'h6c : _GEN_15585; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15587 = 8'he3 == io_state_in_12 ? 8'h67 : _GEN_15586; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15588 = 8'he4 == io_state_in_12 ? 8'h56 : _GEN_15587; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15589 = 8'he5 == io_state_in_12 ? 8'h5d : _GEN_15588; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15590 = 8'he6 == io_state_in_12 ? 8'h40 : _GEN_15589; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15591 = 8'he7 == io_state_in_12 ? 8'h4b : _GEN_15590; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15592 = 8'he8 == io_state_in_12 ? 8'h22 : _GEN_15591; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15593 = 8'he9 == io_state_in_12 ? 8'h29 : _GEN_15592; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15594 = 8'hea == io_state_in_12 ? 8'h34 : _GEN_15593; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15595 = 8'heb == io_state_in_12 ? 8'h3f : _GEN_15594; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15596 = 8'hec == io_state_in_12 ? 8'he : _GEN_15595; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15597 = 8'hed == io_state_in_12 ? 8'h5 : _GEN_15596; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15598 = 8'hee == io_state_in_12 ? 8'h18 : _GEN_15597; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15599 = 8'hef == io_state_in_12 ? 8'h13 : _GEN_15598; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15600 = 8'hf0 == io_state_in_12 ? 8'hca : _GEN_15599; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15601 = 8'hf1 == io_state_in_12 ? 8'hc1 : _GEN_15600; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15602 = 8'hf2 == io_state_in_12 ? 8'hdc : _GEN_15601; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15603 = 8'hf3 == io_state_in_12 ? 8'hd7 : _GEN_15602; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15604 = 8'hf4 == io_state_in_12 ? 8'he6 : _GEN_15603; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15605 = 8'hf5 == io_state_in_12 ? 8'hed : _GEN_15604; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15606 = 8'hf6 == io_state_in_12 ? 8'hf0 : _GEN_15605; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15607 = 8'hf7 == io_state_in_12 ? 8'hfb : _GEN_15606; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15608 = 8'hf8 == io_state_in_12 ? 8'h92 : _GEN_15607; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15609 = 8'hf9 == io_state_in_12 ? 8'h99 : _GEN_15608; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15610 = 8'hfa == io_state_in_12 ? 8'h84 : _GEN_15609; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15611 = 8'hfb == io_state_in_12 ? 8'h8f : _GEN_15610; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15612 = 8'hfc == io_state_in_12 ? 8'hbe : _GEN_15611; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15613 = 8'hfd == io_state_in_12 ? 8'hb5 : _GEN_15612; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15614 = 8'hfe == io_state_in_12 ? 8'ha8 : _GEN_15613; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15615 = 8'hff == io_state_in_12 ? 8'ha3 : _GEN_15614; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15617 = 8'h1 == io_state_in_13 ? 8'hd : 8'h0; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15618 = 8'h2 == io_state_in_13 ? 8'h1a : _GEN_15617; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15619 = 8'h3 == io_state_in_13 ? 8'h17 : _GEN_15618; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15620 = 8'h4 == io_state_in_13 ? 8'h34 : _GEN_15619; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15621 = 8'h5 == io_state_in_13 ? 8'h39 : _GEN_15620; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15622 = 8'h6 == io_state_in_13 ? 8'h2e : _GEN_15621; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15623 = 8'h7 == io_state_in_13 ? 8'h23 : _GEN_15622; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15624 = 8'h8 == io_state_in_13 ? 8'h68 : _GEN_15623; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15625 = 8'h9 == io_state_in_13 ? 8'h65 : _GEN_15624; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15626 = 8'ha == io_state_in_13 ? 8'h72 : _GEN_15625; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15627 = 8'hb == io_state_in_13 ? 8'h7f : _GEN_15626; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15628 = 8'hc == io_state_in_13 ? 8'h5c : _GEN_15627; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15629 = 8'hd == io_state_in_13 ? 8'h51 : _GEN_15628; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15630 = 8'he == io_state_in_13 ? 8'h46 : _GEN_15629; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15631 = 8'hf == io_state_in_13 ? 8'h4b : _GEN_15630; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15632 = 8'h10 == io_state_in_13 ? 8'hd0 : _GEN_15631; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15633 = 8'h11 == io_state_in_13 ? 8'hdd : _GEN_15632; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15634 = 8'h12 == io_state_in_13 ? 8'hca : _GEN_15633; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15635 = 8'h13 == io_state_in_13 ? 8'hc7 : _GEN_15634; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15636 = 8'h14 == io_state_in_13 ? 8'he4 : _GEN_15635; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15637 = 8'h15 == io_state_in_13 ? 8'he9 : _GEN_15636; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15638 = 8'h16 == io_state_in_13 ? 8'hfe : _GEN_15637; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15639 = 8'h17 == io_state_in_13 ? 8'hf3 : _GEN_15638; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15640 = 8'h18 == io_state_in_13 ? 8'hb8 : _GEN_15639; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15641 = 8'h19 == io_state_in_13 ? 8'hb5 : _GEN_15640; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15642 = 8'h1a == io_state_in_13 ? 8'ha2 : _GEN_15641; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15643 = 8'h1b == io_state_in_13 ? 8'haf : _GEN_15642; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15644 = 8'h1c == io_state_in_13 ? 8'h8c : _GEN_15643; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15645 = 8'h1d == io_state_in_13 ? 8'h81 : _GEN_15644; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15646 = 8'h1e == io_state_in_13 ? 8'h96 : _GEN_15645; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15647 = 8'h1f == io_state_in_13 ? 8'h9b : _GEN_15646; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15648 = 8'h20 == io_state_in_13 ? 8'hbb : _GEN_15647; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15649 = 8'h21 == io_state_in_13 ? 8'hb6 : _GEN_15648; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15650 = 8'h22 == io_state_in_13 ? 8'ha1 : _GEN_15649; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15651 = 8'h23 == io_state_in_13 ? 8'hac : _GEN_15650; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15652 = 8'h24 == io_state_in_13 ? 8'h8f : _GEN_15651; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15653 = 8'h25 == io_state_in_13 ? 8'h82 : _GEN_15652; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15654 = 8'h26 == io_state_in_13 ? 8'h95 : _GEN_15653; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15655 = 8'h27 == io_state_in_13 ? 8'h98 : _GEN_15654; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15656 = 8'h28 == io_state_in_13 ? 8'hd3 : _GEN_15655; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15657 = 8'h29 == io_state_in_13 ? 8'hde : _GEN_15656; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15658 = 8'h2a == io_state_in_13 ? 8'hc9 : _GEN_15657; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15659 = 8'h2b == io_state_in_13 ? 8'hc4 : _GEN_15658; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15660 = 8'h2c == io_state_in_13 ? 8'he7 : _GEN_15659; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15661 = 8'h2d == io_state_in_13 ? 8'hea : _GEN_15660; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15662 = 8'h2e == io_state_in_13 ? 8'hfd : _GEN_15661; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15663 = 8'h2f == io_state_in_13 ? 8'hf0 : _GEN_15662; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15664 = 8'h30 == io_state_in_13 ? 8'h6b : _GEN_15663; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15665 = 8'h31 == io_state_in_13 ? 8'h66 : _GEN_15664; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15666 = 8'h32 == io_state_in_13 ? 8'h71 : _GEN_15665; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15667 = 8'h33 == io_state_in_13 ? 8'h7c : _GEN_15666; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15668 = 8'h34 == io_state_in_13 ? 8'h5f : _GEN_15667; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15669 = 8'h35 == io_state_in_13 ? 8'h52 : _GEN_15668; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15670 = 8'h36 == io_state_in_13 ? 8'h45 : _GEN_15669; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15671 = 8'h37 == io_state_in_13 ? 8'h48 : _GEN_15670; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15672 = 8'h38 == io_state_in_13 ? 8'h3 : _GEN_15671; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15673 = 8'h39 == io_state_in_13 ? 8'he : _GEN_15672; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15674 = 8'h3a == io_state_in_13 ? 8'h19 : _GEN_15673; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15675 = 8'h3b == io_state_in_13 ? 8'h14 : _GEN_15674; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15676 = 8'h3c == io_state_in_13 ? 8'h37 : _GEN_15675; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15677 = 8'h3d == io_state_in_13 ? 8'h3a : _GEN_15676; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15678 = 8'h3e == io_state_in_13 ? 8'h2d : _GEN_15677; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15679 = 8'h3f == io_state_in_13 ? 8'h20 : _GEN_15678; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15680 = 8'h40 == io_state_in_13 ? 8'h6d : _GEN_15679; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15681 = 8'h41 == io_state_in_13 ? 8'h60 : _GEN_15680; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15682 = 8'h42 == io_state_in_13 ? 8'h77 : _GEN_15681; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15683 = 8'h43 == io_state_in_13 ? 8'h7a : _GEN_15682; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15684 = 8'h44 == io_state_in_13 ? 8'h59 : _GEN_15683; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15685 = 8'h45 == io_state_in_13 ? 8'h54 : _GEN_15684; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15686 = 8'h46 == io_state_in_13 ? 8'h43 : _GEN_15685; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15687 = 8'h47 == io_state_in_13 ? 8'h4e : _GEN_15686; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15688 = 8'h48 == io_state_in_13 ? 8'h5 : _GEN_15687; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15689 = 8'h49 == io_state_in_13 ? 8'h8 : _GEN_15688; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15690 = 8'h4a == io_state_in_13 ? 8'h1f : _GEN_15689; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15691 = 8'h4b == io_state_in_13 ? 8'h12 : _GEN_15690; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15692 = 8'h4c == io_state_in_13 ? 8'h31 : _GEN_15691; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15693 = 8'h4d == io_state_in_13 ? 8'h3c : _GEN_15692; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15694 = 8'h4e == io_state_in_13 ? 8'h2b : _GEN_15693; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15695 = 8'h4f == io_state_in_13 ? 8'h26 : _GEN_15694; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15696 = 8'h50 == io_state_in_13 ? 8'hbd : _GEN_15695; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15697 = 8'h51 == io_state_in_13 ? 8'hb0 : _GEN_15696; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15698 = 8'h52 == io_state_in_13 ? 8'ha7 : _GEN_15697; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15699 = 8'h53 == io_state_in_13 ? 8'haa : _GEN_15698; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15700 = 8'h54 == io_state_in_13 ? 8'h89 : _GEN_15699; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15701 = 8'h55 == io_state_in_13 ? 8'h84 : _GEN_15700; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15702 = 8'h56 == io_state_in_13 ? 8'h93 : _GEN_15701; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15703 = 8'h57 == io_state_in_13 ? 8'h9e : _GEN_15702; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15704 = 8'h58 == io_state_in_13 ? 8'hd5 : _GEN_15703; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15705 = 8'h59 == io_state_in_13 ? 8'hd8 : _GEN_15704; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15706 = 8'h5a == io_state_in_13 ? 8'hcf : _GEN_15705; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15707 = 8'h5b == io_state_in_13 ? 8'hc2 : _GEN_15706; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15708 = 8'h5c == io_state_in_13 ? 8'he1 : _GEN_15707; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15709 = 8'h5d == io_state_in_13 ? 8'hec : _GEN_15708; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15710 = 8'h5e == io_state_in_13 ? 8'hfb : _GEN_15709; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15711 = 8'h5f == io_state_in_13 ? 8'hf6 : _GEN_15710; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15712 = 8'h60 == io_state_in_13 ? 8'hd6 : _GEN_15711; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15713 = 8'h61 == io_state_in_13 ? 8'hdb : _GEN_15712; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15714 = 8'h62 == io_state_in_13 ? 8'hcc : _GEN_15713; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15715 = 8'h63 == io_state_in_13 ? 8'hc1 : _GEN_15714; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15716 = 8'h64 == io_state_in_13 ? 8'he2 : _GEN_15715; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15717 = 8'h65 == io_state_in_13 ? 8'hef : _GEN_15716; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15718 = 8'h66 == io_state_in_13 ? 8'hf8 : _GEN_15717; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15719 = 8'h67 == io_state_in_13 ? 8'hf5 : _GEN_15718; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15720 = 8'h68 == io_state_in_13 ? 8'hbe : _GEN_15719; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15721 = 8'h69 == io_state_in_13 ? 8'hb3 : _GEN_15720; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15722 = 8'h6a == io_state_in_13 ? 8'ha4 : _GEN_15721; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15723 = 8'h6b == io_state_in_13 ? 8'ha9 : _GEN_15722; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15724 = 8'h6c == io_state_in_13 ? 8'h8a : _GEN_15723; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15725 = 8'h6d == io_state_in_13 ? 8'h87 : _GEN_15724; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15726 = 8'h6e == io_state_in_13 ? 8'h90 : _GEN_15725; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15727 = 8'h6f == io_state_in_13 ? 8'h9d : _GEN_15726; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15728 = 8'h70 == io_state_in_13 ? 8'h6 : _GEN_15727; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15729 = 8'h71 == io_state_in_13 ? 8'hb : _GEN_15728; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15730 = 8'h72 == io_state_in_13 ? 8'h1c : _GEN_15729; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15731 = 8'h73 == io_state_in_13 ? 8'h11 : _GEN_15730; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15732 = 8'h74 == io_state_in_13 ? 8'h32 : _GEN_15731; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15733 = 8'h75 == io_state_in_13 ? 8'h3f : _GEN_15732; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15734 = 8'h76 == io_state_in_13 ? 8'h28 : _GEN_15733; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15735 = 8'h77 == io_state_in_13 ? 8'h25 : _GEN_15734; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15736 = 8'h78 == io_state_in_13 ? 8'h6e : _GEN_15735; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15737 = 8'h79 == io_state_in_13 ? 8'h63 : _GEN_15736; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15738 = 8'h7a == io_state_in_13 ? 8'h74 : _GEN_15737; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15739 = 8'h7b == io_state_in_13 ? 8'h79 : _GEN_15738; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15740 = 8'h7c == io_state_in_13 ? 8'h5a : _GEN_15739; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15741 = 8'h7d == io_state_in_13 ? 8'h57 : _GEN_15740; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15742 = 8'h7e == io_state_in_13 ? 8'h40 : _GEN_15741; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15743 = 8'h7f == io_state_in_13 ? 8'h4d : _GEN_15742; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15744 = 8'h80 == io_state_in_13 ? 8'hda : _GEN_15743; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15745 = 8'h81 == io_state_in_13 ? 8'hd7 : _GEN_15744; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15746 = 8'h82 == io_state_in_13 ? 8'hc0 : _GEN_15745; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15747 = 8'h83 == io_state_in_13 ? 8'hcd : _GEN_15746; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15748 = 8'h84 == io_state_in_13 ? 8'hee : _GEN_15747; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15749 = 8'h85 == io_state_in_13 ? 8'he3 : _GEN_15748; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15750 = 8'h86 == io_state_in_13 ? 8'hf4 : _GEN_15749; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15751 = 8'h87 == io_state_in_13 ? 8'hf9 : _GEN_15750; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15752 = 8'h88 == io_state_in_13 ? 8'hb2 : _GEN_15751; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15753 = 8'h89 == io_state_in_13 ? 8'hbf : _GEN_15752; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15754 = 8'h8a == io_state_in_13 ? 8'ha8 : _GEN_15753; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15755 = 8'h8b == io_state_in_13 ? 8'ha5 : _GEN_15754; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15756 = 8'h8c == io_state_in_13 ? 8'h86 : _GEN_15755; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15757 = 8'h8d == io_state_in_13 ? 8'h8b : _GEN_15756; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15758 = 8'h8e == io_state_in_13 ? 8'h9c : _GEN_15757; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15759 = 8'h8f == io_state_in_13 ? 8'h91 : _GEN_15758; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15760 = 8'h90 == io_state_in_13 ? 8'ha : _GEN_15759; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15761 = 8'h91 == io_state_in_13 ? 8'h7 : _GEN_15760; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15762 = 8'h92 == io_state_in_13 ? 8'h10 : _GEN_15761; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15763 = 8'h93 == io_state_in_13 ? 8'h1d : _GEN_15762; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15764 = 8'h94 == io_state_in_13 ? 8'h3e : _GEN_15763; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15765 = 8'h95 == io_state_in_13 ? 8'h33 : _GEN_15764; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15766 = 8'h96 == io_state_in_13 ? 8'h24 : _GEN_15765; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15767 = 8'h97 == io_state_in_13 ? 8'h29 : _GEN_15766; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15768 = 8'h98 == io_state_in_13 ? 8'h62 : _GEN_15767; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15769 = 8'h99 == io_state_in_13 ? 8'h6f : _GEN_15768; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15770 = 8'h9a == io_state_in_13 ? 8'h78 : _GEN_15769; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15771 = 8'h9b == io_state_in_13 ? 8'h75 : _GEN_15770; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15772 = 8'h9c == io_state_in_13 ? 8'h56 : _GEN_15771; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15773 = 8'h9d == io_state_in_13 ? 8'h5b : _GEN_15772; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15774 = 8'h9e == io_state_in_13 ? 8'h4c : _GEN_15773; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15775 = 8'h9f == io_state_in_13 ? 8'h41 : _GEN_15774; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15776 = 8'ha0 == io_state_in_13 ? 8'h61 : _GEN_15775; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15777 = 8'ha1 == io_state_in_13 ? 8'h6c : _GEN_15776; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15778 = 8'ha2 == io_state_in_13 ? 8'h7b : _GEN_15777; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15779 = 8'ha3 == io_state_in_13 ? 8'h76 : _GEN_15778; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15780 = 8'ha4 == io_state_in_13 ? 8'h55 : _GEN_15779; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15781 = 8'ha5 == io_state_in_13 ? 8'h58 : _GEN_15780; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15782 = 8'ha6 == io_state_in_13 ? 8'h4f : _GEN_15781; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15783 = 8'ha7 == io_state_in_13 ? 8'h42 : _GEN_15782; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15784 = 8'ha8 == io_state_in_13 ? 8'h9 : _GEN_15783; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15785 = 8'ha9 == io_state_in_13 ? 8'h4 : _GEN_15784; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15786 = 8'haa == io_state_in_13 ? 8'h13 : _GEN_15785; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15787 = 8'hab == io_state_in_13 ? 8'h1e : _GEN_15786; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15788 = 8'hac == io_state_in_13 ? 8'h3d : _GEN_15787; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15789 = 8'had == io_state_in_13 ? 8'h30 : _GEN_15788; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15790 = 8'hae == io_state_in_13 ? 8'h27 : _GEN_15789; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15791 = 8'haf == io_state_in_13 ? 8'h2a : _GEN_15790; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15792 = 8'hb0 == io_state_in_13 ? 8'hb1 : _GEN_15791; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15793 = 8'hb1 == io_state_in_13 ? 8'hbc : _GEN_15792; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15794 = 8'hb2 == io_state_in_13 ? 8'hab : _GEN_15793; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15795 = 8'hb3 == io_state_in_13 ? 8'ha6 : _GEN_15794; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15796 = 8'hb4 == io_state_in_13 ? 8'h85 : _GEN_15795; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15797 = 8'hb5 == io_state_in_13 ? 8'h88 : _GEN_15796; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15798 = 8'hb6 == io_state_in_13 ? 8'h9f : _GEN_15797; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15799 = 8'hb7 == io_state_in_13 ? 8'h92 : _GEN_15798; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15800 = 8'hb8 == io_state_in_13 ? 8'hd9 : _GEN_15799; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15801 = 8'hb9 == io_state_in_13 ? 8'hd4 : _GEN_15800; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15802 = 8'hba == io_state_in_13 ? 8'hc3 : _GEN_15801; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15803 = 8'hbb == io_state_in_13 ? 8'hce : _GEN_15802; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15804 = 8'hbc == io_state_in_13 ? 8'hed : _GEN_15803; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15805 = 8'hbd == io_state_in_13 ? 8'he0 : _GEN_15804; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15806 = 8'hbe == io_state_in_13 ? 8'hf7 : _GEN_15805; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15807 = 8'hbf == io_state_in_13 ? 8'hfa : _GEN_15806; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15808 = 8'hc0 == io_state_in_13 ? 8'hb7 : _GEN_15807; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15809 = 8'hc1 == io_state_in_13 ? 8'hba : _GEN_15808; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15810 = 8'hc2 == io_state_in_13 ? 8'had : _GEN_15809; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15811 = 8'hc3 == io_state_in_13 ? 8'ha0 : _GEN_15810; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15812 = 8'hc4 == io_state_in_13 ? 8'h83 : _GEN_15811; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15813 = 8'hc5 == io_state_in_13 ? 8'h8e : _GEN_15812; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15814 = 8'hc6 == io_state_in_13 ? 8'h99 : _GEN_15813; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15815 = 8'hc7 == io_state_in_13 ? 8'h94 : _GEN_15814; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15816 = 8'hc8 == io_state_in_13 ? 8'hdf : _GEN_15815; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15817 = 8'hc9 == io_state_in_13 ? 8'hd2 : _GEN_15816; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15818 = 8'hca == io_state_in_13 ? 8'hc5 : _GEN_15817; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15819 = 8'hcb == io_state_in_13 ? 8'hc8 : _GEN_15818; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15820 = 8'hcc == io_state_in_13 ? 8'heb : _GEN_15819; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15821 = 8'hcd == io_state_in_13 ? 8'he6 : _GEN_15820; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15822 = 8'hce == io_state_in_13 ? 8'hf1 : _GEN_15821; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15823 = 8'hcf == io_state_in_13 ? 8'hfc : _GEN_15822; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15824 = 8'hd0 == io_state_in_13 ? 8'h67 : _GEN_15823; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15825 = 8'hd1 == io_state_in_13 ? 8'h6a : _GEN_15824; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15826 = 8'hd2 == io_state_in_13 ? 8'h7d : _GEN_15825; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15827 = 8'hd3 == io_state_in_13 ? 8'h70 : _GEN_15826; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15828 = 8'hd4 == io_state_in_13 ? 8'h53 : _GEN_15827; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15829 = 8'hd5 == io_state_in_13 ? 8'h5e : _GEN_15828; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15830 = 8'hd6 == io_state_in_13 ? 8'h49 : _GEN_15829; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15831 = 8'hd7 == io_state_in_13 ? 8'h44 : _GEN_15830; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15832 = 8'hd8 == io_state_in_13 ? 8'hf : _GEN_15831; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15833 = 8'hd9 == io_state_in_13 ? 8'h2 : _GEN_15832; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15834 = 8'hda == io_state_in_13 ? 8'h15 : _GEN_15833; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15835 = 8'hdb == io_state_in_13 ? 8'h18 : _GEN_15834; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15836 = 8'hdc == io_state_in_13 ? 8'h3b : _GEN_15835; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15837 = 8'hdd == io_state_in_13 ? 8'h36 : _GEN_15836; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15838 = 8'hde == io_state_in_13 ? 8'h21 : _GEN_15837; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15839 = 8'hdf == io_state_in_13 ? 8'h2c : _GEN_15838; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15840 = 8'he0 == io_state_in_13 ? 8'hc : _GEN_15839; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15841 = 8'he1 == io_state_in_13 ? 8'h1 : _GEN_15840; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15842 = 8'he2 == io_state_in_13 ? 8'h16 : _GEN_15841; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15843 = 8'he3 == io_state_in_13 ? 8'h1b : _GEN_15842; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15844 = 8'he4 == io_state_in_13 ? 8'h38 : _GEN_15843; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15845 = 8'he5 == io_state_in_13 ? 8'h35 : _GEN_15844; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15846 = 8'he6 == io_state_in_13 ? 8'h22 : _GEN_15845; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15847 = 8'he7 == io_state_in_13 ? 8'h2f : _GEN_15846; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15848 = 8'he8 == io_state_in_13 ? 8'h64 : _GEN_15847; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15849 = 8'he9 == io_state_in_13 ? 8'h69 : _GEN_15848; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15850 = 8'hea == io_state_in_13 ? 8'h7e : _GEN_15849; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15851 = 8'heb == io_state_in_13 ? 8'h73 : _GEN_15850; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15852 = 8'hec == io_state_in_13 ? 8'h50 : _GEN_15851; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15853 = 8'hed == io_state_in_13 ? 8'h5d : _GEN_15852; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15854 = 8'hee == io_state_in_13 ? 8'h4a : _GEN_15853; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15855 = 8'hef == io_state_in_13 ? 8'h47 : _GEN_15854; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15856 = 8'hf0 == io_state_in_13 ? 8'hdc : _GEN_15855; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15857 = 8'hf1 == io_state_in_13 ? 8'hd1 : _GEN_15856; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15858 = 8'hf2 == io_state_in_13 ? 8'hc6 : _GEN_15857; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15859 = 8'hf3 == io_state_in_13 ? 8'hcb : _GEN_15858; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15860 = 8'hf4 == io_state_in_13 ? 8'he8 : _GEN_15859; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15861 = 8'hf5 == io_state_in_13 ? 8'he5 : _GEN_15860; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15862 = 8'hf6 == io_state_in_13 ? 8'hf2 : _GEN_15861; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15863 = 8'hf7 == io_state_in_13 ? 8'hff : _GEN_15862; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15864 = 8'hf8 == io_state_in_13 ? 8'hb4 : _GEN_15863; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15865 = 8'hf9 == io_state_in_13 ? 8'hb9 : _GEN_15864; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15866 = 8'hfa == io_state_in_13 ? 8'hae : _GEN_15865; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15867 = 8'hfb == io_state_in_13 ? 8'ha3 : _GEN_15866; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15868 = 8'hfc == io_state_in_13 ? 8'h80 : _GEN_15867; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15869 = 8'hfd == io_state_in_13 ? 8'h8d : _GEN_15868; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15870 = 8'hfe == io_state_in_13 ? 8'h9a : _GEN_15869; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _GEN_15871 = 8'hff == io_state_in_13 ? 8'h97 : _GEN_15870; // @[InvMixColumns.scala 144:{43,43}]
  wire [7:0] _tmp_state_15_T = _GEN_15615 ^ _GEN_15871; // @[InvMixColumns.scala 144:43]
  wire [7:0] _GEN_15873 = 8'h1 == io_state_in_14 ? 8'h9 : 8'h0; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15874 = 8'h2 == io_state_in_14 ? 8'h12 : _GEN_15873; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15875 = 8'h3 == io_state_in_14 ? 8'h1b : _GEN_15874; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15876 = 8'h4 == io_state_in_14 ? 8'h24 : _GEN_15875; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15877 = 8'h5 == io_state_in_14 ? 8'h2d : _GEN_15876; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15878 = 8'h6 == io_state_in_14 ? 8'h36 : _GEN_15877; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15879 = 8'h7 == io_state_in_14 ? 8'h3f : _GEN_15878; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15880 = 8'h8 == io_state_in_14 ? 8'h48 : _GEN_15879; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15881 = 8'h9 == io_state_in_14 ? 8'h41 : _GEN_15880; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15882 = 8'ha == io_state_in_14 ? 8'h5a : _GEN_15881; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15883 = 8'hb == io_state_in_14 ? 8'h53 : _GEN_15882; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15884 = 8'hc == io_state_in_14 ? 8'h6c : _GEN_15883; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15885 = 8'hd == io_state_in_14 ? 8'h65 : _GEN_15884; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15886 = 8'he == io_state_in_14 ? 8'h7e : _GEN_15885; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15887 = 8'hf == io_state_in_14 ? 8'h77 : _GEN_15886; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15888 = 8'h10 == io_state_in_14 ? 8'h90 : _GEN_15887; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15889 = 8'h11 == io_state_in_14 ? 8'h99 : _GEN_15888; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15890 = 8'h12 == io_state_in_14 ? 8'h82 : _GEN_15889; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15891 = 8'h13 == io_state_in_14 ? 8'h8b : _GEN_15890; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15892 = 8'h14 == io_state_in_14 ? 8'hb4 : _GEN_15891; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15893 = 8'h15 == io_state_in_14 ? 8'hbd : _GEN_15892; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15894 = 8'h16 == io_state_in_14 ? 8'ha6 : _GEN_15893; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15895 = 8'h17 == io_state_in_14 ? 8'haf : _GEN_15894; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15896 = 8'h18 == io_state_in_14 ? 8'hd8 : _GEN_15895; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15897 = 8'h19 == io_state_in_14 ? 8'hd1 : _GEN_15896; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15898 = 8'h1a == io_state_in_14 ? 8'hca : _GEN_15897; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15899 = 8'h1b == io_state_in_14 ? 8'hc3 : _GEN_15898; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15900 = 8'h1c == io_state_in_14 ? 8'hfc : _GEN_15899; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15901 = 8'h1d == io_state_in_14 ? 8'hf5 : _GEN_15900; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15902 = 8'h1e == io_state_in_14 ? 8'hee : _GEN_15901; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15903 = 8'h1f == io_state_in_14 ? 8'he7 : _GEN_15902; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15904 = 8'h20 == io_state_in_14 ? 8'h3b : _GEN_15903; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15905 = 8'h21 == io_state_in_14 ? 8'h32 : _GEN_15904; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15906 = 8'h22 == io_state_in_14 ? 8'h29 : _GEN_15905; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15907 = 8'h23 == io_state_in_14 ? 8'h20 : _GEN_15906; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15908 = 8'h24 == io_state_in_14 ? 8'h1f : _GEN_15907; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15909 = 8'h25 == io_state_in_14 ? 8'h16 : _GEN_15908; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15910 = 8'h26 == io_state_in_14 ? 8'hd : _GEN_15909; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15911 = 8'h27 == io_state_in_14 ? 8'h4 : _GEN_15910; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15912 = 8'h28 == io_state_in_14 ? 8'h73 : _GEN_15911; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15913 = 8'h29 == io_state_in_14 ? 8'h7a : _GEN_15912; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15914 = 8'h2a == io_state_in_14 ? 8'h61 : _GEN_15913; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15915 = 8'h2b == io_state_in_14 ? 8'h68 : _GEN_15914; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15916 = 8'h2c == io_state_in_14 ? 8'h57 : _GEN_15915; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15917 = 8'h2d == io_state_in_14 ? 8'h5e : _GEN_15916; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15918 = 8'h2e == io_state_in_14 ? 8'h45 : _GEN_15917; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15919 = 8'h2f == io_state_in_14 ? 8'h4c : _GEN_15918; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15920 = 8'h30 == io_state_in_14 ? 8'hab : _GEN_15919; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15921 = 8'h31 == io_state_in_14 ? 8'ha2 : _GEN_15920; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15922 = 8'h32 == io_state_in_14 ? 8'hb9 : _GEN_15921; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15923 = 8'h33 == io_state_in_14 ? 8'hb0 : _GEN_15922; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15924 = 8'h34 == io_state_in_14 ? 8'h8f : _GEN_15923; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15925 = 8'h35 == io_state_in_14 ? 8'h86 : _GEN_15924; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15926 = 8'h36 == io_state_in_14 ? 8'h9d : _GEN_15925; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15927 = 8'h37 == io_state_in_14 ? 8'h94 : _GEN_15926; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15928 = 8'h38 == io_state_in_14 ? 8'he3 : _GEN_15927; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15929 = 8'h39 == io_state_in_14 ? 8'hea : _GEN_15928; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15930 = 8'h3a == io_state_in_14 ? 8'hf1 : _GEN_15929; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15931 = 8'h3b == io_state_in_14 ? 8'hf8 : _GEN_15930; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15932 = 8'h3c == io_state_in_14 ? 8'hc7 : _GEN_15931; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15933 = 8'h3d == io_state_in_14 ? 8'hce : _GEN_15932; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15934 = 8'h3e == io_state_in_14 ? 8'hd5 : _GEN_15933; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15935 = 8'h3f == io_state_in_14 ? 8'hdc : _GEN_15934; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15936 = 8'h40 == io_state_in_14 ? 8'h76 : _GEN_15935; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15937 = 8'h41 == io_state_in_14 ? 8'h7f : _GEN_15936; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15938 = 8'h42 == io_state_in_14 ? 8'h64 : _GEN_15937; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15939 = 8'h43 == io_state_in_14 ? 8'h6d : _GEN_15938; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15940 = 8'h44 == io_state_in_14 ? 8'h52 : _GEN_15939; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15941 = 8'h45 == io_state_in_14 ? 8'h5b : _GEN_15940; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15942 = 8'h46 == io_state_in_14 ? 8'h40 : _GEN_15941; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15943 = 8'h47 == io_state_in_14 ? 8'h49 : _GEN_15942; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15944 = 8'h48 == io_state_in_14 ? 8'h3e : _GEN_15943; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15945 = 8'h49 == io_state_in_14 ? 8'h37 : _GEN_15944; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15946 = 8'h4a == io_state_in_14 ? 8'h2c : _GEN_15945; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15947 = 8'h4b == io_state_in_14 ? 8'h25 : _GEN_15946; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15948 = 8'h4c == io_state_in_14 ? 8'h1a : _GEN_15947; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15949 = 8'h4d == io_state_in_14 ? 8'h13 : _GEN_15948; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15950 = 8'h4e == io_state_in_14 ? 8'h8 : _GEN_15949; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15951 = 8'h4f == io_state_in_14 ? 8'h1 : _GEN_15950; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15952 = 8'h50 == io_state_in_14 ? 8'he6 : _GEN_15951; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15953 = 8'h51 == io_state_in_14 ? 8'hef : _GEN_15952; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15954 = 8'h52 == io_state_in_14 ? 8'hf4 : _GEN_15953; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15955 = 8'h53 == io_state_in_14 ? 8'hfd : _GEN_15954; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15956 = 8'h54 == io_state_in_14 ? 8'hc2 : _GEN_15955; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15957 = 8'h55 == io_state_in_14 ? 8'hcb : _GEN_15956; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15958 = 8'h56 == io_state_in_14 ? 8'hd0 : _GEN_15957; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15959 = 8'h57 == io_state_in_14 ? 8'hd9 : _GEN_15958; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15960 = 8'h58 == io_state_in_14 ? 8'hae : _GEN_15959; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15961 = 8'h59 == io_state_in_14 ? 8'ha7 : _GEN_15960; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15962 = 8'h5a == io_state_in_14 ? 8'hbc : _GEN_15961; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15963 = 8'h5b == io_state_in_14 ? 8'hb5 : _GEN_15962; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15964 = 8'h5c == io_state_in_14 ? 8'h8a : _GEN_15963; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15965 = 8'h5d == io_state_in_14 ? 8'h83 : _GEN_15964; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15966 = 8'h5e == io_state_in_14 ? 8'h98 : _GEN_15965; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15967 = 8'h5f == io_state_in_14 ? 8'h91 : _GEN_15966; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15968 = 8'h60 == io_state_in_14 ? 8'h4d : _GEN_15967; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15969 = 8'h61 == io_state_in_14 ? 8'h44 : _GEN_15968; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15970 = 8'h62 == io_state_in_14 ? 8'h5f : _GEN_15969; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15971 = 8'h63 == io_state_in_14 ? 8'h56 : _GEN_15970; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15972 = 8'h64 == io_state_in_14 ? 8'h69 : _GEN_15971; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15973 = 8'h65 == io_state_in_14 ? 8'h60 : _GEN_15972; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15974 = 8'h66 == io_state_in_14 ? 8'h7b : _GEN_15973; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15975 = 8'h67 == io_state_in_14 ? 8'h72 : _GEN_15974; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15976 = 8'h68 == io_state_in_14 ? 8'h5 : _GEN_15975; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15977 = 8'h69 == io_state_in_14 ? 8'hc : _GEN_15976; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15978 = 8'h6a == io_state_in_14 ? 8'h17 : _GEN_15977; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15979 = 8'h6b == io_state_in_14 ? 8'h1e : _GEN_15978; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15980 = 8'h6c == io_state_in_14 ? 8'h21 : _GEN_15979; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15981 = 8'h6d == io_state_in_14 ? 8'h28 : _GEN_15980; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15982 = 8'h6e == io_state_in_14 ? 8'h33 : _GEN_15981; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15983 = 8'h6f == io_state_in_14 ? 8'h3a : _GEN_15982; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15984 = 8'h70 == io_state_in_14 ? 8'hdd : _GEN_15983; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15985 = 8'h71 == io_state_in_14 ? 8'hd4 : _GEN_15984; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15986 = 8'h72 == io_state_in_14 ? 8'hcf : _GEN_15985; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15987 = 8'h73 == io_state_in_14 ? 8'hc6 : _GEN_15986; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15988 = 8'h74 == io_state_in_14 ? 8'hf9 : _GEN_15987; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15989 = 8'h75 == io_state_in_14 ? 8'hf0 : _GEN_15988; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15990 = 8'h76 == io_state_in_14 ? 8'heb : _GEN_15989; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15991 = 8'h77 == io_state_in_14 ? 8'he2 : _GEN_15990; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15992 = 8'h78 == io_state_in_14 ? 8'h95 : _GEN_15991; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15993 = 8'h79 == io_state_in_14 ? 8'h9c : _GEN_15992; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15994 = 8'h7a == io_state_in_14 ? 8'h87 : _GEN_15993; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15995 = 8'h7b == io_state_in_14 ? 8'h8e : _GEN_15994; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15996 = 8'h7c == io_state_in_14 ? 8'hb1 : _GEN_15995; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15997 = 8'h7d == io_state_in_14 ? 8'hb8 : _GEN_15996; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15998 = 8'h7e == io_state_in_14 ? 8'ha3 : _GEN_15997; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_15999 = 8'h7f == io_state_in_14 ? 8'haa : _GEN_15998; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16000 = 8'h80 == io_state_in_14 ? 8'hec : _GEN_15999; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16001 = 8'h81 == io_state_in_14 ? 8'he5 : _GEN_16000; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16002 = 8'h82 == io_state_in_14 ? 8'hfe : _GEN_16001; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16003 = 8'h83 == io_state_in_14 ? 8'hf7 : _GEN_16002; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16004 = 8'h84 == io_state_in_14 ? 8'hc8 : _GEN_16003; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16005 = 8'h85 == io_state_in_14 ? 8'hc1 : _GEN_16004; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16006 = 8'h86 == io_state_in_14 ? 8'hda : _GEN_16005; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16007 = 8'h87 == io_state_in_14 ? 8'hd3 : _GEN_16006; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16008 = 8'h88 == io_state_in_14 ? 8'ha4 : _GEN_16007; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16009 = 8'h89 == io_state_in_14 ? 8'had : _GEN_16008; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16010 = 8'h8a == io_state_in_14 ? 8'hb6 : _GEN_16009; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16011 = 8'h8b == io_state_in_14 ? 8'hbf : _GEN_16010; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16012 = 8'h8c == io_state_in_14 ? 8'h80 : _GEN_16011; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16013 = 8'h8d == io_state_in_14 ? 8'h89 : _GEN_16012; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16014 = 8'h8e == io_state_in_14 ? 8'h92 : _GEN_16013; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16015 = 8'h8f == io_state_in_14 ? 8'h9b : _GEN_16014; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16016 = 8'h90 == io_state_in_14 ? 8'h7c : _GEN_16015; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16017 = 8'h91 == io_state_in_14 ? 8'h75 : _GEN_16016; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16018 = 8'h92 == io_state_in_14 ? 8'h6e : _GEN_16017; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16019 = 8'h93 == io_state_in_14 ? 8'h67 : _GEN_16018; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16020 = 8'h94 == io_state_in_14 ? 8'h58 : _GEN_16019; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16021 = 8'h95 == io_state_in_14 ? 8'h51 : _GEN_16020; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16022 = 8'h96 == io_state_in_14 ? 8'h4a : _GEN_16021; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16023 = 8'h97 == io_state_in_14 ? 8'h43 : _GEN_16022; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16024 = 8'h98 == io_state_in_14 ? 8'h34 : _GEN_16023; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16025 = 8'h99 == io_state_in_14 ? 8'h3d : _GEN_16024; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16026 = 8'h9a == io_state_in_14 ? 8'h26 : _GEN_16025; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16027 = 8'h9b == io_state_in_14 ? 8'h2f : _GEN_16026; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16028 = 8'h9c == io_state_in_14 ? 8'h10 : _GEN_16027; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16029 = 8'h9d == io_state_in_14 ? 8'h19 : _GEN_16028; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16030 = 8'h9e == io_state_in_14 ? 8'h2 : _GEN_16029; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16031 = 8'h9f == io_state_in_14 ? 8'hb : _GEN_16030; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16032 = 8'ha0 == io_state_in_14 ? 8'hd7 : _GEN_16031; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16033 = 8'ha1 == io_state_in_14 ? 8'hde : _GEN_16032; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16034 = 8'ha2 == io_state_in_14 ? 8'hc5 : _GEN_16033; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16035 = 8'ha3 == io_state_in_14 ? 8'hcc : _GEN_16034; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16036 = 8'ha4 == io_state_in_14 ? 8'hf3 : _GEN_16035; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16037 = 8'ha5 == io_state_in_14 ? 8'hfa : _GEN_16036; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16038 = 8'ha6 == io_state_in_14 ? 8'he1 : _GEN_16037; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16039 = 8'ha7 == io_state_in_14 ? 8'he8 : _GEN_16038; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16040 = 8'ha8 == io_state_in_14 ? 8'h9f : _GEN_16039; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16041 = 8'ha9 == io_state_in_14 ? 8'h96 : _GEN_16040; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16042 = 8'haa == io_state_in_14 ? 8'h8d : _GEN_16041; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16043 = 8'hab == io_state_in_14 ? 8'h84 : _GEN_16042; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16044 = 8'hac == io_state_in_14 ? 8'hbb : _GEN_16043; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16045 = 8'had == io_state_in_14 ? 8'hb2 : _GEN_16044; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16046 = 8'hae == io_state_in_14 ? 8'ha9 : _GEN_16045; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16047 = 8'haf == io_state_in_14 ? 8'ha0 : _GEN_16046; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16048 = 8'hb0 == io_state_in_14 ? 8'h47 : _GEN_16047; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16049 = 8'hb1 == io_state_in_14 ? 8'h4e : _GEN_16048; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16050 = 8'hb2 == io_state_in_14 ? 8'h55 : _GEN_16049; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16051 = 8'hb3 == io_state_in_14 ? 8'h5c : _GEN_16050; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16052 = 8'hb4 == io_state_in_14 ? 8'h63 : _GEN_16051; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16053 = 8'hb5 == io_state_in_14 ? 8'h6a : _GEN_16052; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16054 = 8'hb6 == io_state_in_14 ? 8'h71 : _GEN_16053; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16055 = 8'hb7 == io_state_in_14 ? 8'h78 : _GEN_16054; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16056 = 8'hb8 == io_state_in_14 ? 8'hf : _GEN_16055; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16057 = 8'hb9 == io_state_in_14 ? 8'h6 : _GEN_16056; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16058 = 8'hba == io_state_in_14 ? 8'h1d : _GEN_16057; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16059 = 8'hbb == io_state_in_14 ? 8'h14 : _GEN_16058; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16060 = 8'hbc == io_state_in_14 ? 8'h2b : _GEN_16059; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16061 = 8'hbd == io_state_in_14 ? 8'h22 : _GEN_16060; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16062 = 8'hbe == io_state_in_14 ? 8'h39 : _GEN_16061; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16063 = 8'hbf == io_state_in_14 ? 8'h30 : _GEN_16062; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16064 = 8'hc0 == io_state_in_14 ? 8'h9a : _GEN_16063; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16065 = 8'hc1 == io_state_in_14 ? 8'h93 : _GEN_16064; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16066 = 8'hc2 == io_state_in_14 ? 8'h88 : _GEN_16065; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16067 = 8'hc3 == io_state_in_14 ? 8'h81 : _GEN_16066; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16068 = 8'hc4 == io_state_in_14 ? 8'hbe : _GEN_16067; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16069 = 8'hc5 == io_state_in_14 ? 8'hb7 : _GEN_16068; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16070 = 8'hc6 == io_state_in_14 ? 8'hac : _GEN_16069; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16071 = 8'hc7 == io_state_in_14 ? 8'ha5 : _GEN_16070; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16072 = 8'hc8 == io_state_in_14 ? 8'hd2 : _GEN_16071; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16073 = 8'hc9 == io_state_in_14 ? 8'hdb : _GEN_16072; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16074 = 8'hca == io_state_in_14 ? 8'hc0 : _GEN_16073; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16075 = 8'hcb == io_state_in_14 ? 8'hc9 : _GEN_16074; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16076 = 8'hcc == io_state_in_14 ? 8'hf6 : _GEN_16075; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16077 = 8'hcd == io_state_in_14 ? 8'hff : _GEN_16076; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16078 = 8'hce == io_state_in_14 ? 8'he4 : _GEN_16077; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16079 = 8'hcf == io_state_in_14 ? 8'hed : _GEN_16078; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16080 = 8'hd0 == io_state_in_14 ? 8'ha : _GEN_16079; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16081 = 8'hd1 == io_state_in_14 ? 8'h3 : _GEN_16080; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16082 = 8'hd2 == io_state_in_14 ? 8'h18 : _GEN_16081; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16083 = 8'hd3 == io_state_in_14 ? 8'h11 : _GEN_16082; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16084 = 8'hd4 == io_state_in_14 ? 8'h2e : _GEN_16083; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16085 = 8'hd5 == io_state_in_14 ? 8'h27 : _GEN_16084; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16086 = 8'hd6 == io_state_in_14 ? 8'h3c : _GEN_16085; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16087 = 8'hd7 == io_state_in_14 ? 8'h35 : _GEN_16086; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16088 = 8'hd8 == io_state_in_14 ? 8'h42 : _GEN_16087; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16089 = 8'hd9 == io_state_in_14 ? 8'h4b : _GEN_16088; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16090 = 8'hda == io_state_in_14 ? 8'h50 : _GEN_16089; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16091 = 8'hdb == io_state_in_14 ? 8'h59 : _GEN_16090; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16092 = 8'hdc == io_state_in_14 ? 8'h66 : _GEN_16091; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16093 = 8'hdd == io_state_in_14 ? 8'h6f : _GEN_16092; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16094 = 8'hde == io_state_in_14 ? 8'h74 : _GEN_16093; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16095 = 8'hdf == io_state_in_14 ? 8'h7d : _GEN_16094; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16096 = 8'he0 == io_state_in_14 ? 8'ha1 : _GEN_16095; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16097 = 8'he1 == io_state_in_14 ? 8'ha8 : _GEN_16096; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16098 = 8'he2 == io_state_in_14 ? 8'hb3 : _GEN_16097; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16099 = 8'he3 == io_state_in_14 ? 8'hba : _GEN_16098; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16100 = 8'he4 == io_state_in_14 ? 8'h85 : _GEN_16099; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16101 = 8'he5 == io_state_in_14 ? 8'h8c : _GEN_16100; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16102 = 8'he6 == io_state_in_14 ? 8'h97 : _GEN_16101; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16103 = 8'he7 == io_state_in_14 ? 8'h9e : _GEN_16102; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16104 = 8'he8 == io_state_in_14 ? 8'he9 : _GEN_16103; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16105 = 8'he9 == io_state_in_14 ? 8'he0 : _GEN_16104; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16106 = 8'hea == io_state_in_14 ? 8'hfb : _GEN_16105; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16107 = 8'heb == io_state_in_14 ? 8'hf2 : _GEN_16106; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16108 = 8'hec == io_state_in_14 ? 8'hcd : _GEN_16107; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16109 = 8'hed == io_state_in_14 ? 8'hc4 : _GEN_16108; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16110 = 8'hee == io_state_in_14 ? 8'hdf : _GEN_16109; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16111 = 8'hef == io_state_in_14 ? 8'hd6 : _GEN_16110; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16112 = 8'hf0 == io_state_in_14 ? 8'h31 : _GEN_16111; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16113 = 8'hf1 == io_state_in_14 ? 8'h38 : _GEN_16112; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16114 = 8'hf2 == io_state_in_14 ? 8'h23 : _GEN_16113; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16115 = 8'hf3 == io_state_in_14 ? 8'h2a : _GEN_16114; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16116 = 8'hf4 == io_state_in_14 ? 8'h15 : _GEN_16115; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16117 = 8'hf5 == io_state_in_14 ? 8'h1c : _GEN_16116; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16118 = 8'hf6 == io_state_in_14 ? 8'h7 : _GEN_16117; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16119 = 8'hf7 == io_state_in_14 ? 8'he : _GEN_16118; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16120 = 8'hf8 == io_state_in_14 ? 8'h79 : _GEN_16119; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16121 = 8'hf9 == io_state_in_14 ? 8'h70 : _GEN_16120; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16122 = 8'hfa == io_state_in_14 ? 8'h6b : _GEN_16121; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16123 = 8'hfb == io_state_in_14 ? 8'h62 : _GEN_16122; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16124 = 8'hfc == io_state_in_14 ? 8'h5d : _GEN_16123; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16125 = 8'hfd == io_state_in_14 ? 8'h54 : _GEN_16124; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16126 = 8'hfe == io_state_in_14 ? 8'h4f : _GEN_16125; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _GEN_16127 = 8'hff == io_state_in_14 ? 8'h46 : _GEN_16126; // @[InvMixColumns.scala 144:{68,68}]
  wire [7:0] _tmp_state_15_T_1 = _tmp_state_15_T ^ _GEN_16127; // @[InvMixColumns.scala 144:68]
  wire [7:0] _GEN_16129 = 8'h1 == io_state_in_15 ? 8'he : 8'h0; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16130 = 8'h2 == io_state_in_15 ? 8'h1c : _GEN_16129; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16131 = 8'h3 == io_state_in_15 ? 8'h12 : _GEN_16130; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16132 = 8'h4 == io_state_in_15 ? 8'h38 : _GEN_16131; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16133 = 8'h5 == io_state_in_15 ? 8'h36 : _GEN_16132; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16134 = 8'h6 == io_state_in_15 ? 8'h24 : _GEN_16133; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16135 = 8'h7 == io_state_in_15 ? 8'h2a : _GEN_16134; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16136 = 8'h8 == io_state_in_15 ? 8'h70 : _GEN_16135; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16137 = 8'h9 == io_state_in_15 ? 8'h7e : _GEN_16136; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16138 = 8'ha == io_state_in_15 ? 8'h6c : _GEN_16137; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16139 = 8'hb == io_state_in_15 ? 8'h62 : _GEN_16138; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16140 = 8'hc == io_state_in_15 ? 8'h48 : _GEN_16139; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16141 = 8'hd == io_state_in_15 ? 8'h46 : _GEN_16140; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16142 = 8'he == io_state_in_15 ? 8'h54 : _GEN_16141; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16143 = 8'hf == io_state_in_15 ? 8'h5a : _GEN_16142; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16144 = 8'h10 == io_state_in_15 ? 8'he0 : _GEN_16143; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16145 = 8'h11 == io_state_in_15 ? 8'hee : _GEN_16144; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16146 = 8'h12 == io_state_in_15 ? 8'hfc : _GEN_16145; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16147 = 8'h13 == io_state_in_15 ? 8'hf2 : _GEN_16146; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16148 = 8'h14 == io_state_in_15 ? 8'hd8 : _GEN_16147; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16149 = 8'h15 == io_state_in_15 ? 8'hd6 : _GEN_16148; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16150 = 8'h16 == io_state_in_15 ? 8'hc4 : _GEN_16149; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16151 = 8'h17 == io_state_in_15 ? 8'hca : _GEN_16150; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16152 = 8'h18 == io_state_in_15 ? 8'h90 : _GEN_16151; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16153 = 8'h19 == io_state_in_15 ? 8'h9e : _GEN_16152; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16154 = 8'h1a == io_state_in_15 ? 8'h8c : _GEN_16153; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16155 = 8'h1b == io_state_in_15 ? 8'h82 : _GEN_16154; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16156 = 8'h1c == io_state_in_15 ? 8'ha8 : _GEN_16155; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16157 = 8'h1d == io_state_in_15 ? 8'ha6 : _GEN_16156; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16158 = 8'h1e == io_state_in_15 ? 8'hb4 : _GEN_16157; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16159 = 8'h1f == io_state_in_15 ? 8'hba : _GEN_16158; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16160 = 8'h20 == io_state_in_15 ? 8'hdb : _GEN_16159; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16161 = 8'h21 == io_state_in_15 ? 8'hd5 : _GEN_16160; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16162 = 8'h22 == io_state_in_15 ? 8'hc7 : _GEN_16161; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16163 = 8'h23 == io_state_in_15 ? 8'hc9 : _GEN_16162; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16164 = 8'h24 == io_state_in_15 ? 8'he3 : _GEN_16163; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16165 = 8'h25 == io_state_in_15 ? 8'hed : _GEN_16164; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16166 = 8'h26 == io_state_in_15 ? 8'hff : _GEN_16165; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16167 = 8'h27 == io_state_in_15 ? 8'hf1 : _GEN_16166; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16168 = 8'h28 == io_state_in_15 ? 8'hab : _GEN_16167; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16169 = 8'h29 == io_state_in_15 ? 8'ha5 : _GEN_16168; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16170 = 8'h2a == io_state_in_15 ? 8'hb7 : _GEN_16169; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16171 = 8'h2b == io_state_in_15 ? 8'hb9 : _GEN_16170; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16172 = 8'h2c == io_state_in_15 ? 8'h93 : _GEN_16171; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16173 = 8'h2d == io_state_in_15 ? 8'h9d : _GEN_16172; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16174 = 8'h2e == io_state_in_15 ? 8'h8f : _GEN_16173; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16175 = 8'h2f == io_state_in_15 ? 8'h81 : _GEN_16174; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16176 = 8'h30 == io_state_in_15 ? 8'h3b : _GEN_16175; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16177 = 8'h31 == io_state_in_15 ? 8'h35 : _GEN_16176; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16178 = 8'h32 == io_state_in_15 ? 8'h27 : _GEN_16177; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16179 = 8'h33 == io_state_in_15 ? 8'h29 : _GEN_16178; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16180 = 8'h34 == io_state_in_15 ? 8'h3 : _GEN_16179; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16181 = 8'h35 == io_state_in_15 ? 8'hd : _GEN_16180; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16182 = 8'h36 == io_state_in_15 ? 8'h1f : _GEN_16181; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16183 = 8'h37 == io_state_in_15 ? 8'h11 : _GEN_16182; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16184 = 8'h38 == io_state_in_15 ? 8'h4b : _GEN_16183; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16185 = 8'h39 == io_state_in_15 ? 8'h45 : _GEN_16184; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16186 = 8'h3a == io_state_in_15 ? 8'h57 : _GEN_16185; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16187 = 8'h3b == io_state_in_15 ? 8'h59 : _GEN_16186; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16188 = 8'h3c == io_state_in_15 ? 8'h73 : _GEN_16187; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16189 = 8'h3d == io_state_in_15 ? 8'h7d : _GEN_16188; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16190 = 8'h3e == io_state_in_15 ? 8'h6f : _GEN_16189; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16191 = 8'h3f == io_state_in_15 ? 8'h61 : _GEN_16190; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16192 = 8'h40 == io_state_in_15 ? 8'had : _GEN_16191; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16193 = 8'h41 == io_state_in_15 ? 8'ha3 : _GEN_16192; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16194 = 8'h42 == io_state_in_15 ? 8'hb1 : _GEN_16193; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16195 = 8'h43 == io_state_in_15 ? 8'hbf : _GEN_16194; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16196 = 8'h44 == io_state_in_15 ? 8'h95 : _GEN_16195; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16197 = 8'h45 == io_state_in_15 ? 8'h9b : _GEN_16196; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16198 = 8'h46 == io_state_in_15 ? 8'h89 : _GEN_16197; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16199 = 8'h47 == io_state_in_15 ? 8'h87 : _GEN_16198; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16200 = 8'h48 == io_state_in_15 ? 8'hdd : _GEN_16199; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16201 = 8'h49 == io_state_in_15 ? 8'hd3 : _GEN_16200; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16202 = 8'h4a == io_state_in_15 ? 8'hc1 : _GEN_16201; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16203 = 8'h4b == io_state_in_15 ? 8'hcf : _GEN_16202; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16204 = 8'h4c == io_state_in_15 ? 8'he5 : _GEN_16203; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16205 = 8'h4d == io_state_in_15 ? 8'heb : _GEN_16204; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16206 = 8'h4e == io_state_in_15 ? 8'hf9 : _GEN_16205; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16207 = 8'h4f == io_state_in_15 ? 8'hf7 : _GEN_16206; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16208 = 8'h50 == io_state_in_15 ? 8'h4d : _GEN_16207; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16209 = 8'h51 == io_state_in_15 ? 8'h43 : _GEN_16208; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16210 = 8'h52 == io_state_in_15 ? 8'h51 : _GEN_16209; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16211 = 8'h53 == io_state_in_15 ? 8'h5f : _GEN_16210; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16212 = 8'h54 == io_state_in_15 ? 8'h75 : _GEN_16211; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16213 = 8'h55 == io_state_in_15 ? 8'h7b : _GEN_16212; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16214 = 8'h56 == io_state_in_15 ? 8'h69 : _GEN_16213; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16215 = 8'h57 == io_state_in_15 ? 8'h67 : _GEN_16214; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16216 = 8'h58 == io_state_in_15 ? 8'h3d : _GEN_16215; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16217 = 8'h59 == io_state_in_15 ? 8'h33 : _GEN_16216; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16218 = 8'h5a == io_state_in_15 ? 8'h21 : _GEN_16217; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16219 = 8'h5b == io_state_in_15 ? 8'h2f : _GEN_16218; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16220 = 8'h5c == io_state_in_15 ? 8'h5 : _GEN_16219; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16221 = 8'h5d == io_state_in_15 ? 8'hb : _GEN_16220; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16222 = 8'h5e == io_state_in_15 ? 8'h19 : _GEN_16221; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16223 = 8'h5f == io_state_in_15 ? 8'h17 : _GEN_16222; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16224 = 8'h60 == io_state_in_15 ? 8'h76 : _GEN_16223; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16225 = 8'h61 == io_state_in_15 ? 8'h78 : _GEN_16224; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16226 = 8'h62 == io_state_in_15 ? 8'h6a : _GEN_16225; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16227 = 8'h63 == io_state_in_15 ? 8'h64 : _GEN_16226; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16228 = 8'h64 == io_state_in_15 ? 8'h4e : _GEN_16227; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16229 = 8'h65 == io_state_in_15 ? 8'h40 : _GEN_16228; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16230 = 8'h66 == io_state_in_15 ? 8'h52 : _GEN_16229; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16231 = 8'h67 == io_state_in_15 ? 8'h5c : _GEN_16230; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16232 = 8'h68 == io_state_in_15 ? 8'h6 : _GEN_16231; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16233 = 8'h69 == io_state_in_15 ? 8'h8 : _GEN_16232; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16234 = 8'h6a == io_state_in_15 ? 8'h1a : _GEN_16233; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16235 = 8'h6b == io_state_in_15 ? 8'h14 : _GEN_16234; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16236 = 8'h6c == io_state_in_15 ? 8'h3e : _GEN_16235; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16237 = 8'h6d == io_state_in_15 ? 8'h30 : _GEN_16236; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16238 = 8'h6e == io_state_in_15 ? 8'h22 : _GEN_16237; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16239 = 8'h6f == io_state_in_15 ? 8'h2c : _GEN_16238; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16240 = 8'h70 == io_state_in_15 ? 8'h96 : _GEN_16239; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16241 = 8'h71 == io_state_in_15 ? 8'h98 : _GEN_16240; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16242 = 8'h72 == io_state_in_15 ? 8'h8a : _GEN_16241; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16243 = 8'h73 == io_state_in_15 ? 8'h84 : _GEN_16242; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16244 = 8'h74 == io_state_in_15 ? 8'hae : _GEN_16243; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16245 = 8'h75 == io_state_in_15 ? 8'ha0 : _GEN_16244; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16246 = 8'h76 == io_state_in_15 ? 8'hb2 : _GEN_16245; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16247 = 8'h77 == io_state_in_15 ? 8'hbc : _GEN_16246; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16248 = 8'h78 == io_state_in_15 ? 8'he6 : _GEN_16247; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16249 = 8'h79 == io_state_in_15 ? 8'he8 : _GEN_16248; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16250 = 8'h7a == io_state_in_15 ? 8'hfa : _GEN_16249; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16251 = 8'h7b == io_state_in_15 ? 8'hf4 : _GEN_16250; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16252 = 8'h7c == io_state_in_15 ? 8'hde : _GEN_16251; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16253 = 8'h7d == io_state_in_15 ? 8'hd0 : _GEN_16252; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16254 = 8'h7e == io_state_in_15 ? 8'hc2 : _GEN_16253; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16255 = 8'h7f == io_state_in_15 ? 8'hcc : _GEN_16254; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16256 = 8'h80 == io_state_in_15 ? 8'h41 : _GEN_16255; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16257 = 8'h81 == io_state_in_15 ? 8'h4f : _GEN_16256; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16258 = 8'h82 == io_state_in_15 ? 8'h5d : _GEN_16257; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16259 = 8'h83 == io_state_in_15 ? 8'h53 : _GEN_16258; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16260 = 8'h84 == io_state_in_15 ? 8'h79 : _GEN_16259; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16261 = 8'h85 == io_state_in_15 ? 8'h77 : _GEN_16260; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16262 = 8'h86 == io_state_in_15 ? 8'h65 : _GEN_16261; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16263 = 8'h87 == io_state_in_15 ? 8'h6b : _GEN_16262; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16264 = 8'h88 == io_state_in_15 ? 8'h31 : _GEN_16263; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16265 = 8'h89 == io_state_in_15 ? 8'h3f : _GEN_16264; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16266 = 8'h8a == io_state_in_15 ? 8'h2d : _GEN_16265; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16267 = 8'h8b == io_state_in_15 ? 8'h23 : _GEN_16266; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16268 = 8'h8c == io_state_in_15 ? 8'h9 : _GEN_16267; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16269 = 8'h8d == io_state_in_15 ? 8'h7 : _GEN_16268; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16270 = 8'h8e == io_state_in_15 ? 8'h15 : _GEN_16269; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16271 = 8'h8f == io_state_in_15 ? 8'h1b : _GEN_16270; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16272 = 8'h90 == io_state_in_15 ? 8'ha1 : _GEN_16271; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16273 = 8'h91 == io_state_in_15 ? 8'haf : _GEN_16272; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16274 = 8'h92 == io_state_in_15 ? 8'hbd : _GEN_16273; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16275 = 8'h93 == io_state_in_15 ? 8'hb3 : _GEN_16274; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16276 = 8'h94 == io_state_in_15 ? 8'h99 : _GEN_16275; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16277 = 8'h95 == io_state_in_15 ? 8'h97 : _GEN_16276; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16278 = 8'h96 == io_state_in_15 ? 8'h85 : _GEN_16277; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16279 = 8'h97 == io_state_in_15 ? 8'h8b : _GEN_16278; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16280 = 8'h98 == io_state_in_15 ? 8'hd1 : _GEN_16279; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16281 = 8'h99 == io_state_in_15 ? 8'hdf : _GEN_16280; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16282 = 8'h9a == io_state_in_15 ? 8'hcd : _GEN_16281; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16283 = 8'h9b == io_state_in_15 ? 8'hc3 : _GEN_16282; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16284 = 8'h9c == io_state_in_15 ? 8'he9 : _GEN_16283; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16285 = 8'h9d == io_state_in_15 ? 8'he7 : _GEN_16284; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16286 = 8'h9e == io_state_in_15 ? 8'hf5 : _GEN_16285; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16287 = 8'h9f == io_state_in_15 ? 8'hfb : _GEN_16286; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16288 = 8'ha0 == io_state_in_15 ? 8'h9a : _GEN_16287; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16289 = 8'ha1 == io_state_in_15 ? 8'h94 : _GEN_16288; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16290 = 8'ha2 == io_state_in_15 ? 8'h86 : _GEN_16289; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16291 = 8'ha3 == io_state_in_15 ? 8'h88 : _GEN_16290; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16292 = 8'ha4 == io_state_in_15 ? 8'ha2 : _GEN_16291; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16293 = 8'ha5 == io_state_in_15 ? 8'hac : _GEN_16292; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16294 = 8'ha6 == io_state_in_15 ? 8'hbe : _GEN_16293; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16295 = 8'ha7 == io_state_in_15 ? 8'hb0 : _GEN_16294; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16296 = 8'ha8 == io_state_in_15 ? 8'hea : _GEN_16295; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16297 = 8'ha9 == io_state_in_15 ? 8'he4 : _GEN_16296; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16298 = 8'haa == io_state_in_15 ? 8'hf6 : _GEN_16297; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16299 = 8'hab == io_state_in_15 ? 8'hf8 : _GEN_16298; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16300 = 8'hac == io_state_in_15 ? 8'hd2 : _GEN_16299; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16301 = 8'had == io_state_in_15 ? 8'hdc : _GEN_16300; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16302 = 8'hae == io_state_in_15 ? 8'hce : _GEN_16301; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16303 = 8'haf == io_state_in_15 ? 8'hc0 : _GEN_16302; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16304 = 8'hb0 == io_state_in_15 ? 8'h7a : _GEN_16303; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16305 = 8'hb1 == io_state_in_15 ? 8'h74 : _GEN_16304; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16306 = 8'hb2 == io_state_in_15 ? 8'h66 : _GEN_16305; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16307 = 8'hb3 == io_state_in_15 ? 8'h68 : _GEN_16306; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16308 = 8'hb4 == io_state_in_15 ? 8'h42 : _GEN_16307; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16309 = 8'hb5 == io_state_in_15 ? 8'h4c : _GEN_16308; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16310 = 8'hb6 == io_state_in_15 ? 8'h5e : _GEN_16309; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16311 = 8'hb7 == io_state_in_15 ? 8'h50 : _GEN_16310; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16312 = 8'hb8 == io_state_in_15 ? 8'ha : _GEN_16311; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16313 = 8'hb9 == io_state_in_15 ? 8'h4 : _GEN_16312; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16314 = 8'hba == io_state_in_15 ? 8'h16 : _GEN_16313; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16315 = 8'hbb == io_state_in_15 ? 8'h18 : _GEN_16314; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16316 = 8'hbc == io_state_in_15 ? 8'h32 : _GEN_16315; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16317 = 8'hbd == io_state_in_15 ? 8'h3c : _GEN_16316; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16318 = 8'hbe == io_state_in_15 ? 8'h2e : _GEN_16317; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16319 = 8'hbf == io_state_in_15 ? 8'h20 : _GEN_16318; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16320 = 8'hc0 == io_state_in_15 ? 8'hec : _GEN_16319; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16321 = 8'hc1 == io_state_in_15 ? 8'he2 : _GEN_16320; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16322 = 8'hc2 == io_state_in_15 ? 8'hf0 : _GEN_16321; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16323 = 8'hc3 == io_state_in_15 ? 8'hfe : _GEN_16322; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16324 = 8'hc4 == io_state_in_15 ? 8'hd4 : _GEN_16323; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16325 = 8'hc5 == io_state_in_15 ? 8'hda : _GEN_16324; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16326 = 8'hc6 == io_state_in_15 ? 8'hc8 : _GEN_16325; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16327 = 8'hc7 == io_state_in_15 ? 8'hc6 : _GEN_16326; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16328 = 8'hc8 == io_state_in_15 ? 8'h9c : _GEN_16327; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16329 = 8'hc9 == io_state_in_15 ? 8'h92 : _GEN_16328; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16330 = 8'hca == io_state_in_15 ? 8'h80 : _GEN_16329; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16331 = 8'hcb == io_state_in_15 ? 8'h8e : _GEN_16330; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16332 = 8'hcc == io_state_in_15 ? 8'ha4 : _GEN_16331; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16333 = 8'hcd == io_state_in_15 ? 8'haa : _GEN_16332; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16334 = 8'hce == io_state_in_15 ? 8'hb8 : _GEN_16333; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16335 = 8'hcf == io_state_in_15 ? 8'hb6 : _GEN_16334; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16336 = 8'hd0 == io_state_in_15 ? 8'hc : _GEN_16335; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16337 = 8'hd1 == io_state_in_15 ? 8'h2 : _GEN_16336; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16338 = 8'hd2 == io_state_in_15 ? 8'h10 : _GEN_16337; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16339 = 8'hd3 == io_state_in_15 ? 8'h1e : _GEN_16338; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16340 = 8'hd4 == io_state_in_15 ? 8'h34 : _GEN_16339; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16341 = 8'hd5 == io_state_in_15 ? 8'h3a : _GEN_16340; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16342 = 8'hd6 == io_state_in_15 ? 8'h28 : _GEN_16341; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16343 = 8'hd7 == io_state_in_15 ? 8'h26 : _GEN_16342; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16344 = 8'hd8 == io_state_in_15 ? 8'h7c : _GEN_16343; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16345 = 8'hd9 == io_state_in_15 ? 8'h72 : _GEN_16344; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16346 = 8'hda == io_state_in_15 ? 8'h60 : _GEN_16345; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16347 = 8'hdb == io_state_in_15 ? 8'h6e : _GEN_16346; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16348 = 8'hdc == io_state_in_15 ? 8'h44 : _GEN_16347; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16349 = 8'hdd == io_state_in_15 ? 8'h4a : _GEN_16348; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16350 = 8'hde == io_state_in_15 ? 8'h58 : _GEN_16349; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16351 = 8'hdf == io_state_in_15 ? 8'h56 : _GEN_16350; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16352 = 8'he0 == io_state_in_15 ? 8'h37 : _GEN_16351; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16353 = 8'he1 == io_state_in_15 ? 8'h39 : _GEN_16352; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16354 = 8'he2 == io_state_in_15 ? 8'h2b : _GEN_16353; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16355 = 8'he3 == io_state_in_15 ? 8'h25 : _GEN_16354; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16356 = 8'he4 == io_state_in_15 ? 8'hf : _GEN_16355; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16357 = 8'he5 == io_state_in_15 ? 8'h1 : _GEN_16356; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16358 = 8'he6 == io_state_in_15 ? 8'h13 : _GEN_16357; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16359 = 8'he7 == io_state_in_15 ? 8'h1d : _GEN_16358; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16360 = 8'he8 == io_state_in_15 ? 8'h47 : _GEN_16359; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16361 = 8'he9 == io_state_in_15 ? 8'h49 : _GEN_16360; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16362 = 8'hea == io_state_in_15 ? 8'h5b : _GEN_16361; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16363 = 8'heb == io_state_in_15 ? 8'h55 : _GEN_16362; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16364 = 8'hec == io_state_in_15 ? 8'h7f : _GEN_16363; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16365 = 8'hed == io_state_in_15 ? 8'h71 : _GEN_16364; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16366 = 8'hee == io_state_in_15 ? 8'h63 : _GEN_16365; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16367 = 8'hef == io_state_in_15 ? 8'h6d : _GEN_16366; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16368 = 8'hf0 == io_state_in_15 ? 8'hd7 : _GEN_16367; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16369 = 8'hf1 == io_state_in_15 ? 8'hd9 : _GEN_16368; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16370 = 8'hf2 == io_state_in_15 ? 8'hcb : _GEN_16369; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16371 = 8'hf3 == io_state_in_15 ? 8'hc5 : _GEN_16370; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16372 = 8'hf4 == io_state_in_15 ? 8'hef : _GEN_16371; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16373 = 8'hf5 == io_state_in_15 ? 8'he1 : _GEN_16372; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16374 = 8'hf6 == io_state_in_15 ? 8'hf3 : _GEN_16373; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16375 = 8'hf7 == io_state_in_15 ? 8'hfd : _GEN_16374; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16376 = 8'hf8 == io_state_in_15 ? 8'ha7 : _GEN_16375; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16377 = 8'hf9 == io_state_in_15 ? 8'ha9 : _GEN_16376; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16378 = 8'hfa == io_state_in_15 ? 8'hbb : _GEN_16377; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16379 = 8'hfb == io_state_in_15 ? 8'hb5 : _GEN_16378; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16380 = 8'hfc == io_state_in_15 ? 8'h9f : _GEN_16379; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16381 = 8'hfd == io_state_in_15 ? 8'h91 : _GEN_16380; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16382 = 8'hfe == io_state_in_15 ? 8'h83 : _GEN_16381; // @[InvMixColumns.scala 144:{93,93}]
  wire [7:0] _GEN_16383 = 8'hff == io_state_in_15 ? 8'h8d : _GEN_16382; // @[InvMixColumns.scala 144:{93,93}]
  assign io_state_out_0 = _tmp_state_0_T_1 ^ _GEN_1023; // @[InvMixColumns.scala 126:89]
  assign io_state_out_1 = _tmp_state_1_T_1 ^ _GEN_2047; // @[InvMixColumns.scala 127:89]
  assign io_state_out_2 = _tmp_state_2_T_1 ^ _GEN_3071; // @[InvMixColumns.scala 128:89]
  assign io_state_out_3 = _tmp_state_3_T_1 ^ _GEN_4095; // @[InvMixColumns.scala 129:89]
  assign io_state_out_4 = _tmp_state_4_T_1 ^ _GEN_5119; // @[InvMixColumns.scala 131:89]
  assign io_state_out_5 = _tmp_state_5_T_1 ^ _GEN_6143; // @[InvMixColumns.scala 132:89]
  assign io_state_out_6 = _tmp_state_6_T_1 ^ _GEN_7167; // @[InvMixColumns.scala 133:89]
  assign io_state_out_7 = _tmp_state_7_T_1 ^ _GEN_8191; // @[InvMixColumns.scala 134:89]
  assign io_state_out_8 = _tmp_state_8_T_1 ^ _GEN_9215; // @[InvMixColumns.scala 136:90]
  assign io_state_out_9 = _tmp_state_9_T_1 ^ _GEN_10239; // @[InvMixColumns.scala 137:90]
  assign io_state_out_10 = _tmp_state_10_T_1 ^ _GEN_11263; // @[InvMixColumns.scala 138:91]
  assign io_state_out_11 = _tmp_state_11_T_1 ^ _GEN_12287; // @[InvMixColumns.scala 139:91]
  assign io_state_out_12 = _tmp_state_12_T_1 ^ _GEN_13311; // @[InvMixColumns.scala 141:93]
  assign io_state_out_13 = _tmp_state_13_T_1 ^ _GEN_14335; // @[InvMixColumns.scala 142:93]
  assign io_state_out_14 = _tmp_state_14_T_1 ^ _GEN_15359; // @[InvMixColumns.scala 143:93]
  assign io_state_out_15 = _tmp_state_15_T_1 ^ _GEN_16383; // @[InvMixColumns.scala 144:93]
endmodule
module InvCipher(
  input        clock,
  input        reset,
  input  [7:0] io_ciphertext_0,
  input  [7:0] io_ciphertext_1,
  input  [7:0] io_ciphertext_2,
  input  [7:0] io_ciphertext_3,
  input  [7:0] io_ciphertext_4,
  input  [7:0] io_ciphertext_5,
  input  [7:0] io_ciphertext_6,
  input  [7:0] io_ciphertext_7,
  input  [7:0] io_ciphertext_8,
  input  [7:0] io_ciphertext_9,
  input  [7:0] io_ciphertext_10,
  input  [7:0] io_ciphertext_11,
  input  [7:0] io_ciphertext_12,
  input  [7:0] io_ciphertext_13,
  input  [7:0] io_ciphertext_14,
  input  [7:0] io_ciphertext_15,
  input  [7:0] io_roundKey_0,
  input  [7:0] io_roundKey_1,
  input  [7:0] io_roundKey_2,
  input  [7:0] io_roundKey_3,
  input  [7:0] io_roundKey_4,
  input  [7:0] io_roundKey_5,
  input  [7:0] io_roundKey_6,
  input  [7:0] io_roundKey_7,
  input  [7:0] io_roundKey_8,
  input  [7:0] io_roundKey_9,
  input  [7:0] io_roundKey_10,
  input  [7:0] io_roundKey_11,
  input  [7:0] io_roundKey_12,
  input  [7:0] io_roundKey_13,
  input  [7:0] io_roundKey_14,
  input  [7:0] io_roundKey_15,
  input        io_start,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15,
  output       io_state_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] AddRoundKeyModule_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] InvSubBytesModule_io_state_in_0; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_1; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_2; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_3; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_4; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_5; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_6; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_7; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_8; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_9; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_10; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_11; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_12; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_13; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_14; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_15; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_0; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_1; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_2; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_3; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_4; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_5; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_6; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_7; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_8; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_9; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_10; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_11; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_12; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_13; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_14; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_15; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvShiftRowsModule_io_state_in_0; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_1; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_2; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_3; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_4; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_5; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_6; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_7; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_8; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_9; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_10; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_11; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_12; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_13; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_14; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_15; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_0; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_1; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_2; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_3; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_4; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_5; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_6; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_7; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_8; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_9; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_10; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_11; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_12; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_13; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_14; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_15; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvMixColumnsModule_io_state_in_0; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_1; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_2; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_3; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_4; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_5; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_6; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_7; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_8; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_9; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_10; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_11; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_12; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_13; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_14; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_15; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_0; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_1; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_2; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_3; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_4; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_5; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_6; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_7; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_8; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_9; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_10; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_11; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_12; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_13; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_14; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_15; // @[InvMixColumns.scala 154:64]
  reg [7:0] state_0; // @[InvCipher.scala 31:22]
  reg [7:0] state_1; // @[InvCipher.scala 31:22]
  reg [7:0] state_2; // @[InvCipher.scala 31:22]
  reg [7:0] state_3; // @[InvCipher.scala 31:22]
  reg [7:0] state_4; // @[InvCipher.scala 31:22]
  reg [7:0] state_5; // @[InvCipher.scala 31:22]
  reg [7:0] state_6; // @[InvCipher.scala 31:22]
  reg [7:0] state_7; // @[InvCipher.scala 31:22]
  reg [7:0] state_8; // @[InvCipher.scala 31:22]
  reg [7:0] state_9; // @[InvCipher.scala 31:22]
  reg [7:0] state_10; // @[InvCipher.scala 31:22]
  reg [7:0] state_11; // @[InvCipher.scala 31:22]
  reg [7:0] state_12; // @[InvCipher.scala 31:22]
  reg [7:0] state_13; // @[InvCipher.scala 31:22]
  reg [7:0] state_14; // @[InvCipher.scala 31:22]
  reg [7:0] state_15; // @[InvCipher.scala 31:22]
  reg [3:0] rounds; // @[InvCipher.scala 32:23]
  reg [1:0] STM; // @[InvCipher.scala 36:20]
  wire [3:0] _rounds_T_1 = rounds + 4'h1; // @[InvCipher.scala 46:24]
  wire [1:0] _GEN_1 = rounds == 4'ha ? 2'h0 : STM; // @[InvCipher.scala 51:29 52:13 36:20]
  wire  _io_state_out_valid_T = rounds == 4'hb; // @[InvCipher.scala 73:32]
  AddRoundKey AddRoundKeyModule ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKeyModule_io_state_in_0),
    .io_state_in_1(AddRoundKeyModule_io_state_in_1),
    .io_state_in_2(AddRoundKeyModule_io_state_in_2),
    .io_state_in_3(AddRoundKeyModule_io_state_in_3),
    .io_state_in_4(AddRoundKeyModule_io_state_in_4),
    .io_state_in_5(AddRoundKeyModule_io_state_in_5),
    .io_state_in_6(AddRoundKeyModule_io_state_in_6),
    .io_state_in_7(AddRoundKeyModule_io_state_in_7),
    .io_state_in_8(AddRoundKeyModule_io_state_in_8),
    .io_state_in_9(AddRoundKeyModule_io_state_in_9),
    .io_state_in_10(AddRoundKeyModule_io_state_in_10),
    .io_state_in_11(AddRoundKeyModule_io_state_in_11),
    .io_state_in_12(AddRoundKeyModule_io_state_in_12),
    .io_state_in_13(AddRoundKeyModule_io_state_in_13),
    .io_state_in_14(AddRoundKeyModule_io_state_in_14),
    .io_state_in_15(AddRoundKeyModule_io_state_in_15),
    .io_roundKey_0(AddRoundKeyModule_io_roundKey_0),
    .io_roundKey_1(AddRoundKeyModule_io_roundKey_1),
    .io_roundKey_2(AddRoundKeyModule_io_roundKey_2),
    .io_roundKey_3(AddRoundKeyModule_io_roundKey_3),
    .io_roundKey_4(AddRoundKeyModule_io_roundKey_4),
    .io_roundKey_5(AddRoundKeyModule_io_roundKey_5),
    .io_roundKey_6(AddRoundKeyModule_io_roundKey_6),
    .io_roundKey_7(AddRoundKeyModule_io_roundKey_7),
    .io_roundKey_8(AddRoundKeyModule_io_roundKey_8),
    .io_roundKey_9(AddRoundKeyModule_io_roundKey_9),
    .io_roundKey_10(AddRoundKeyModule_io_roundKey_10),
    .io_roundKey_11(AddRoundKeyModule_io_roundKey_11),
    .io_roundKey_12(AddRoundKeyModule_io_roundKey_12),
    .io_roundKey_13(AddRoundKeyModule_io_roundKey_13),
    .io_roundKey_14(AddRoundKeyModule_io_roundKey_14),
    .io_roundKey_15(AddRoundKeyModule_io_roundKey_15),
    .io_state_out_0(AddRoundKeyModule_io_state_out_0),
    .io_state_out_1(AddRoundKeyModule_io_state_out_1),
    .io_state_out_2(AddRoundKeyModule_io_state_out_2),
    .io_state_out_3(AddRoundKeyModule_io_state_out_3),
    .io_state_out_4(AddRoundKeyModule_io_state_out_4),
    .io_state_out_5(AddRoundKeyModule_io_state_out_5),
    .io_state_out_6(AddRoundKeyModule_io_state_out_6),
    .io_state_out_7(AddRoundKeyModule_io_state_out_7),
    .io_state_out_8(AddRoundKeyModule_io_state_out_8),
    .io_state_out_9(AddRoundKeyModule_io_state_out_9),
    .io_state_out_10(AddRoundKeyModule_io_state_out_10),
    .io_state_out_11(AddRoundKeyModule_io_state_out_11),
    .io_state_out_12(AddRoundKeyModule_io_state_out_12),
    .io_state_out_13(AddRoundKeyModule_io_state_out_13),
    .io_state_out_14(AddRoundKeyModule_io_state_out_14),
    .io_state_out_15(AddRoundKeyModule_io_state_out_15)
  );
  InvSubBytes InvSubBytesModule ( // @[InvSubBytes.scala 43:84]
    .io_state_in_0(InvSubBytesModule_io_state_in_0),
    .io_state_in_1(InvSubBytesModule_io_state_in_1),
    .io_state_in_2(InvSubBytesModule_io_state_in_2),
    .io_state_in_3(InvSubBytesModule_io_state_in_3),
    .io_state_in_4(InvSubBytesModule_io_state_in_4),
    .io_state_in_5(InvSubBytesModule_io_state_in_5),
    .io_state_in_6(InvSubBytesModule_io_state_in_6),
    .io_state_in_7(InvSubBytesModule_io_state_in_7),
    .io_state_in_8(InvSubBytesModule_io_state_in_8),
    .io_state_in_9(InvSubBytesModule_io_state_in_9),
    .io_state_in_10(InvSubBytesModule_io_state_in_10),
    .io_state_in_11(InvSubBytesModule_io_state_in_11),
    .io_state_in_12(InvSubBytesModule_io_state_in_12),
    .io_state_in_13(InvSubBytesModule_io_state_in_13),
    .io_state_in_14(InvSubBytesModule_io_state_in_14),
    .io_state_in_15(InvSubBytesModule_io_state_in_15),
    .io_state_out_0(InvSubBytesModule_io_state_out_0),
    .io_state_out_1(InvSubBytesModule_io_state_out_1),
    .io_state_out_2(InvSubBytesModule_io_state_out_2),
    .io_state_out_3(InvSubBytesModule_io_state_out_3),
    .io_state_out_4(InvSubBytesModule_io_state_out_4),
    .io_state_out_5(InvSubBytesModule_io_state_out_5),
    .io_state_out_6(InvSubBytesModule_io_state_out_6),
    .io_state_out_7(InvSubBytesModule_io_state_out_7),
    .io_state_out_8(InvSubBytesModule_io_state_out_8),
    .io_state_out_9(InvSubBytesModule_io_state_out_9),
    .io_state_out_10(InvSubBytesModule_io_state_out_10),
    .io_state_out_11(InvSubBytesModule_io_state_out_11),
    .io_state_out_12(InvSubBytesModule_io_state_out_12),
    .io_state_out_13(InvSubBytesModule_io_state_out_13),
    .io_state_out_14(InvSubBytesModule_io_state_out_14),
    .io_state_out_15(InvSubBytesModule_io_state_out_15)
  );
  InvShiftRows InvShiftRowsModule ( // @[InvShiftRows.scala 35:37]
    .io_state_in_0(InvShiftRowsModule_io_state_in_0),
    .io_state_in_1(InvShiftRowsModule_io_state_in_1),
    .io_state_in_2(InvShiftRowsModule_io_state_in_2),
    .io_state_in_3(InvShiftRowsModule_io_state_in_3),
    .io_state_in_4(InvShiftRowsModule_io_state_in_4),
    .io_state_in_5(InvShiftRowsModule_io_state_in_5),
    .io_state_in_6(InvShiftRowsModule_io_state_in_6),
    .io_state_in_7(InvShiftRowsModule_io_state_in_7),
    .io_state_in_8(InvShiftRowsModule_io_state_in_8),
    .io_state_in_9(InvShiftRowsModule_io_state_in_9),
    .io_state_in_10(InvShiftRowsModule_io_state_in_10),
    .io_state_in_11(InvShiftRowsModule_io_state_in_11),
    .io_state_in_12(InvShiftRowsModule_io_state_in_12),
    .io_state_in_13(InvShiftRowsModule_io_state_in_13),
    .io_state_in_14(InvShiftRowsModule_io_state_in_14),
    .io_state_in_15(InvShiftRowsModule_io_state_in_15),
    .io_state_out_0(InvShiftRowsModule_io_state_out_0),
    .io_state_out_1(InvShiftRowsModule_io_state_out_1),
    .io_state_out_2(InvShiftRowsModule_io_state_out_2),
    .io_state_out_3(InvShiftRowsModule_io_state_out_3),
    .io_state_out_4(InvShiftRowsModule_io_state_out_4),
    .io_state_out_5(InvShiftRowsModule_io_state_out_5),
    .io_state_out_6(InvShiftRowsModule_io_state_out_6),
    .io_state_out_7(InvShiftRowsModule_io_state_out_7),
    .io_state_out_8(InvShiftRowsModule_io_state_out_8),
    .io_state_out_9(InvShiftRowsModule_io_state_out_9),
    .io_state_out_10(InvShiftRowsModule_io_state_out_10),
    .io_state_out_11(InvShiftRowsModule_io_state_out_11),
    .io_state_out_12(InvShiftRowsModule_io_state_out_12),
    .io_state_out_13(InvShiftRowsModule_io_state_out_13),
    .io_state_out_14(InvShiftRowsModule_io_state_out_14),
    .io_state_out_15(InvShiftRowsModule_io_state_out_15)
  );
  InvMixColumns InvMixColumnsModule ( // @[InvMixColumns.scala 154:64]
    .io_state_in_0(InvMixColumnsModule_io_state_in_0),
    .io_state_in_1(InvMixColumnsModule_io_state_in_1),
    .io_state_in_2(InvMixColumnsModule_io_state_in_2),
    .io_state_in_3(InvMixColumnsModule_io_state_in_3),
    .io_state_in_4(InvMixColumnsModule_io_state_in_4),
    .io_state_in_5(InvMixColumnsModule_io_state_in_5),
    .io_state_in_6(InvMixColumnsModule_io_state_in_6),
    .io_state_in_7(InvMixColumnsModule_io_state_in_7),
    .io_state_in_8(InvMixColumnsModule_io_state_in_8),
    .io_state_in_9(InvMixColumnsModule_io_state_in_9),
    .io_state_in_10(InvMixColumnsModule_io_state_in_10),
    .io_state_in_11(InvMixColumnsModule_io_state_in_11),
    .io_state_in_12(InvMixColumnsModule_io_state_in_12),
    .io_state_in_13(InvMixColumnsModule_io_state_in_13),
    .io_state_in_14(InvMixColumnsModule_io_state_in_14),
    .io_state_in_15(InvMixColumnsModule_io_state_in_15),
    .io_state_out_0(InvMixColumnsModule_io_state_out_0),
    .io_state_out_1(InvMixColumnsModule_io_state_out_1),
    .io_state_out_2(InvMixColumnsModule_io_state_out_2),
    .io_state_out_3(InvMixColumnsModule_io_state_out_3),
    .io_state_out_4(InvMixColumnsModule_io_state_out_4),
    .io_state_out_5(InvMixColumnsModule_io_state_out_5),
    .io_state_out_6(InvMixColumnsModule_io_state_out_6),
    .io_state_out_7(InvMixColumnsModule_io_state_out_7),
    .io_state_out_8(InvMixColumnsModule_io_state_out_8),
    .io_state_out_9(InvMixColumnsModule_io_state_out_9),
    .io_state_out_10(InvMixColumnsModule_io_state_out_10),
    .io_state_out_11(InvMixColumnsModule_io_state_out_11),
    .io_state_out_12(InvMixColumnsModule_io_state_out_12),
    .io_state_out_13(InvMixColumnsModule_io_state_out_13),
    .io_state_out_14(InvMixColumnsModule_io_state_out_14),
    .io_state_out_15(InvMixColumnsModule_io_state_out_15)
  );
  assign io_state_out_0 = _io_state_out_valid_T ? state_0 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_1 = _io_state_out_valid_T ? state_1 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_2 = _io_state_out_valid_T ? state_2 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_3 = _io_state_out_valid_T ? state_3 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_4 = _io_state_out_valid_T ? state_4 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_5 = _io_state_out_valid_T ? state_5 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_6 = _io_state_out_valid_T ? state_6 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_7 = _io_state_out_valid_T ? state_7 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_8 = _io_state_out_valid_T ? state_8 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_9 = _io_state_out_valid_T ? state_9 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_10 = _io_state_out_valid_T ? state_10 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_11 = _io_state_out_valid_T ? state_11 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_12 = _io_state_out_valid_T ? state_12 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_13 = _io_state_out_valid_T ? state_13 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_14 = _io_state_out_valid_T ? state_14 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_15 = _io_state_out_valid_T ? state_15 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_valid = rounds == 4'hb; // @[InvCipher.scala 73:32]
  assign AddRoundKeyModule_io_state_in_0 = STM == 2'h1 ? io_ciphertext_0 : InvSubBytesModule_io_state_out_0; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_1 = STM == 2'h1 ? io_ciphertext_1 : InvSubBytesModule_io_state_out_1; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_2 = STM == 2'h1 ? io_ciphertext_2 : InvSubBytesModule_io_state_out_2; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_3 = STM == 2'h1 ? io_ciphertext_3 : InvSubBytesModule_io_state_out_3; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_4 = STM == 2'h1 ? io_ciphertext_4 : InvSubBytesModule_io_state_out_4; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_5 = STM == 2'h1 ? io_ciphertext_5 : InvSubBytesModule_io_state_out_5; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_6 = STM == 2'h1 ? io_ciphertext_6 : InvSubBytesModule_io_state_out_6; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_7 = STM == 2'h1 ? io_ciphertext_7 : InvSubBytesModule_io_state_out_7; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_8 = STM == 2'h1 ? io_ciphertext_8 : InvSubBytesModule_io_state_out_8; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_9 = STM == 2'h1 ? io_ciphertext_9 : InvSubBytesModule_io_state_out_9; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_10 = STM == 2'h1 ? io_ciphertext_10 : InvSubBytesModule_io_state_out_10; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_11 = STM == 2'h1 ? io_ciphertext_11 : InvSubBytesModule_io_state_out_11; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_12 = STM == 2'h1 ? io_ciphertext_12 : InvSubBytesModule_io_state_out_12; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_13 = STM == 2'h1 ? io_ciphertext_13 : InvSubBytesModule_io_state_out_13; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_14 = STM == 2'h1 ? io_ciphertext_14 : InvSubBytesModule_io_state_out_14; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_15 = STM == 2'h1 ? io_ciphertext_15 : InvSubBytesModule_io_state_out_15; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_roundKey_0 = io_roundKey_0; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_1 = io_roundKey_1; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_2 = io_roundKey_2; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_3 = io_roundKey_3; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_4 = io_roundKey_4; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_5 = io_roundKey_5; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_6 = io_roundKey_6; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_7 = io_roundKey_7; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_8 = io_roundKey_8; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_9 = io_roundKey_9; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_10 = io_roundKey_10; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_11 = io_roundKey_11; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_12 = io_roundKey_12; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_13 = io_roundKey_13; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_14 = io_roundKey_14; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_15 = io_roundKey_15; // @[InvCipher.scala 65:33]
  assign InvSubBytesModule_io_state_in_0 = InvShiftRowsModule_io_state_out_0; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_1 = InvShiftRowsModule_io_state_out_1; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_2 = InvShiftRowsModule_io_state_out_2; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_3 = InvShiftRowsModule_io_state_out_3; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_4 = InvShiftRowsModule_io_state_out_4; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_5 = InvShiftRowsModule_io_state_out_5; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_6 = InvShiftRowsModule_io_state_out_6; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_7 = InvShiftRowsModule_io_state_out_7; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_8 = InvShiftRowsModule_io_state_out_8; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_9 = InvShiftRowsModule_io_state_out_9; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_10 = InvShiftRowsModule_io_state_out_10; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_11 = InvShiftRowsModule_io_state_out_11; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_12 = InvShiftRowsModule_io_state_out_12; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_13 = InvShiftRowsModule_io_state_out_13; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_14 = InvShiftRowsModule_io_state_out_14; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_15 = InvShiftRowsModule_io_state_out_15; // @[InvCipher.scala 61:33]
  assign InvShiftRowsModule_io_state_in_0 = state_0; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_1 = state_1; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_2 = state_2; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_3 = state_3; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_4 = state_4; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_5 = state_5; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_6 = state_6; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_7 = state_7; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_8 = state_8; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_9 = state_9; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_10 = state_10; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_11 = state_11; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_12 = state_12; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_13 = state_13; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_14 = state_14; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_15 = state_15; // @[InvCipher.scala 58:34]
  assign InvMixColumnsModule_io_state_in_0 = AddRoundKeyModule_io_state_out_0; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_1 = AddRoundKeyModule_io_state_out_1; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_2 = AddRoundKeyModule_io_state_out_2; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_3 = AddRoundKeyModule_io_state_out_3; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_4 = AddRoundKeyModule_io_state_out_4; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_5 = AddRoundKeyModule_io_state_out_5; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_6 = AddRoundKeyModule_io_state_out_6; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_7 = AddRoundKeyModule_io_state_out_7; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_8 = AddRoundKeyModule_io_state_out_8; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_9 = AddRoundKeyModule_io_state_out_9; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_10 = AddRoundKeyModule_io_state_out_10; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_11 = AddRoundKeyModule_io_state_out_11; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_12 = AddRoundKeyModule_io_state_out_12; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_13 = AddRoundKeyModule_io_state_out_13; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_14 = AddRoundKeyModule_io_state_out_14; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_15 = AddRoundKeyModule_io_state_out_15; // @[InvCipher.scala 68:35]
  always @(posedge clock) begin
    if (reset) begin // @[InvCipher.scala 31:22]
      state_0 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_0 <= InvMixColumnsModule_io_state_out_0;
      end else begin
        state_0 <= AddRoundKeyModule_io_state_out_0;
      end
    end else begin
      state_0 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_1 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_1 <= InvMixColumnsModule_io_state_out_1;
      end else begin
        state_1 <= AddRoundKeyModule_io_state_out_1;
      end
    end else begin
      state_1 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_2 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_2 <= InvMixColumnsModule_io_state_out_2;
      end else begin
        state_2 <= AddRoundKeyModule_io_state_out_2;
      end
    end else begin
      state_2 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_3 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_3 <= InvMixColumnsModule_io_state_out_3;
      end else begin
        state_3 <= AddRoundKeyModule_io_state_out_3;
      end
    end else begin
      state_3 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_4 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_4 <= InvMixColumnsModule_io_state_out_4;
      end else begin
        state_4 <= AddRoundKeyModule_io_state_out_4;
      end
    end else begin
      state_4 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_5 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_5 <= InvMixColumnsModule_io_state_out_5;
      end else begin
        state_5 <= AddRoundKeyModule_io_state_out_5;
      end
    end else begin
      state_5 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_6 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_6 <= InvMixColumnsModule_io_state_out_6;
      end else begin
        state_6 <= AddRoundKeyModule_io_state_out_6;
      end
    end else begin
      state_6 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_7 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_7 <= InvMixColumnsModule_io_state_out_7;
      end else begin
        state_7 <= AddRoundKeyModule_io_state_out_7;
      end
    end else begin
      state_7 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_8 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_8 <= InvMixColumnsModule_io_state_out_8;
      end else begin
        state_8 <= AddRoundKeyModule_io_state_out_8;
      end
    end else begin
      state_8 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_9 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_9 <= InvMixColumnsModule_io_state_out_9;
      end else begin
        state_9 <= AddRoundKeyModule_io_state_out_9;
      end
    end else begin
      state_9 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_10 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_10 <= InvMixColumnsModule_io_state_out_10;
      end else begin
        state_10 <= AddRoundKeyModule_io_state_out_10;
      end
    end else begin
      state_10 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_11 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_11 <= InvMixColumnsModule_io_state_out_11;
      end else begin
        state_11 <= AddRoundKeyModule_io_state_out_11;
      end
    end else begin
      state_11 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_12 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_12 <= InvMixColumnsModule_io_state_out_12;
      end else begin
        state_12 <= AddRoundKeyModule_io_state_out_12;
      end
    end else begin
      state_12 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_13 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_13 <= InvMixColumnsModule_io_state_out_13;
      end else begin
        state_13 <= AddRoundKeyModule_io_state_out_13;
      end
    end else begin
      state_13 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_14 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_14 <= InvMixColumnsModule_io_state_out_14;
      end else begin
        state_14 <= AddRoundKeyModule_io_state_out_14;
      end
    end else begin
      state_14 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_15 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_15 <= InvMixColumnsModule_io_state_out_15;
      end else begin
        state_15 <= AddRoundKeyModule_io_state_out_15;
      end
    end else begin
      state_15 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 32:23]
      rounds <= 4'h0; // @[InvCipher.scala 32:23]
    end else if (2'h0 == STM) begin // @[InvCipher.scala 38:15]
      rounds <= 4'h0; // @[InvCipher.scala 43:14]
    end else if (2'h1 == STM) begin // @[InvCipher.scala 38:15]
      rounds <= _rounds_T_1; // @[InvCipher.scala 46:14]
    end else if (2'h2 == STM) begin // @[InvCipher.scala 38:15]
      rounds <= _rounds_T_1; // @[InvCipher.scala 50:14]
    end
    if (reset) begin // @[InvCipher.scala 36:20]
      STM <= 2'h0; // @[InvCipher.scala 36:20]
    end else if (2'h0 == STM) begin // @[InvCipher.scala 38:15]
      if (io_start) begin // @[InvCipher.scala 40:22]
        STM <= 2'h1; // @[InvCipher.scala 41:13]
      end
    end else if (2'h1 == STM) begin // @[InvCipher.scala 38:15]
      STM <= 2'h2; // @[InvCipher.scala 47:11]
    end else if (2'h2 == STM) begin // @[InvCipher.scala 38:15]
      STM <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  rounds = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  STM = _RAND_17[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AESDecrypt(
  input          clock,
  input          reset,
  input          io_input_valid,
  input  [255:0] io_input_text,
  output [255:0] io_output_text,
  output         io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  invcipher_A_clock; // @[InvCipher.scala 101:78]
  wire  invcipher_A_reset; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_15; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_15; // @[InvCipher.scala 101:78]
  wire  invcipher_A_io_start; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_15; // @[InvCipher.scala 101:78]
  wire  invcipher_A_io_state_out_valid; // @[InvCipher.scala 101:78]
  wire  invcipher_B_clock; // @[InvCipher.scala 101:78]
  wire  invcipher_B_reset; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_15; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_15; // @[InvCipher.scala 101:78]
  wire  invcipher_B_io_start; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_15; // @[InvCipher.scala 101:78]
  wire  invcipher_B_io_state_out_valid; // @[InvCipher.scala 101:78]
  reg [3:0] address; // @[AESDecrypt.scala 95:26]
  reg  tmp; // @[AESDecrypt.scala 97:22]
  wire [3:0] _address_T_1 = address - 4'h1; // @[AESDecrypt.scala 102:26]
  wire  _GEN_2 = io_input_valid & ~tmp | tmp; // @[AESDecrypt.scala 100:15 97:22 98:34]
  wire [7:0] _GEN_4 = 4'h1 == address ? 8'hd6 : 8'h0; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_5 = 4'h2 == address ? 8'hb6 : _GEN_4; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_6 = 4'h3 == address ? 8'hb6 : _GEN_5; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_7 = 4'h4 == address ? 8'h47 : _GEN_6; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_8 = 4'h5 == address ? 8'h3c : _GEN_7; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_9 = 4'h6 == address ? 8'h5e : _GEN_8; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_10 = 4'h7 == address ? 8'h14 : _GEN_9; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_11 = 4'h8 == address ? 8'h47 : _GEN_10; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_12 = 4'h9 == address ? 8'h54 : _GEN_11; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_15 = 4'h1 == address ? 8'haa : 8'h1; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_16 = 4'h2 == address ? 8'h92 : _GEN_15; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_17 = 4'h3 == address ? 8'hff : _GEN_16; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_18 = 4'h4 == address ? 8'hf7 : _GEN_17; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_19 = 4'h5 == address ? 8'haa : _GEN_18; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_20 = 4'h6 == address ? 8'h39 : _GEN_19; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_21 = 4'h7 == address ? 8'hf9 : _GEN_20; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_22 = 4'h8 == address ? 8'h43 : _GEN_21; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_23 = 4'h9 == address ? 8'h99 : _GEN_22; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_26 = 4'h1 == address ? 8'h74 : 8'h2; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_27 = 4'h2 == address ? 8'hcf : _GEN_26; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_28 = 4'h3 == address ? 8'h74 : _GEN_27; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_29 = 4'h4 == address ? 8'hf7 : _GEN_28; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_30 = 4'h5 == address ? 8'ha3 : _GEN_29; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_31 = 4'h6 == address ? 8'hf : _GEN_30; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_32 = 4'h7 == address ? 8'h70 : _GEN_31; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_33 = 4'h8 == address ? 8'h87 : _GEN_32; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_34 = 4'h9 == address ? 8'h32 : _GEN_33; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_37 = 4'h1 == address ? 8'hfd : 8'h3; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_38 = 4'h2 == address ? 8'hb : _GEN_37; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_39 = 4'h3 == address ? 8'h4e : _GEN_38; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_40 = 4'h4 == address ? 8'hbc : _GEN_39; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_41 = 4'h5 == address ? 8'he8 : _GEN_40; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_42 = 4'h6 == address ? 8'h7d : _GEN_41; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_43 = 4'h7 == address ? 8'h1a : _GEN_42; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_44 = 4'h8 == address ? 8'h35 : _GEN_43; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_45 = 4'h9 == address ? 8'hd1 : _GEN_44; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_48 = 4'h1 == address ? 8'hd2 : 8'h4; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_49 = 4'h2 == address ? 8'h64 : _GEN_48; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_50 = 4'h3 == address ? 8'hd2 : _GEN_49; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_51 = 4'h4 == address ? 8'h95 : _GEN_50; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_52 = 4'h5 == address ? 8'ha9 : _GEN_51; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_53 = 4'h6 == address ? 8'hf7 : _GEN_52; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_54 = 4'h7 == address ? 8'he3 : _GEN_53; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_55 = 4'h8 == address ? 8'ha4 : _GEN_54; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_56 = 4'h9 == address ? 8'hf0 : _GEN_55; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_59 = 4'h1 == address ? 8'haf : 8'h5; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_60 = 4'h2 == address ? 8'h3d : _GEN_59; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_61 = 4'h3 == address ? 8'hc2 : _GEN_60; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_62 = 4'h4 == address ? 8'h35 : _GEN_61; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_63 = 4'h5 == address ? 8'h9f : _GEN_62; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_64 = 4'h6 == address ? 8'ha6 : _GEN_63; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_65 = 4'h7 == address ? 8'h5f : _GEN_64; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_66 = 4'h8 == address ? 8'h1c : _GEN_65; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_67 = 4'h9 == address ? 8'h85 : _GEN_66; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_70 = 4'h1 == address ? 8'h72 : 8'h6; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_71 = 4'h2 == address ? 8'hbd : _GEN_70; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_72 = 4'h3 == address ? 8'hc9 : _GEN_71; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_73 = 4'h4 == address ? 8'h3e : _GEN_72; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_74 = 4'h5 == address ? 8'h9d : _GEN_73; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_75 = 4'h6 == address ? 8'h92 : _GEN_74; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_76 = 4'h7 == address ? 8'he2 : _GEN_75; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_77 = 4'h8 == address ? 8'h65 : _GEN_76; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_78 = 4'h9 == address ? 8'h57 : _GEN_77; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_81 = 4'h1 == address ? 8'hfa : 8'h7; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_82 = 4'h2 == address ? 8'hf1 : _GEN_81; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_83 = 4'h3 == address ? 8'hbf : _GEN_82; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_84 = 4'h4 == address ? 8'h3 : _GEN_83; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_85 = 4'h5 == address ? 8'heb : _GEN_84; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_86 = 4'h6 == address ? 8'h96 : _GEN_85; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_87 = 4'h7 == address ? 8'h8c : _GEN_86; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_88 = 4'h8 == address ? 8'hb9 : _GEN_87; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_89 = 4'h9 == address ? 8'h68 : _GEN_88; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_92 = 4'h1 == address ? 8'hda : 8'h8; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_93 = 4'h2 == address ? 8'hbe : _GEN_92; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_94 = 4'h3 == address ? 8'h6c : _GEN_93; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_95 = 4'h4 == address ? 8'hf9 : _GEN_94; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_96 = 4'h5 == address ? 8'h50 : _GEN_95; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_97 = 4'h6 == address ? 8'ha7 : _GEN_96; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_98 = 4'h7 == address ? 8'h44 : _GEN_97; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_99 = 4'h8 == address ? 8'he0 : _GEN_98; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_100 = 4'h9 == address ? 8'h10 : _GEN_99; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_103 = 4'h1 == address ? 8'ha6 : 8'h9; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_104 = 4'h2 == address ? 8'h9b : _GEN_103; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_105 = 4'h3 == address ? 8'h59 : _GEN_104; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_106 = 4'h4 == address ? 8'h6c : _GEN_105; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_107 = 4'h5 == address ? 8'hf3 : _GEN_106; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_108 = 4'h6 == address ? 8'h55 : _GEN_107; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_109 = 4'h7 == address ? 8'ha : _GEN_108; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_110 = 4'h8 == address ? 8'h16 : _GEN_109; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_111 = 4'h9 == address ? 8'h93 : _GEN_110; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_114 = 4'h1 == address ? 8'h78 : 8'ha; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_115 = 4'h2 == address ? 8'hc5 : _GEN_114; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_116 = 4'h3 == address ? 8'hc : _GEN_115; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_117 = 4'h4 == address ? 8'h32 : _GEN_116; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_118 = 4'h5 == address ? 8'haf : _GEN_117; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_119 = 4'h6 == address ? 8'h3d : _GEN_118; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_120 = 4'h7 == address ? 8'hdf : _GEN_119; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_121 = 4'h8 == address ? 8'hba : _GEN_120; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_122 = 4'h9 == address ? 8'hed : _GEN_121; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_125 = 4'h1 == address ? 8'hf1 : 8'hb; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_126 = 4'h2 == address ? 8'h0 : _GEN_125; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_127 = 4'h3 == address ? 8'hbf : _GEN_126; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_128 = 4'h4 == address ? 8'hbc : _GEN_127; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_129 = 4'h5 == address ? 8'h57 : _GEN_128; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_130 = 4'h6 == address ? 8'hc1 : _GEN_129; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_131 = 4'h7 == address ? 8'h4d : _GEN_130; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_132 = 4'h8 == address ? 8'hf4 : _GEN_131; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_133 = 4'h9 == address ? 8'h9c : _GEN_132; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_136 = 4'h1 == address ? 8'hd6 : 8'hc; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_137 = 4'h2 == address ? 8'h68 : _GEN_136; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_138 = 4'h3 == address ? 8'h4 : _GEN_137; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_139 = 4'h4 == address ? 8'hfd : _GEN_138; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_140 = 4'h5 == address ? 8'had : _GEN_139; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_141 = 4'h6 == address ? 8'ha : _GEN_140; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_142 = 4'h7 == address ? 8'h4e : _GEN_141; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_143 = 4'h8 == address ? 8'hae : _GEN_142; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_144 = 4'h9 == address ? 8'hbe : _GEN_143; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_147 = 4'h1 == address ? 8'hab : 8'hd; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_148 = 4'h2 == address ? 8'h30 : _GEN_147; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_149 = 4'h3 == address ? 8'h69 : _GEN_148; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_150 = 4'h4 == address ? 8'h5 : _GEN_149; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_151 = 4'h5 == address ? 8'hf6 : _GEN_150; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_152 = 4'h6 == address ? 8'ha3 : _GEN_151; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_153 = 4'h7 == address ? 8'ha9 : _GEN_152; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_154 = 4'h8 == address ? 8'hbf : _GEN_153; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_155 = 4'h9 == address ? 8'h2c : _GEN_154; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_158 = 4'h1 == address ? 8'h76 : 8'he; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_159 = 4'h2 == address ? 8'hb3 : _GEN_158; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_160 = 4'h3 == address ? 8'hbf : _GEN_159; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_161 = 4'h4 == address ? 8'h8d : _GEN_160; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_162 = 4'h5 == address ? 8'h22 : _GEN_161; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_163 = 4'h6 == address ? 8'h1f : _GEN_162; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_164 = 4'h7 == address ? 8'hc0 : _GEN_163; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_165 = 4'h8 == address ? 8'h7a : _GEN_164; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_166 = 4'h9 == address ? 8'h97 : _GEN_165; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_169 = 4'h1 == address ? 8'hfe : 8'hf; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_170 = 4'h2 == address ? 8'hfe : _GEN_169; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_171 = 4'h3 == address ? 8'h41 : _GEN_170; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_172 = 4'h4 == address ? 8'hfd : _GEN_171; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_173 = 4'h5 == address ? 8'haa : _GEN_172; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_174 = 4'h6 == address ? 8'h6b : _GEN_173; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_175 = 4'h7 == address ? 8'h26 : _GEN_174; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_176 = 4'h8 == address ? 8'hd2 : _GEN_175; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_177 = 4'h9 == address ? 8'h4e : _GEN_176; // @[AESDecrypt.scala 106:{29,29}]
  wire [63:0] io_output_text_lo = {invcipher_A_io_state_out_8,invcipher_A_io_state_out_9,invcipher_A_io_state_out_10,
    invcipher_A_io_state_out_11,invcipher_A_io_state_out_12,invcipher_A_io_state_out_13,invcipher_A_io_state_out_14,
    invcipher_A_io_state_out_15}; // @[Cat.scala 31:58]
  wire [127:0] _io_output_text_T = {invcipher_A_io_state_out_0,invcipher_A_io_state_out_1,invcipher_A_io_state_out_2,
    invcipher_A_io_state_out_3,invcipher_A_io_state_out_4,invcipher_A_io_state_out_5,invcipher_A_io_state_out_6,
    invcipher_A_io_state_out_7,io_output_text_lo}; // @[Cat.scala 31:58]
  wire [63:0] io_output_text_lo_1 = {invcipher_B_io_state_out_8,invcipher_B_io_state_out_9,invcipher_B_io_state_out_10,
    invcipher_B_io_state_out_11,invcipher_B_io_state_out_12,invcipher_B_io_state_out_13,invcipher_B_io_state_out_14,
    invcipher_B_io_state_out_15}; // @[Cat.scala 31:58]
  wire [127:0] _io_output_text_T_1 = {invcipher_B_io_state_out_0,invcipher_B_io_state_out_1,invcipher_B_io_state_out_2,
    invcipher_B_io_state_out_3,invcipher_B_io_state_out_4,invcipher_B_io_state_out_5,invcipher_B_io_state_out_6,
    invcipher_B_io_state_out_7,io_output_text_lo_1}; // @[Cat.scala 31:58]
  InvCipher invcipher_A ( // @[InvCipher.scala 101:78]
    .clock(invcipher_A_clock),
    .reset(invcipher_A_reset),
    .io_ciphertext_0(invcipher_A_io_ciphertext_0),
    .io_ciphertext_1(invcipher_A_io_ciphertext_1),
    .io_ciphertext_2(invcipher_A_io_ciphertext_2),
    .io_ciphertext_3(invcipher_A_io_ciphertext_3),
    .io_ciphertext_4(invcipher_A_io_ciphertext_4),
    .io_ciphertext_5(invcipher_A_io_ciphertext_5),
    .io_ciphertext_6(invcipher_A_io_ciphertext_6),
    .io_ciphertext_7(invcipher_A_io_ciphertext_7),
    .io_ciphertext_8(invcipher_A_io_ciphertext_8),
    .io_ciphertext_9(invcipher_A_io_ciphertext_9),
    .io_ciphertext_10(invcipher_A_io_ciphertext_10),
    .io_ciphertext_11(invcipher_A_io_ciphertext_11),
    .io_ciphertext_12(invcipher_A_io_ciphertext_12),
    .io_ciphertext_13(invcipher_A_io_ciphertext_13),
    .io_ciphertext_14(invcipher_A_io_ciphertext_14),
    .io_ciphertext_15(invcipher_A_io_ciphertext_15),
    .io_roundKey_0(invcipher_A_io_roundKey_0),
    .io_roundKey_1(invcipher_A_io_roundKey_1),
    .io_roundKey_2(invcipher_A_io_roundKey_2),
    .io_roundKey_3(invcipher_A_io_roundKey_3),
    .io_roundKey_4(invcipher_A_io_roundKey_4),
    .io_roundKey_5(invcipher_A_io_roundKey_5),
    .io_roundKey_6(invcipher_A_io_roundKey_6),
    .io_roundKey_7(invcipher_A_io_roundKey_7),
    .io_roundKey_8(invcipher_A_io_roundKey_8),
    .io_roundKey_9(invcipher_A_io_roundKey_9),
    .io_roundKey_10(invcipher_A_io_roundKey_10),
    .io_roundKey_11(invcipher_A_io_roundKey_11),
    .io_roundKey_12(invcipher_A_io_roundKey_12),
    .io_roundKey_13(invcipher_A_io_roundKey_13),
    .io_roundKey_14(invcipher_A_io_roundKey_14),
    .io_roundKey_15(invcipher_A_io_roundKey_15),
    .io_start(invcipher_A_io_start),
    .io_state_out_0(invcipher_A_io_state_out_0),
    .io_state_out_1(invcipher_A_io_state_out_1),
    .io_state_out_2(invcipher_A_io_state_out_2),
    .io_state_out_3(invcipher_A_io_state_out_3),
    .io_state_out_4(invcipher_A_io_state_out_4),
    .io_state_out_5(invcipher_A_io_state_out_5),
    .io_state_out_6(invcipher_A_io_state_out_6),
    .io_state_out_7(invcipher_A_io_state_out_7),
    .io_state_out_8(invcipher_A_io_state_out_8),
    .io_state_out_9(invcipher_A_io_state_out_9),
    .io_state_out_10(invcipher_A_io_state_out_10),
    .io_state_out_11(invcipher_A_io_state_out_11),
    .io_state_out_12(invcipher_A_io_state_out_12),
    .io_state_out_13(invcipher_A_io_state_out_13),
    .io_state_out_14(invcipher_A_io_state_out_14),
    .io_state_out_15(invcipher_A_io_state_out_15),
    .io_state_out_valid(invcipher_A_io_state_out_valid)
  );
  InvCipher invcipher_B ( // @[InvCipher.scala 101:78]
    .clock(invcipher_B_clock),
    .reset(invcipher_B_reset),
    .io_ciphertext_0(invcipher_B_io_ciphertext_0),
    .io_ciphertext_1(invcipher_B_io_ciphertext_1),
    .io_ciphertext_2(invcipher_B_io_ciphertext_2),
    .io_ciphertext_3(invcipher_B_io_ciphertext_3),
    .io_ciphertext_4(invcipher_B_io_ciphertext_4),
    .io_ciphertext_5(invcipher_B_io_ciphertext_5),
    .io_ciphertext_6(invcipher_B_io_ciphertext_6),
    .io_ciphertext_7(invcipher_B_io_ciphertext_7),
    .io_ciphertext_8(invcipher_B_io_ciphertext_8),
    .io_ciphertext_9(invcipher_B_io_ciphertext_9),
    .io_ciphertext_10(invcipher_B_io_ciphertext_10),
    .io_ciphertext_11(invcipher_B_io_ciphertext_11),
    .io_ciphertext_12(invcipher_B_io_ciphertext_12),
    .io_ciphertext_13(invcipher_B_io_ciphertext_13),
    .io_ciphertext_14(invcipher_B_io_ciphertext_14),
    .io_ciphertext_15(invcipher_B_io_ciphertext_15),
    .io_roundKey_0(invcipher_B_io_roundKey_0),
    .io_roundKey_1(invcipher_B_io_roundKey_1),
    .io_roundKey_2(invcipher_B_io_roundKey_2),
    .io_roundKey_3(invcipher_B_io_roundKey_3),
    .io_roundKey_4(invcipher_B_io_roundKey_4),
    .io_roundKey_5(invcipher_B_io_roundKey_5),
    .io_roundKey_6(invcipher_B_io_roundKey_6),
    .io_roundKey_7(invcipher_B_io_roundKey_7),
    .io_roundKey_8(invcipher_B_io_roundKey_8),
    .io_roundKey_9(invcipher_B_io_roundKey_9),
    .io_roundKey_10(invcipher_B_io_roundKey_10),
    .io_roundKey_11(invcipher_B_io_roundKey_11),
    .io_roundKey_12(invcipher_B_io_roundKey_12),
    .io_roundKey_13(invcipher_B_io_roundKey_13),
    .io_roundKey_14(invcipher_B_io_roundKey_14),
    .io_roundKey_15(invcipher_B_io_roundKey_15),
    .io_start(invcipher_B_io_start),
    .io_state_out_0(invcipher_B_io_state_out_0),
    .io_state_out_1(invcipher_B_io_state_out_1),
    .io_state_out_2(invcipher_B_io_state_out_2),
    .io_state_out_3(invcipher_B_io_state_out_3),
    .io_state_out_4(invcipher_B_io_state_out_4),
    .io_state_out_5(invcipher_B_io_state_out_5),
    .io_state_out_6(invcipher_B_io_state_out_6),
    .io_state_out_7(invcipher_B_io_state_out_7),
    .io_state_out_8(invcipher_B_io_state_out_8),
    .io_state_out_9(invcipher_B_io_state_out_9),
    .io_state_out_10(invcipher_B_io_state_out_10),
    .io_state_out_11(invcipher_B_io_state_out_11),
    .io_state_out_12(invcipher_B_io_state_out_12),
    .io_state_out_13(invcipher_B_io_state_out_13),
    .io_state_out_14(invcipher_B_io_state_out_14),
    .io_state_out_15(invcipher_B_io_state_out_15),
    .io_state_out_valid(invcipher_B_io_state_out_valid)
  );
  assign io_output_text = {_io_output_text_T,_io_output_text_T_1}; // @[Cat.scala 31:58]
  assign io_output_valid = invcipher_A_io_state_out_valid & invcipher_B_io_state_out_valid; // @[AESDecrypt.scala 116:55]
  assign invcipher_A_clock = clock;
  assign invcipher_A_reset = reset;
  assign invcipher_A_io_ciphertext_0 = io_input_text[255:248]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_1 = io_input_text[247:240]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_2 = io_input_text[239:232]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_3 = io_input_text[231:224]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_4 = io_input_text[223:216]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_5 = io_input_text[215:208]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_6 = io_input_text[207:200]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_7 = io_input_text[199:192]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_8 = io_input_text[191:184]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_9 = io_input_text[183:176]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_10 = io_input_text[175:168]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_11 = io_input_text[167:160]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_12 = io_input_text[159:152]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_13 = io_input_text[151:144]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_14 = io_input_text[143:136]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_15 = io_input_text[135:128]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_start = io_input_valid; // @[AESDecrypt.scala 104:26]
  assign invcipher_B_clock = clock;
  assign invcipher_B_reset = reset;
  assign invcipher_B_io_ciphertext_0 = io_input_text[127:120]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_1 = io_input_text[119:112]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_2 = io_input_text[111:104]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_3 = io_input_text[103:96]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_4 = io_input_text[95:88]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_5 = io_input_text[87:80]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_6 = io_input_text[79:72]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_7 = io_input_text[71:64]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_8 = io_input_text[63:56]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_9 = io_input_text[55:48]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_10 = io_input_text[47:40]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_11 = io_input_text[39:32]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_12 = io_input_text[31:24]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_13 = io_input_text[23:16]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_14 = io_input_text[15:8]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_15 = io_input_text[7:0]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_start = io_input_valid; // @[AESDecrypt.scala 108:26]
  always @(posedge clock) begin
    if (reset) begin // @[AESDecrypt.scala 95:26]
      address <= 4'h0; // @[AESDecrypt.scala 95:26]
    end else if (io_input_valid & ~tmp) begin // @[AESDecrypt.scala 98:34]
      address <= 4'ha; // @[AESDecrypt.scala 99:15]
    end else if (address != 4'h0) begin // @[AESDecrypt.scala 101:32]
      address <= _address_T_1; // @[AESDecrypt.scala 102:15]
    end
    if (reset) begin // @[AESDecrypt.scala 97:22]
      tmp <= 1'h0; // @[AESDecrypt.scala 97:22]
    end else begin
      tmp <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  address = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  tmp = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InvCipher_2(
  input        clock,
  input        reset,
  input  [7:0] io_ciphertext_0,
  input  [7:0] io_ciphertext_1,
  input  [7:0] io_ciphertext_2,
  input  [7:0] io_ciphertext_3,
  input  [7:0] io_ciphertext_4,
  input  [7:0] io_ciphertext_5,
  input  [7:0] io_ciphertext_6,
  input  [7:0] io_ciphertext_7,
  input  [7:0] io_ciphertext_8,
  input  [7:0] io_ciphertext_9,
  input  [7:0] io_ciphertext_10,
  input  [7:0] io_ciphertext_11,
  input  [7:0] io_ciphertext_12,
  input  [7:0] io_ciphertext_13,
  input  [7:0] io_ciphertext_14,
  input  [7:0] io_ciphertext_15,
  input  [7:0] io_roundKey_0,
  input  [7:0] io_roundKey_1,
  input  [7:0] io_roundKey_2,
  input  [7:0] io_roundKey_3,
  input  [7:0] io_roundKey_4,
  input  [7:0] io_roundKey_5,
  input  [7:0] io_roundKey_6,
  input  [7:0] io_roundKey_7,
  input  [7:0] io_roundKey_8,
  input  [7:0] io_roundKey_9,
  input  [7:0] io_roundKey_10,
  input  [7:0] io_roundKey_11,
  input  [7:0] io_roundKey_12,
  input  [7:0] io_roundKey_13,
  input  [7:0] io_roundKey_14,
  input  [7:0] io_roundKey_15,
  input        io_start,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15,
  output       io_state_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] AddRoundKeyModule_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] InvSubBytesModule_io_state_in_0; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_1; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_2; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_3; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_4; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_5; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_6; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_7; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_8; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_9; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_10; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_11; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_12; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_13; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_14; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_in_15; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_0; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_1; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_2; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_3; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_4; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_5; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_6; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_7; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_8; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_9; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_10; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_11; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_12; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_13; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_14; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvSubBytesModule_io_state_out_15; // @[InvSubBytes.scala 43:84]
  wire [7:0] InvShiftRowsModule_io_state_in_0; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_1; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_2; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_3; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_4; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_5; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_6; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_7; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_8; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_9; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_10; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_11; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_12; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_13; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_14; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_in_15; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_0; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_1; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_2; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_3; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_4; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_5; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_6; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_7; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_8; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_9; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_10; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_11; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_12; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_13; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_14; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvShiftRowsModule_io_state_out_15; // @[InvShiftRows.scala 35:37]
  wire [7:0] InvMixColumnsModule_io_state_in_0; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_1; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_2; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_3; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_4; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_5; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_6; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_7; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_8; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_9; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_10; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_11; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_12; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_13; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_14; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_in_15; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_0; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_1; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_2; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_3; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_4; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_5; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_6; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_7; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_8; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_9; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_10; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_11; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_12; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_13; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_14; // @[InvMixColumns.scala 154:64]
  wire [7:0] InvMixColumnsModule_io_state_out_15; // @[InvMixColumns.scala 154:64]
  reg [7:0] state_0; // @[InvCipher.scala 31:22]
  reg [7:0] state_1; // @[InvCipher.scala 31:22]
  reg [7:0] state_2; // @[InvCipher.scala 31:22]
  reg [7:0] state_3; // @[InvCipher.scala 31:22]
  reg [7:0] state_4; // @[InvCipher.scala 31:22]
  reg [7:0] state_5; // @[InvCipher.scala 31:22]
  reg [7:0] state_6; // @[InvCipher.scala 31:22]
  reg [7:0] state_7; // @[InvCipher.scala 31:22]
  reg [7:0] state_8; // @[InvCipher.scala 31:22]
  reg [7:0] state_9; // @[InvCipher.scala 31:22]
  reg [7:0] state_10; // @[InvCipher.scala 31:22]
  reg [7:0] state_11; // @[InvCipher.scala 31:22]
  reg [7:0] state_12; // @[InvCipher.scala 31:22]
  reg [7:0] state_13; // @[InvCipher.scala 31:22]
  reg [7:0] state_14; // @[InvCipher.scala 31:22]
  reg [7:0] state_15; // @[InvCipher.scala 31:22]
  reg [3:0] rounds; // @[InvCipher.scala 32:23]
  reg [1:0] STM; // @[InvCipher.scala 36:20]
  wire [3:0] _rounds_T_1 = rounds + 4'h1; // @[InvCipher.scala 46:24]
  wire [1:0] _GEN_1 = rounds == 4'ha ? 2'h0 : STM; // @[InvCipher.scala 51:29 52:13 36:20]
  wire  _io_state_out_valid_T = rounds == 4'hb; // @[InvCipher.scala 73:32]
  AddRoundKey AddRoundKeyModule ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKeyModule_io_state_in_0),
    .io_state_in_1(AddRoundKeyModule_io_state_in_1),
    .io_state_in_2(AddRoundKeyModule_io_state_in_2),
    .io_state_in_3(AddRoundKeyModule_io_state_in_3),
    .io_state_in_4(AddRoundKeyModule_io_state_in_4),
    .io_state_in_5(AddRoundKeyModule_io_state_in_5),
    .io_state_in_6(AddRoundKeyModule_io_state_in_6),
    .io_state_in_7(AddRoundKeyModule_io_state_in_7),
    .io_state_in_8(AddRoundKeyModule_io_state_in_8),
    .io_state_in_9(AddRoundKeyModule_io_state_in_9),
    .io_state_in_10(AddRoundKeyModule_io_state_in_10),
    .io_state_in_11(AddRoundKeyModule_io_state_in_11),
    .io_state_in_12(AddRoundKeyModule_io_state_in_12),
    .io_state_in_13(AddRoundKeyModule_io_state_in_13),
    .io_state_in_14(AddRoundKeyModule_io_state_in_14),
    .io_state_in_15(AddRoundKeyModule_io_state_in_15),
    .io_roundKey_0(AddRoundKeyModule_io_roundKey_0),
    .io_roundKey_1(AddRoundKeyModule_io_roundKey_1),
    .io_roundKey_2(AddRoundKeyModule_io_roundKey_2),
    .io_roundKey_3(AddRoundKeyModule_io_roundKey_3),
    .io_roundKey_4(AddRoundKeyModule_io_roundKey_4),
    .io_roundKey_5(AddRoundKeyModule_io_roundKey_5),
    .io_roundKey_6(AddRoundKeyModule_io_roundKey_6),
    .io_roundKey_7(AddRoundKeyModule_io_roundKey_7),
    .io_roundKey_8(AddRoundKeyModule_io_roundKey_8),
    .io_roundKey_9(AddRoundKeyModule_io_roundKey_9),
    .io_roundKey_10(AddRoundKeyModule_io_roundKey_10),
    .io_roundKey_11(AddRoundKeyModule_io_roundKey_11),
    .io_roundKey_12(AddRoundKeyModule_io_roundKey_12),
    .io_roundKey_13(AddRoundKeyModule_io_roundKey_13),
    .io_roundKey_14(AddRoundKeyModule_io_roundKey_14),
    .io_roundKey_15(AddRoundKeyModule_io_roundKey_15),
    .io_state_out_0(AddRoundKeyModule_io_state_out_0),
    .io_state_out_1(AddRoundKeyModule_io_state_out_1),
    .io_state_out_2(AddRoundKeyModule_io_state_out_2),
    .io_state_out_3(AddRoundKeyModule_io_state_out_3),
    .io_state_out_4(AddRoundKeyModule_io_state_out_4),
    .io_state_out_5(AddRoundKeyModule_io_state_out_5),
    .io_state_out_6(AddRoundKeyModule_io_state_out_6),
    .io_state_out_7(AddRoundKeyModule_io_state_out_7),
    .io_state_out_8(AddRoundKeyModule_io_state_out_8),
    .io_state_out_9(AddRoundKeyModule_io_state_out_9),
    .io_state_out_10(AddRoundKeyModule_io_state_out_10),
    .io_state_out_11(AddRoundKeyModule_io_state_out_11),
    .io_state_out_12(AddRoundKeyModule_io_state_out_12),
    .io_state_out_13(AddRoundKeyModule_io_state_out_13),
    .io_state_out_14(AddRoundKeyModule_io_state_out_14),
    .io_state_out_15(AddRoundKeyModule_io_state_out_15)
  );
  InvSubBytes InvSubBytesModule ( // @[InvSubBytes.scala 43:84]
    .io_state_in_0(InvSubBytesModule_io_state_in_0),
    .io_state_in_1(InvSubBytesModule_io_state_in_1),
    .io_state_in_2(InvSubBytesModule_io_state_in_2),
    .io_state_in_3(InvSubBytesModule_io_state_in_3),
    .io_state_in_4(InvSubBytesModule_io_state_in_4),
    .io_state_in_5(InvSubBytesModule_io_state_in_5),
    .io_state_in_6(InvSubBytesModule_io_state_in_6),
    .io_state_in_7(InvSubBytesModule_io_state_in_7),
    .io_state_in_8(InvSubBytesModule_io_state_in_8),
    .io_state_in_9(InvSubBytesModule_io_state_in_9),
    .io_state_in_10(InvSubBytesModule_io_state_in_10),
    .io_state_in_11(InvSubBytesModule_io_state_in_11),
    .io_state_in_12(InvSubBytesModule_io_state_in_12),
    .io_state_in_13(InvSubBytesModule_io_state_in_13),
    .io_state_in_14(InvSubBytesModule_io_state_in_14),
    .io_state_in_15(InvSubBytesModule_io_state_in_15),
    .io_state_out_0(InvSubBytesModule_io_state_out_0),
    .io_state_out_1(InvSubBytesModule_io_state_out_1),
    .io_state_out_2(InvSubBytesModule_io_state_out_2),
    .io_state_out_3(InvSubBytesModule_io_state_out_3),
    .io_state_out_4(InvSubBytesModule_io_state_out_4),
    .io_state_out_5(InvSubBytesModule_io_state_out_5),
    .io_state_out_6(InvSubBytesModule_io_state_out_6),
    .io_state_out_7(InvSubBytesModule_io_state_out_7),
    .io_state_out_8(InvSubBytesModule_io_state_out_8),
    .io_state_out_9(InvSubBytesModule_io_state_out_9),
    .io_state_out_10(InvSubBytesModule_io_state_out_10),
    .io_state_out_11(InvSubBytesModule_io_state_out_11),
    .io_state_out_12(InvSubBytesModule_io_state_out_12),
    .io_state_out_13(InvSubBytesModule_io_state_out_13),
    .io_state_out_14(InvSubBytesModule_io_state_out_14),
    .io_state_out_15(InvSubBytesModule_io_state_out_15)
  );
  InvShiftRows InvShiftRowsModule ( // @[InvShiftRows.scala 35:37]
    .io_state_in_0(InvShiftRowsModule_io_state_in_0),
    .io_state_in_1(InvShiftRowsModule_io_state_in_1),
    .io_state_in_2(InvShiftRowsModule_io_state_in_2),
    .io_state_in_3(InvShiftRowsModule_io_state_in_3),
    .io_state_in_4(InvShiftRowsModule_io_state_in_4),
    .io_state_in_5(InvShiftRowsModule_io_state_in_5),
    .io_state_in_6(InvShiftRowsModule_io_state_in_6),
    .io_state_in_7(InvShiftRowsModule_io_state_in_7),
    .io_state_in_8(InvShiftRowsModule_io_state_in_8),
    .io_state_in_9(InvShiftRowsModule_io_state_in_9),
    .io_state_in_10(InvShiftRowsModule_io_state_in_10),
    .io_state_in_11(InvShiftRowsModule_io_state_in_11),
    .io_state_in_12(InvShiftRowsModule_io_state_in_12),
    .io_state_in_13(InvShiftRowsModule_io_state_in_13),
    .io_state_in_14(InvShiftRowsModule_io_state_in_14),
    .io_state_in_15(InvShiftRowsModule_io_state_in_15),
    .io_state_out_0(InvShiftRowsModule_io_state_out_0),
    .io_state_out_1(InvShiftRowsModule_io_state_out_1),
    .io_state_out_2(InvShiftRowsModule_io_state_out_2),
    .io_state_out_3(InvShiftRowsModule_io_state_out_3),
    .io_state_out_4(InvShiftRowsModule_io_state_out_4),
    .io_state_out_5(InvShiftRowsModule_io_state_out_5),
    .io_state_out_6(InvShiftRowsModule_io_state_out_6),
    .io_state_out_7(InvShiftRowsModule_io_state_out_7),
    .io_state_out_8(InvShiftRowsModule_io_state_out_8),
    .io_state_out_9(InvShiftRowsModule_io_state_out_9),
    .io_state_out_10(InvShiftRowsModule_io_state_out_10),
    .io_state_out_11(InvShiftRowsModule_io_state_out_11),
    .io_state_out_12(InvShiftRowsModule_io_state_out_12),
    .io_state_out_13(InvShiftRowsModule_io_state_out_13),
    .io_state_out_14(InvShiftRowsModule_io_state_out_14),
    .io_state_out_15(InvShiftRowsModule_io_state_out_15)
  );
  InvMixColumns InvMixColumnsModule ( // @[InvMixColumns.scala 154:64]
    .io_state_in_0(InvMixColumnsModule_io_state_in_0),
    .io_state_in_1(InvMixColumnsModule_io_state_in_1),
    .io_state_in_2(InvMixColumnsModule_io_state_in_2),
    .io_state_in_3(InvMixColumnsModule_io_state_in_3),
    .io_state_in_4(InvMixColumnsModule_io_state_in_4),
    .io_state_in_5(InvMixColumnsModule_io_state_in_5),
    .io_state_in_6(InvMixColumnsModule_io_state_in_6),
    .io_state_in_7(InvMixColumnsModule_io_state_in_7),
    .io_state_in_8(InvMixColumnsModule_io_state_in_8),
    .io_state_in_9(InvMixColumnsModule_io_state_in_9),
    .io_state_in_10(InvMixColumnsModule_io_state_in_10),
    .io_state_in_11(InvMixColumnsModule_io_state_in_11),
    .io_state_in_12(InvMixColumnsModule_io_state_in_12),
    .io_state_in_13(InvMixColumnsModule_io_state_in_13),
    .io_state_in_14(InvMixColumnsModule_io_state_in_14),
    .io_state_in_15(InvMixColumnsModule_io_state_in_15),
    .io_state_out_0(InvMixColumnsModule_io_state_out_0),
    .io_state_out_1(InvMixColumnsModule_io_state_out_1),
    .io_state_out_2(InvMixColumnsModule_io_state_out_2),
    .io_state_out_3(InvMixColumnsModule_io_state_out_3),
    .io_state_out_4(InvMixColumnsModule_io_state_out_4),
    .io_state_out_5(InvMixColumnsModule_io_state_out_5),
    .io_state_out_6(InvMixColumnsModule_io_state_out_6),
    .io_state_out_7(InvMixColumnsModule_io_state_out_7),
    .io_state_out_8(InvMixColumnsModule_io_state_out_8),
    .io_state_out_9(InvMixColumnsModule_io_state_out_9),
    .io_state_out_10(InvMixColumnsModule_io_state_out_10),
    .io_state_out_11(InvMixColumnsModule_io_state_out_11),
    .io_state_out_12(InvMixColumnsModule_io_state_out_12),
    .io_state_out_13(InvMixColumnsModule_io_state_out_13),
    .io_state_out_14(InvMixColumnsModule_io_state_out_14),
    .io_state_out_15(InvMixColumnsModule_io_state_out_15)
  );
  assign io_state_out_0 = _io_state_out_valid_T ? state_0 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_1 = _io_state_out_valid_T ? state_1 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_2 = _io_state_out_valid_T ? state_2 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_3 = _io_state_out_valid_T ? state_3 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_4 = _io_state_out_valid_T ? state_4 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_5 = _io_state_out_valid_T ? state_5 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_6 = _io_state_out_valid_T ? state_6 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_7 = _io_state_out_valid_T ? state_7 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_8 = _io_state_out_valid_T ? state_8 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_9 = _io_state_out_valid_T ? state_9 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_10 = _io_state_out_valid_T ? state_10 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_11 = _io_state_out_valid_T ? state_11 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_12 = _io_state_out_valid_T ? state_12 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_13 = _io_state_out_valid_T ? state_13 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_14 = _io_state_out_valid_T ? state_14 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_15 = _io_state_out_valid_T ? state_15 : 8'h0; // @[InvCipher.scala 74:22]
  assign io_state_out_valid = rounds == 4'hb; // @[InvCipher.scala 73:32]
  assign AddRoundKeyModule_io_state_in_0 = STM == 2'h1 ? io_ciphertext_0 : InvSubBytesModule_io_state_out_0; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_1 = STM == 2'h1 ? io_ciphertext_1 : InvSubBytesModule_io_state_out_1; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_2 = STM == 2'h1 ? io_ciphertext_2 : InvSubBytesModule_io_state_out_2; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_3 = STM == 2'h1 ? io_ciphertext_3 : InvSubBytesModule_io_state_out_3; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_4 = STM == 2'h1 ? io_ciphertext_4 : InvSubBytesModule_io_state_out_4; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_5 = STM == 2'h1 ? io_ciphertext_5 : InvSubBytesModule_io_state_out_5; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_6 = STM == 2'h1 ? io_ciphertext_6 : InvSubBytesModule_io_state_out_6; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_7 = STM == 2'h1 ? io_ciphertext_7 : InvSubBytesModule_io_state_out_7; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_8 = STM == 2'h1 ? io_ciphertext_8 : InvSubBytesModule_io_state_out_8; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_9 = STM == 2'h1 ? io_ciphertext_9 : InvSubBytesModule_io_state_out_9; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_10 = STM == 2'h1 ? io_ciphertext_10 : InvSubBytesModule_io_state_out_10; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_11 = STM == 2'h1 ? io_ciphertext_11 : InvSubBytesModule_io_state_out_11; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_12 = STM == 2'h1 ? io_ciphertext_12 : InvSubBytesModule_io_state_out_12; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_13 = STM == 2'h1 ? io_ciphertext_13 : InvSubBytesModule_io_state_out_13; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_14 = STM == 2'h1 ? io_ciphertext_14 : InvSubBytesModule_io_state_out_14; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_state_in_15 = STM == 2'h1 ? io_ciphertext_15 : InvSubBytesModule_io_state_out_15; // @[InvCipher.scala 64:39]
  assign AddRoundKeyModule_io_roundKey_0 = io_roundKey_0; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_1 = io_roundKey_1; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_2 = io_roundKey_2; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_3 = io_roundKey_3; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_4 = io_roundKey_4; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_5 = io_roundKey_5; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_6 = io_roundKey_6; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_7 = io_roundKey_7; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_8 = io_roundKey_8; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_9 = io_roundKey_9; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_10 = io_roundKey_10; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_11 = io_roundKey_11; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_12 = io_roundKey_12; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_13 = io_roundKey_13; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_14 = io_roundKey_14; // @[InvCipher.scala 65:33]
  assign AddRoundKeyModule_io_roundKey_15 = io_roundKey_15; // @[InvCipher.scala 65:33]
  assign InvSubBytesModule_io_state_in_0 = InvShiftRowsModule_io_state_out_0; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_1 = InvShiftRowsModule_io_state_out_1; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_2 = InvShiftRowsModule_io_state_out_2; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_3 = InvShiftRowsModule_io_state_out_3; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_4 = InvShiftRowsModule_io_state_out_4; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_5 = InvShiftRowsModule_io_state_out_5; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_6 = InvShiftRowsModule_io_state_out_6; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_7 = InvShiftRowsModule_io_state_out_7; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_8 = InvShiftRowsModule_io_state_out_8; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_9 = InvShiftRowsModule_io_state_out_9; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_10 = InvShiftRowsModule_io_state_out_10; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_11 = InvShiftRowsModule_io_state_out_11; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_12 = InvShiftRowsModule_io_state_out_12; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_13 = InvShiftRowsModule_io_state_out_13; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_14 = InvShiftRowsModule_io_state_out_14; // @[InvCipher.scala 61:33]
  assign InvSubBytesModule_io_state_in_15 = InvShiftRowsModule_io_state_out_15; // @[InvCipher.scala 61:33]
  assign InvShiftRowsModule_io_state_in_0 = state_0; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_1 = state_1; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_2 = state_2; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_3 = state_3; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_4 = state_4; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_5 = state_5; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_6 = state_6; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_7 = state_7; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_8 = state_8; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_9 = state_9; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_10 = state_10; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_11 = state_11; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_12 = state_12; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_13 = state_13; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_14 = state_14; // @[InvCipher.scala 58:34]
  assign InvShiftRowsModule_io_state_in_15 = state_15; // @[InvCipher.scala 58:34]
  assign InvMixColumnsModule_io_state_in_0 = AddRoundKeyModule_io_state_out_0; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_1 = AddRoundKeyModule_io_state_out_1; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_2 = AddRoundKeyModule_io_state_out_2; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_3 = AddRoundKeyModule_io_state_out_3; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_4 = AddRoundKeyModule_io_state_out_4; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_5 = AddRoundKeyModule_io_state_out_5; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_6 = AddRoundKeyModule_io_state_out_6; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_7 = AddRoundKeyModule_io_state_out_7; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_8 = AddRoundKeyModule_io_state_out_8; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_9 = AddRoundKeyModule_io_state_out_9; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_10 = AddRoundKeyModule_io_state_out_10; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_11 = AddRoundKeyModule_io_state_out_11; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_12 = AddRoundKeyModule_io_state_out_12; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_13 = AddRoundKeyModule_io_state_out_13; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_14 = AddRoundKeyModule_io_state_out_14; // @[InvCipher.scala 68:35]
  assign InvMixColumnsModule_io_state_in_15 = AddRoundKeyModule_io_state_out_15; // @[InvCipher.scala 68:35]
  always @(posedge clock) begin
    if (reset) begin // @[InvCipher.scala 31:22]
      state_0 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_0 <= InvMixColumnsModule_io_state_out_0;
      end else begin
        state_0 <= AddRoundKeyModule_io_state_out_0;
      end
    end else begin
      state_0 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_1 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_1 <= InvMixColumnsModule_io_state_out_1;
      end else begin
        state_1 <= AddRoundKeyModule_io_state_out_1;
      end
    end else begin
      state_1 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_2 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_2 <= InvMixColumnsModule_io_state_out_2;
      end else begin
        state_2 <= AddRoundKeyModule_io_state_out_2;
      end
    end else begin
      state_2 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_3 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_3 <= InvMixColumnsModule_io_state_out_3;
      end else begin
        state_3 <= AddRoundKeyModule_io_state_out_3;
      end
    end else begin
      state_3 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_4 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_4 <= InvMixColumnsModule_io_state_out_4;
      end else begin
        state_4 <= AddRoundKeyModule_io_state_out_4;
      end
    end else begin
      state_4 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_5 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_5 <= InvMixColumnsModule_io_state_out_5;
      end else begin
        state_5 <= AddRoundKeyModule_io_state_out_5;
      end
    end else begin
      state_5 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_6 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_6 <= InvMixColumnsModule_io_state_out_6;
      end else begin
        state_6 <= AddRoundKeyModule_io_state_out_6;
      end
    end else begin
      state_6 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_7 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_7 <= InvMixColumnsModule_io_state_out_7;
      end else begin
        state_7 <= AddRoundKeyModule_io_state_out_7;
      end
    end else begin
      state_7 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_8 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_8 <= InvMixColumnsModule_io_state_out_8;
      end else begin
        state_8 <= AddRoundKeyModule_io_state_out_8;
      end
    end else begin
      state_8 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_9 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_9 <= InvMixColumnsModule_io_state_out_9;
      end else begin
        state_9 <= AddRoundKeyModule_io_state_out_9;
      end
    end else begin
      state_9 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_10 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_10 <= InvMixColumnsModule_io_state_out_10;
      end else begin
        state_10 <= AddRoundKeyModule_io_state_out_10;
      end
    end else begin
      state_10 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_11 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_11 <= InvMixColumnsModule_io_state_out_11;
      end else begin
        state_11 <= AddRoundKeyModule_io_state_out_11;
      end
    end else begin
      state_11 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_12 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_12 <= InvMixColumnsModule_io_state_out_12;
      end else begin
        state_12 <= AddRoundKeyModule_io_state_out_12;
      end
    end else begin
      state_12 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_13 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_13 <= InvMixColumnsModule_io_state_out_13;
      end else begin
        state_13 <= AddRoundKeyModule_io_state_out_13;
      end
    end else begin
      state_13 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_14 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_14 <= InvMixColumnsModule_io_state_out_14;
      end else begin
        state_14 <= AddRoundKeyModule_io_state_out_14;
      end
    end else begin
      state_14 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 31:22]
      state_15 <= 8'h0; // @[InvCipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[InvCipher.scala 70:15]
      if (rounds > 4'h0 & rounds < 4'ha) begin // @[InvCipher.scala 70:34]
        state_15 <= InvMixColumnsModule_io_state_out_15;
      end else begin
        state_15 <= AddRoundKeyModule_io_state_out_15;
      end
    end else begin
      state_15 <= 8'h0;
    end
    if (reset) begin // @[InvCipher.scala 32:23]
      rounds <= 4'h0; // @[InvCipher.scala 32:23]
    end else if (2'h0 == STM) begin // @[InvCipher.scala 38:15]
      rounds <= 4'h0; // @[InvCipher.scala 43:14]
    end else if (2'h1 == STM) begin // @[InvCipher.scala 38:15]
      rounds <= _rounds_T_1; // @[InvCipher.scala 46:14]
    end else if (2'h2 == STM) begin // @[InvCipher.scala 38:15]
      rounds <= _rounds_T_1; // @[InvCipher.scala 50:14]
    end
    if (reset) begin // @[InvCipher.scala 36:20]
      STM <= 2'h0; // @[InvCipher.scala 36:20]
    end else if (2'h0 == STM) begin // @[InvCipher.scala 38:15]
      if (io_start) begin // @[InvCipher.scala 40:22]
        STM <= 2'h1; // @[InvCipher.scala 41:13]
      end
    end else if (2'h1 == STM) begin // @[InvCipher.scala 38:15]
      STM <= 2'h2; // @[InvCipher.scala 47:11]
    end else if (2'h2 == STM) begin // @[InvCipher.scala 38:15]
      STM <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  rounds = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  STM = _RAND_17[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AESDecrypt_1(
  input          clock,
  input          reset,
  input          io_input_valid,
  input  [255:0] io_input_text,
  output [255:0] io_output_text,
  output         io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  invcipher_A_clock; // @[InvCipher.scala 101:78]
  wire  invcipher_A_reset; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_ciphertext_15; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_roundKey_15; // @[InvCipher.scala 101:78]
  wire  invcipher_A_io_start; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_A_io_state_out_15; // @[InvCipher.scala 101:78]
  wire  invcipher_A_io_state_out_valid; // @[InvCipher.scala 101:78]
  wire  invcipher_B_clock; // @[InvCipher.scala 101:78]
  wire  invcipher_B_reset; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_ciphertext_15; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_roundKey_15; // @[InvCipher.scala 101:78]
  wire  invcipher_B_io_start; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_0; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_1; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_2; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_3; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_4; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_5; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_6; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_7; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_8; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_9; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_10; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_11; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_12; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_13; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_14; // @[InvCipher.scala 101:78]
  wire [7:0] invcipher_B_io_state_out_15; // @[InvCipher.scala 101:78]
  wire  invcipher_B_io_state_out_valid; // @[InvCipher.scala 101:78]
  reg [3:0] address; // @[AESDecrypt.scala 95:26]
  reg  tmp; // @[AESDecrypt.scala 97:22]
  wire [3:0] _address_T_1 = address - 4'h1; // @[AESDecrypt.scala 102:26]
  wire  _GEN_2 = io_input_valid & ~tmp | tmp; // @[AESDecrypt.scala 100:15 97:22 98:34]
  wire [7:0] _GEN_4 = 4'h1 == address ? 8'hd6 : 8'h0; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_5 = 4'h2 == address ? 8'hb6 : _GEN_4; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_6 = 4'h3 == address ? 8'hb6 : _GEN_5; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_7 = 4'h4 == address ? 8'h47 : _GEN_6; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_8 = 4'h5 == address ? 8'h3c : _GEN_7; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_9 = 4'h6 == address ? 8'h5e : _GEN_8; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_10 = 4'h7 == address ? 8'h14 : _GEN_9; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_11 = 4'h8 == address ? 8'h47 : _GEN_10; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_12 = 4'h9 == address ? 8'h54 : _GEN_11; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_15 = 4'h1 == address ? 8'haa : 8'h1; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_16 = 4'h2 == address ? 8'h92 : _GEN_15; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_17 = 4'h3 == address ? 8'hff : _GEN_16; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_18 = 4'h4 == address ? 8'hf7 : _GEN_17; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_19 = 4'h5 == address ? 8'haa : _GEN_18; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_20 = 4'h6 == address ? 8'h39 : _GEN_19; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_21 = 4'h7 == address ? 8'hf9 : _GEN_20; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_22 = 4'h8 == address ? 8'h43 : _GEN_21; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_23 = 4'h9 == address ? 8'h99 : _GEN_22; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_26 = 4'h1 == address ? 8'h74 : 8'h2; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_27 = 4'h2 == address ? 8'hcf : _GEN_26; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_28 = 4'h3 == address ? 8'h74 : _GEN_27; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_29 = 4'h4 == address ? 8'hf7 : _GEN_28; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_30 = 4'h5 == address ? 8'ha3 : _GEN_29; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_31 = 4'h6 == address ? 8'hf : _GEN_30; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_32 = 4'h7 == address ? 8'h70 : _GEN_31; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_33 = 4'h8 == address ? 8'h87 : _GEN_32; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_34 = 4'h9 == address ? 8'h32 : _GEN_33; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_37 = 4'h1 == address ? 8'hfd : 8'h3; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_38 = 4'h2 == address ? 8'hb : _GEN_37; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_39 = 4'h3 == address ? 8'h4e : _GEN_38; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_40 = 4'h4 == address ? 8'hbc : _GEN_39; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_41 = 4'h5 == address ? 8'he8 : _GEN_40; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_42 = 4'h6 == address ? 8'h7d : _GEN_41; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_43 = 4'h7 == address ? 8'h1a : _GEN_42; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_44 = 4'h8 == address ? 8'h35 : _GEN_43; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_45 = 4'h9 == address ? 8'hd1 : _GEN_44; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_48 = 4'h1 == address ? 8'hd2 : 8'h4; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_49 = 4'h2 == address ? 8'h64 : _GEN_48; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_50 = 4'h3 == address ? 8'hd2 : _GEN_49; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_51 = 4'h4 == address ? 8'h95 : _GEN_50; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_52 = 4'h5 == address ? 8'ha9 : _GEN_51; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_53 = 4'h6 == address ? 8'hf7 : _GEN_52; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_54 = 4'h7 == address ? 8'he3 : _GEN_53; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_55 = 4'h8 == address ? 8'ha4 : _GEN_54; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_56 = 4'h9 == address ? 8'hf0 : _GEN_55; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_59 = 4'h1 == address ? 8'haf : 8'h5; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_60 = 4'h2 == address ? 8'h3d : _GEN_59; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_61 = 4'h3 == address ? 8'hc2 : _GEN_60; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_62 = 4'h4 == address ? 8'h35 : _GEN_61; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_63 = 4'h5 == address ? 8'h9f : _GEN_62; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_64 = 4'h6 == address ? 8'ha6 : _GEN_63; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_65 = 4'h7 == address ? 8'h5f : _GEN_64; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_66 = 4'h8 == address ? 8'h1c : _GEN_65; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_67 = 4'h9 == address ? 8'h85 : _GEN_66; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_70 = 4'h1 == address ? 8'h72 : 8'h6; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_71 = 4'h2 == address ? 8'hbd : _GEN_70; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_72 = 4'h3 == address ? 8'hc9 : _GEN_71; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_73 = 4'h4 == address ? 8'h3e : _GEN_72; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_74 = 4'h5 == address ? 8'h9d : _GEN_73; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_75 = 4'h6 == address ? 8'h92 : _GEN_74; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_76 = 4'h7 == address ? 8'he2 : _GEN_75; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_77 = 4'h8 == address ? 8'h65 : _GEN_76; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_78 = 4'h9 == address ? 8'h57 : _GEN_77; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_81 = 4'h1 == address ? 8'hfa : 8'h7; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_82 = 4'h2 == address ? 8'hf1 : _GEN_81; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_83 = 4'h3 == address ? 8'hbf : _GEN_82; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_84 = 4'h4 == address ? 8'h3 : _GEN_83; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_85 = 4'h5 == address ? 8'heb : _GEN_84; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_86 = 4'h6 == address ? 8'h96 : _GEN_85; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_87 = 4'h7 == address ? 8'h8c : _GEN_86; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_88 = 4'h8 == address ? 8'hb9 : _GEN_87; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_89 = 4'h9 == address ? 8'h68 : _GEN_88; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_92 = 4'h1 == address ? 8'hda : 8'h8; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_93 = 4'h2 == address ? 8'hbe : _GEN_92; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_94 = 4'h3 == address ? 8'h6c : _GEN_93; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_95 = 4'h4 == address ? 8'hf9 : _GEN_94; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_96 = 4'h5 == address ? 8'h50 : _GEN_95; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_97 = 4'h6 == address ? 8'ha7 : _GEN_96; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_98 = 4'h7 == address ? 8'h44 : _GEN_97; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_99 = 4'h8 == address ? 8'he0 : _GEN_98; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_100 = 4'h9 == address ? 8'h10 : _GEN_99; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_103 = 4'h1 == address ? 8'ha6 : 8'h9; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_104 = 4'h2 == address ? 8'h9b : _GEN_103; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_105 = 4'h3 == address ? 8'h59 : _GEN_104; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_106 = 4'h4 == address ? 8'h6c : _GEN_105; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_107 = 4'h5 == address ? 8'hf3 : _GEN_106; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_108 = 4'h6 == address ? 8'h55 : _GEN_107; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_109 = 4'h7 == address ? 8'ha : _GEN_108; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_110 = 4'h8 == address ? 8'h16 : _GEN_109; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_111 = 4'h9 == address ? 8'h93 : _GEN_110; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_114 = 4'h1 == address ? 8'h78 : 8'ha; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_115 = 4'h2 == address ? 8'hc5 : _GEN_114; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_116 = 4'h3 == address ? 8'hc : _GEN_115; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_117 = 4'h4 == address ? 8'h32 : _GEN_116; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_118 = 4'h5 == address ? 8'haf : _GEN_117; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_119 = 4'h6 == address ? 8'h3d : _GEN_118; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_120 = 4'h7 == address ? 8'hdf : _GEN_119; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_121 = 4'h8 == address ? 8'hba : _GEN_120; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_122 = 4'h9 == address ? 8'hed : _GEN_121; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_125 = 4'h1 == address ? 8'hf1 : 8'hb; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_126 = 4'h2 == address ? 8'h0 : _GEN_125; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_127 = 4'h3 == address ? 8'hbf : _GEN_126; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_128 = 4'h4 == address ? 8'hbc : _GEN_127; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_129 = 4'h5 == address ? 8'h57 : _GEN_128; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_130 = 4'h6 == address ? 8'hc1 : _GEN_129; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_131 = 4'h7 == address ? 8'h4d : _GEN_130; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_132 = 4'h8 == address ? 8'hf4 : _GEN_131; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_133 = 4'h9 == address ? 8'h9c : _GEN_132; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_136 = 4'h1 == address ? 8'hd6 : 8'hc; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_137 = 4'h2 == address ? 8'h68 : _GEN_136; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_138 = 4'h3 == address ? 8'h4 : _GEN_137; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_139 = 4'h4 == address ? 8'hfd : _GEN_138; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_140 = 4'h5 == address ? 8'had : _GEN_139; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_141 = 4'h6 == address ? 8'ha : _GEN_140; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_142 = 4'h7 == address ? 8'h4e : _GEN_141; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_143 = 4'h8 == address ? 8'hae : _GEN_142; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_144 = 4'h9 == address ? 8'hbe : _GEN_143; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_147 = 4'h1 == address ? 8'hab : 8'hd; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_148 = 4'h2 == address ? 8'h30 : _GEN_147; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_149 = 4'h3 == address ? 8'h69 : _GEN_148; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_150 = 4'h4 == address ? 8'h5 : _GEN_149; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_151 = 4'h5 == address ? 8'hf6 : _GEN_150; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_152 = 4'h6 == address ? 8'ha3 : _GEN_151; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_153 = 4'h7 == address ? 8'ha9 : _GEN_152; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_154 = 4'h8 == address ? 8'hbf : _GEN_153; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_155 = 4'h9 == address ? 8'h2c : _GEN_154; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_158 = 4'h1 == address ? 8'h76 : 8'he; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_159 = 4'h2 == address ? 8'hb3 : _GEN_158; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_160 = 4'h3 == address ? 8'hbf : _GEN_159; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_161 = 4'h4 == address ? 8'h8d : _GEN_160; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_162 = 4'h5 == address ? 8'h22 : _GEN_161; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_163 = 4'h6 == address ? 8'h1f : _GEN_162; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_164 = 4'h7 == address ? 8'hc0 : _GEN_163; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_165 = 4'h8 == address ? 8'h7a : _GEN_164; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_166 = 4'h9 == address ? 8'h97 : _GEN_165; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_169 = 4'h1 == address ? 8'hfe : 8'hf; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_170 = 4'h2 == address ? 8'hfe : _GEN_169; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_171 = 4'h3 == address ? 8'h41 : _GEN_170; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_172 = 4'h4 == address ? 8'hfd : _GEN_171; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_173 = 4'h5 == address ? 8'haa : _GEN_172; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_174 = 4'h6 == address ? 8'h6b : _GEN_173; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_175 = 4'h7 == address ? 8'h26 : _GEN_174; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_176 = 4'h8 == address ? 8'hd2 : _GEN_175; // @[AESDecrypt.scala 106:{29,29}]
  wire [7:0] _GEN_177 = 4'h9 == address ? 8'h4e : _GEN_176; // @[AESDecrypt.scala 106:{29,29}]
  wire [63:0] io_output_text_lo = {invcipher_A_io_state_out_8,invcipher_A_io_state_out_9,invcipher_A_io_state_out_10,
    invcipher_A_io_state_out_11,invcipher_A_io_state_out_12,invcipher_A_io_state_out_13,invcipher_A_io_state_out_14,
    invcipher_A_io_state_out_15}; // @[Cat.scala 31:58]
  wire [127:0] _io_output_text_T = {invcipher_A_io_state_out_0,invcipher_A_io_state_out_1,invcipher_A_io_state_out_2,
    invcipher_A_io_state_out_3,invcipher_A_io_state_out_4,invcipher_A_io_state_out_5,invcipher_A_io_state_out_6,
    invcipher_A_io_state_out_7,io_output_text_lo}; // @[Cat.scala 31:58]
  wire [63:0] io_output_text_lo_1 = {invcipher_B_io_state_out_8,invcipher_B_io_state_out_9,invcipher_B_io_state_out_10,
    invcipher_B_io_state_out_11,invcipher_B_io_state_out_12,invcipher_B_io_state_out_13,invcipher_B_io_state_out_14,
    invcipher_B_io_state_out_15}; // @[Cat.scala 31:58]
  wire [127:0] _io_output_text_T_1 = {invcipher_B_io_state_out_0,invcipher_B_io_state_out_1,invcipher_B_io_state_out_2,
    invcipher_B_io_state_out_3,invcipher_B_io_state_out_4,invcipher_B_io_state_out_5,invcipher_B_io_state_out_6,
    invcipher_B_io_state_out_7,io_output_text_lo_1}; // @[Cat.scala 31:58]
  InvCipher_2 invcipher_A ( // @[InvCipher.scala 101:78]
    .clock(invcipher_A_clock),
    .reset(invcipher_A_reset),
    .io_ciphertext_0(invcipher_A_io_ciphertext_0),
    .io_ciphertext_1(invcipher_A_io_ciphertext_1),
    .io_ciphertext_2(invcipher_A_io_ciphertext_2),
    .io_ciphertext_3(invcipher_A_io_ciphertext_3),
    .io_ciphertext_4(invcipher_A_io_ciphertext_4),
    .io_ciphertext_5(invcipher_A_io_ciphertext_5),
    .io_ciphertext_6(invcipher_A_io_ciphertext_6),
    .io_ciphertext_7(invcipher_A_io_ciphertext_7),
    .io_ciphertext_8(invcipher_A_io_ciphertext_8),
    .io_ciphertext_9(invcipher_A_io_ciphertext_9),
    .io_ciphertext_10(invcipher_A_io_ciphertext_10),
    .io_ciphertext_11(invcipher_A_io_ciphertext_11),
    .io_ciphertext_12(invcipher_A_io_ciphertext_12),
    .io_ciphertext_13(invcipher_A_io_ciphertext_13),
    .io_ciphertext_14(invcipher_A_io_ciphertext_14),
    .io_ciphertext_15(invcipher_A_io_ciphertext_15),
    .io_roundKey_0(invcipher_A_io_roundKey_0),
    .io_roundKey_1(invcipher_A_io_roundKey_1),
    .io_roundKey_2(invcipher_A_io_roundKey_2),
    .io_roundKey_3(invcipher_A_io_roundKey_3),
    .io_roundKey_4(invcipher_A_io_roundKey_4),
    .io_roundKey_5(invcipher_A_io_roundKey_5),
    .io_roundKey_6(invcipher_A_io_roundKey_6),
    .io_roundKey_7(invcipher_A_io_roundKey_7),
    .io_roundKey_8(invcipher_A_io_roundKey_8),
    .io_roundKey_9(invcipher_A_io_roundKey_9),
    .io_roundKey_10(invcipher_A_io_roundKey_10),
    .io_roundKey_11(invcipher_A_io_roundKey_11),
    .io_roundKey_12(invcipher_A_io_roundKey_12),
    .io_roundKey_13(invcipher_A_io_roundKey_13),
    .io_roundKey_14(invcipher_A_io_roundKey_14),
    .io_roundKey_15(invcipher_A_io_roundKey_15),
    .io_start(invcipher_A_io_start),
    .io_state_out_0(invcipher_A_io_state_out_0),
    .io_state_out_1(invcipher_A_io_state_out_1),
    .io_state_out_2(invcipher_A_io_state_out_2),
    .io_state_out_3(invcipher_A_io_state_out_3),
    .io_state_out_4(invcipher_A_io_state_out_4),
    .io_state_out_5(invcipher_A_io_state_out_5),
    .io_state_out_6(invcipher_A_io_state_out_6),
    .io_state_out_7(invcipher_A_io_state_out_7),
    .io_state_out_8(invcipher_A_io_state_out_8),
    .io_state_out_9(invcipher_A_io_state_out_9),
    .io_state_out_10(invcipher_A_io_state_out_10),
    .io_state_out_11(invcipher_A_io_state_out_11),
    .io_state_out_12(invcipher_A_io_state_out_12),
    .io_state_out_13(invcipher_A_io_state_out_13),
    .io_state_out_14(invcipher_A_io_state_out_14),
    .io_state_out_15(invcipher_A_io_state_out_15),
    .io_state_out_valid(invcipher_A_io_state_out_valid)
  );
  InvCipher invcipher_B ( // @[InvCipher.scala 101:78]
    .clock(invcipher_B_clock),
    .reset(invcipher_B_reset),
    .io_ciphertext_0(invcipher_B_io_ciphertext_0),
    .io_ciphertext_1(invcipher_B_io_ciphertext_1),
    .io_ciphertext_2(invcipher_B_io_ciphertext_2),
    .io_ciphertext_3(invcipher_B_io_ciphertext_3),
    .io_ciphertext_4(invcipher_B_io_ciphertext_4),
    .io_ciphertext_5(invcipher_B_io_ciphertext_5),
    .io_ciphertext_6(invcipher_B_io_ciphertext_6),
    .io_ciphertext_7(invcipher_B_io_ciphertext_7),
    .io_ciphertext_8(invcipher_B_io_ciphertext_8),
    .io_ciphertext_9(invcipher_B_io_ciphertext_9),
    .io_ciphertext_10(invcipher_B_io_ciphertext_10),
    .io_ciphertext_11(invcipher_B_io_ciphertext_11),
    .io_ciphertext_12(invcipher_B_io_ciphertext_12),
    .io_ciphertext_13(invcipher_B_io_ciphertext_13),
    .io_ciphertext_14(invcipher_B_io_ciphertext_14),
    .io_ciphertext_15(invcipher_B_io_ciphertext_15),
    .io_roundKey_0(invcipher_B_io_roundKey_0),
    .io_roundKey_1(invcipher_B_io_roundKey_1),
    .io_roundKey_2(invcipher_B_io_roundKey_2),
    .io_roundKey_3(invcipher_B_io_roundKey_3),
    .io_roundKey_4(invcipher_B_io_roundKey_4),
    .io_roundKey_5(invcipher_B_io_roundKey_5),
    .io_roundKey_6(invcipher_B_io_roundKey_6),
    .io_roundKey_7(invcipher_B_io_roundKey_7),
    .io_roundKey_8(invcipher_B_io_roundKey_8),
    .io_roundKey_9(invcipher_B_io_roundKey_9),
    .io_roundKey_10(invcipher_B_io_roundKey_10),
    .io_roundKey_11(invcipher_B_io_roundKey_11),
    .io_roundKey_12(invcipher_B_io_roundKey_12),
    .io_roundKey_13(invcipher_B_io_roundKey_13),
    .io_roundKey_14(invcipher_B_io_roundKey_14),
    .io_roundKey_15(invcipher_B_io_roundKey_15),
    .io_start(invcipher_B_io_start),
    .io_state_out_0(invcipher_B_io_state_out_0),
    .io_state_out_1(invcipher_B_io_state_out_1),
    .io_state_out_2(invcipher_B_io_state_out_2),
    .io_state_out_3(invcipher_B_io_state_out_3),
    .io_state_out_4(invcipher_B_io_state_out_4),
    .io_state_out_5(invcipher_B_io_state_out_5),
    .io_state_out_6(invcipher_B_io_state_out_6),
    .io_state_out_7(invcipher_B_io_state_out_7),
    .io_state_out_8(invcipher_B_io_state_out_8),
    .io_state_out_9(invcipher_B_io_state_out_9),
    .io_state_out_10(invcipher_B_io_state_out_10),
    .io_state_out_11(invcipher_B_io_state_out_11),
    .io_state_out_12(invcipher_B_io_state_out_12),
    .io_state_out_13(invcipher_B_io_state_out_13),
    .io_state_out_14(invcipher_B_io_state_out_14),
    .io_state_out_15(invcipher_B_io_state_out_15),
    .io_state_out_valid(invcipher_B_io_state_out_valid)
  );
  assign io_output_text = {_io_output_text_T,_io_output_text_T_1}; // @[Cat.scala 31:58]
  assign io_output_valid = invcipher_A_io_state_out_valid & invcipher_B_io_state_out_valid; // @[AESDecrypt.scala 116:55]
  assign invcipher_A_clock = clock;
  assign invcipher_A_reset = reset;
  assign invcipher_A_io_ciphertext_0 = io_input_text[255:248]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_1 = io_input_text[247:240]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_2 = io_input_text[239:232]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_3 = io_input_text[231:224]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_4 = io_input_text[223:216]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_5 = io_input_text[215:208]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_6 = io_input_text[207:200]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_7 = io_input_text[199:192]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_8 = io_input_text[191:184]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_9 = io_input_text[183:176]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_10 = io_input_text[175:168]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_11 = io_input_text[167:160]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_12 = io_input_text[159:152]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_13 = io_input_text[151:144]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_14 = io_input_text[143:136]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_ciphertext_15 = io_input_text[135:128]; // @[AESDecrypt.scala 36:44]
  assign invcipher_A_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_A_io_start = io_input_valid; // @[AESDecrypt.scala 104:26]
  assign invcipher_B_clock = clock;
  assign invcipher_B_reset = reset;
  assign invcipher_B_io_ciphertext_0 = io_input_text[127:120]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_1 = io_input_text[119:112]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_2 = io_input_text[111:104]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_3 = io_input_text[103:96]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_4 = io_input_text[95:88]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_5 = io_input_text[87:80]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_6 = io_input_text[79:72]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_7 = io_input_text[71:64]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_8 = io_input_text[63:56]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_9 = io_input_text[55:48]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_10 = io_input_text[47:40]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_11 = io_input_text[39:32]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_12 = io_input_text[31:24]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_13 = io_input_text[23:16]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_14 = io_input_text[15:8]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_ciphertext_15 = io_input_text[7:0]; // @[AESDecrypt.scala 37:44]
  assign invcipher_B_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESDecrypt.scala 106:{29,29}]
  assign invcipher_B_io_start = io_input_valid; // @[AESDecrypt.scala 108:26]
  always @(posedge clock) begin
    if (reset) begin // @[AESDecrypt.scala 95:26]
      address <= 4'h0; // @[AESDecrypt.scala 95:26]
    end else if (io_input_valid & ~tmp) begin // @[AESDecrypt.scala 98:34]
      address <= 4'ha; // @[AESDecrypt.scala 99:15]
    end else if (address != 4'h0) begin // @[AESDecrypt.scala 101:32]
      address <= _address_T_1; // @[AESDecrypt.scala 102:15]
    end
    if (reset) begin // @[AESDecrypt.scala 97:22]
      tmp <= 1'h0; // @[AESDecrypt.scala 97:22]
    end else begin
      tmp <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  address = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  tmp = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SubBytes(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  wire [7:0] _GEN_1 = 8'h1 == io_state_in_0 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2 = 8'h2 == io_state_in_0 ? 8'h77 : _GEN_1; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3 = 8'h3 == io_state_in_0 ? 8'h7b : _GEN_2; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4 = 8'h4 == io_state_in_0 ? 8'hf2 : _GEN_3; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_5 = 8'h5 == io_state_in_0 ? 8'h6b : _GEN_4; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_6 = 8'h6 == io_state_in_0 ? 8'h6f : _GEN_5; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_7 = 8'h7 == io_state_in_0 ? 8'hc5 : _GEN_6; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_8 = 8'h8 == io_state_in_0 ? 8'h30 : _GEN_7; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_9 = 8'h9 == io_state_in_0 ? 8'h1 : _GEN_8; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_10 = 8'ha == io_state_in_0 ? 8'h67 : _GEN_9; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_11 = 8'hb == io_state_in_0 ? 8'h2b : _GEN_10; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_12 = 8'hc == io_state_in_0 ? 8'hfe : _GEN_11; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_13 = 8'hd == io_state_in_0 ? 8'hd7 : _GEN_12; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_14 = 8'he == io_state_in_0 ? 8'hab : _GEN_13; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_15 = 8'hf == io_state_in_0 ? 8'h76 : _GEN_14; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_16 = 8'h10 == io_state_in_0 ? 8'hca : _GEN_15; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_17 = 8'h11 == io_state_in_0 ? 8'h82 : _GEN_16; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_18 = 8'h12 == io_state_in_0 ? 8'hc9 : _GEN_17; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_19 = 8'h13 == io_state_in_0 ? 8'h7d : _GEN_18; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_20 = 8'h14 == io_state_in_0 ? 8'hfa : _GEN_19; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_21 = 8'h15 == io_state_in_0 ? 8'h59 : _GEN_20; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_22 = 8'h16 == io_state_in_0 ? 8'h47 : _GEN_21; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_23 = 8'h17 == io_state_in_0 ? 8'hf0 : _GEN_22; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_24 = 8'h18 == io_state_in_0 ? 8'had : _GEN_23; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_25 = 8'h19 == io_state_in_0 ? 8'hd4 : _GEN_24; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_26 = 8'h1a == io_state_in_0 ? 8'ha2 : _GEN_25; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_27 = 8'h1b == io_state_in_0 ? 8'haf : _GEN_26; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_28 = 8'h1c == io_state_in_0 ? 8'h9c : _GEN_27; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_29 = 8'h1d == io_state_in_0 ? 8'ha4 : _GEN_28; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_30 = 8'h1e == io_state_in_0 ? 8'h72 : _GEN_29; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_31 = 8'h1f == io_state_in_0 ? 8'hc0 : _GEN_30; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_32 = 8'h20 == io_state_in_0 ? 8'hb7 : _GEN_31; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_33 = 8'h21 == io_state_in_0 ? 8'hfd : _GEN_32; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_34 = 8'h22 == io_state_in_0 ? 8'h93 : _GEN_33; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_35 = 8'h23 == io_state_in_0 ? 8'h26 : _GEN_34; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_36 = 8'h24 == io_state_in_0 ? 8'h36 : _GEN_35; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_37 = 8'h25 == io_state_in_0 ? 8'h3f : _GEN_36; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_38 = 8'h26 == io_state_in_0 ? 8'hf7 : _GEN_37; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_39 = 8'h27 == io_state_in_0 ? 8'hcc : _GEN_38; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_40 = 8'h28 == io_state_in_0 ? 8'h34 : _GEN_39; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_41 = 8'h29 == io_state_in_0 ? 8'ha5 : _GEN_40; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_42 = 8'h2a == io_state_in_0 ? 8'he5 : _GEN_41; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_43 = 8'h2b == io_state_in_0 ? 8'hf1 : _GEN_42; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_44 = 8'h2c == io_state_in_0 ? 8'h71 : _GEN_43; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_45 = 8'h2d == io_state_in_0 ? 8'hd8 : _GEN_44; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_46 = 8'h2e == io_state_in_0 ? 8'h31 : _GEN_45; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_47 = 8'h2f == io_state_in_0 ? 8'h15 : _GEN_46; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_48 = 8'h30 == io_state_in_0 ? 8'h4 : _GEN_47; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_49 = 8'h31 == io_state_in_0 ? 8'hc7 : _GEN_48; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_50 = 8'h32 == io_state_in_0 ? 8'h23 : _GEN_49; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_51 = 8'h33 == io_state_in_0 ? 8'hc3 : _GEN_50; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_52 = 8'h34 == io_state_in_0 ? 8'h18 : _GEN_51; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_53 = 8'h35 == io_state_in_0 ? 8'h96 : _GEN_52; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_54 = 8'h36 == io_state_in_0 ? 8'h5 : _GEN_53; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_55 = 8'h37 == io_state_in_0 ? 8'h9a : _GEN_54; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_56 = 8'h38 == io_state_in_0 ? 8'h7 : _GEN_55; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_57 = 8'h39 == io_state_in_0 ? 8'h12 : _GEN_56; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_58 = 8'h3a == io_state_in_0 ? 8'h80 : _GEN_57; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_59 = 8'h3b == io_state_in_0 ? 8'he2 : _GEN_58; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_60 = 8'h3c == io_state_in_0 ? 8'heb : _GEN_59; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_61 = 8'h3d == io_state_in_0 ? 8'h27 : _GEN_60; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_62 = 8'h3e == io_state_in_0 ? 8'hb2 : _GEN_61; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_63 = 8'h3f == io_state_in_0 ? 8'h75 : _GEN_62; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_64 = 8'h40 == io_state_in_0 ? 8'h9 : _GEN_63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_65 = 8'h41 == io_state_in_0 ? 8'h83 : _GEN_64; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_66 = 8'h42 == io_state_in_0 ? 8'h2c : _GEN_65; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_67 = 8'h43 == io_state_in_0 ? 8'h1a : _GEN_66; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_68 = 8'h44 == io_state_in_0 ? 8'h1b : _GEN_67; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_69 = 8'h45 == io_state_in_0 ? 8'h6e : _GEN_68; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_70 = 8'h46 == io_state_in_0 ? 8'h5a : _GEN_69; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_71 = 8'h47 == io_state_in_0 ? 8'ha0 : _GEN_70; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_72 = 8'h48 == io_state_in_0 ? 8'h52 : _GEN_71; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_73 = 8'h49 == io_state_in_0 ? 8'h3b : _GEN_72; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_74 = 8'h4a == io_state_in_0 ? 8'hd6 : _GEN_73; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_75 = 8'h4b == io_state_in_0 ? 8'hb3 : _GEN_74; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_76 = 8'h4c == io_state_in_0 ? 8'h29 : _GEN_75; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_77 = 8'h4d == io_state_in_0 ? 8'he3 : _GEN_76; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_78 = 8'h4e == io_state_in_0 ? 8'h2f : _GEN_77; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_79 = 8'h4f == io_state_in_0 ? 8'h84 : _GEN_78; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_80 = 8'h50 == io_state_in_0 ? 8'h53 : _GEN_79; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_81 = 8'h51 == io_state_in_0 ? 8'hd1 : _GEN_80; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_82 = 8'h52 == io_state_in_0 ? 8'h0 : _GEN_81; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_83 = 8'h53 == io_state_in_0 ? 8'hed : _GEN_82; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_84 = 8'h54 == io_state_in_0 ? 8'h20 : _GEN_83; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_85 = 8'h55 == io_state_in_0 ? 8'hfc : _GEN_84; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_86 = 8'h56 == io_state_in_0 ? 8'hb1 : _GEN_85; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_87 = 8'h57 == io_state_in_0 ? 8'h5b : _GEN_86; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_88 = 8'h58 == io_state_in_0 ? 8'h6a : _GEN_87; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_89 = 8'h59 == io_state_in_0 ? 8'hcb : _GEN_88; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_90 = 8'h5a == io_state_in_0 ? 8'hbe : _GEN_89; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_91 = 8'h5b == io_state_in_0 ? 8'h39 : _GEN_90; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_92 = 8'h5c == io_state_in_0 ? 8'h4a : _GEN_91; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_93 = 8'h5d == io_state_in_0 ? 8'h4c : _GEN_92; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_94 = 8'h5e == io_state_in_0 ? 8'h58 : _GEN_93; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_95 = 8'h5f == io_state_in_0 ? 8'hcf : _GEN_94; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_96 = 8'h60 == io_state_in_0 ? 8'hd0 : _GEN_95; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_97 = 8'h61 == io_state_in_0 ? 8'hef : _GEN_96; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_98 = 8'h62 == io_state_in_0 ? 8'haa : _GEN_97; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_99 = 8'h63 == io_state_in_0 ? 8'hfb : _GEN_98; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_100 = 8'h64 == io_state_in_0 ? 8'h43 : _GEN_99; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_101 = 8'h65 == io_state_in_0 ? 8'h4d : _GEN_100; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_102 = 8'h66 == io_state_in_0 ? 8'h33 : _GEN_101; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_103 = 8'h67 == io_state_in_0 ? 8'h85 : _GEN_102; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_104 = 8'h68 == io_state_in_0 ? 8'h45 : _GEN_103; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_105 = 8'h69 == io_state_in_0 ? 8'hf9 : _GEN_104; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_106 = 8'h6a == io_state_in_0 ? 8'h2 : _GEN_105; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_107 = 8'h6b == io_state_in_0 ? 8'h7f : _GEN_106; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_108 = 8'h6c == io_state_in_0 ? 8'h50 : _GEN_107; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_109 = 8'h6d == io_state_in_0 ? 8'h3c : _GEN_108; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_110 = 8'h6e == io_state_in_0 ? 8'h9f : _GEN_109; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_111 = 8'h6f == io_state_in_0 ? 8'ha8 : _GEN_110; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_112 = 8'h70 == io_state_in_0 ? 8'h51 : _GEN_111; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_113 = 8'h71 == io_state_in_0 ? 8'ha3 : _GEN_112; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_114 = 8'h72 == io_state_in_0 ? 8'h40 : _GEN_113; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_115 = 8'h73 == io_state_in_0 ? 8'h8f : _GEN_114; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_116 = 8'h74 == io_state_in_0 ? 8'h92 : _GEN_115; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_117 = 8'h75 == io_state_in_0 ? 8'h9d : _GEN_116; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_118 = 8'h76 == io_state_in_0 ? 8'h38 : _GEN_117; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_119 = 8'h77 == io_state_in_0 ? 8'hf5 : _GEN_118; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_120 = 8'h78 == io_state_in_0 ? 8'hbc : _GEN_119; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_121 = 8'h79 == io_state_in_0 ? 8'hb6 : _GEN_120; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_122 = 8'h7a == io_state_in_0 ? 8'hda : _GEN_121; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_123 = 8'h7b == io_state_in_0 ? 8'h21 : _GEN_122; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_124 = 8'h7c == io_state_in_0 ? 8'h10 : _GEN_123; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_125 = 8'h7d == io_state_in_0 ? 8'hff : _GEN_124; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_126 = 8'h7e == io_state_in_0 ? 8'hf3 : _GEN_125; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_127 = 8'h7f == io_state_in_0 ? 8'hd2 : _GEN_126; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_128 = 8'h80 == io_state_in_0 ? 8'hcd : _GEN_127; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_129 = 8'h81 == io_state_in_0 ? 8'hc : _GEN_128; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_130 = 8'h82 == io_state_in_0 ? 8'h13 : _GEN_129; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_131 = 8'h83 == io_state_in_0 ? 8'hec : _GEN_130; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_132 = 8'h84 == io_state_in_0 ? 8'h5f : _GEN_131; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_133 = 8'h85 == io_state_in_0 ? 8'h97 : _GEN_132; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_134 = 8'h86 == io_state_in_0 ? 8'h44 : _GEN_133; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_135 = 8'h87 == io_state_in_0 ? 8'h17 : _GEN_134; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_136 = 8'h88 == io_state_in_0 ? 8'hc4 : _GEN_135; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_137 = 8'h89 == io_state_in_0 ? 8'ha7 : _GEN_136; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_138 = 8'h8a == io_state_in_0 ? 8'h7e : _GEN_137; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_139 = 8'h8b == io_state_in_0 ? 8'h3d : _GEN_138; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_140 = 8'h8c == io_state_in_0 ? 8'h64 : _GEN_139; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_141 = 8'h8d == io_state_in_0 ? 8'h5d : _GEN_140; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_142 = 8'h8e == io_state_in_0 ? 8'h19 : _GEN_141; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_143 = 8'h8f == io_state_in_0 ? 8'h73 : _GEN_142; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_144 = 8'h90 == io_state_in_0 ? 8'h60 : _GEN_143; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_145 = 8'h91 == io_state_in_0 ? 8'h81 : _GEN_144; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_146 = 8'h92 == io_state_in_0 ? 8'h4f : _GEN_145; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_147 = 8'h93 == io_state_in_0 ? 8'hdc : _GEN_146; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_148 = 8'h94 == io_state_in_0 ? 8'h22 : _GEN_147; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_149 = 8'h95 == io_state_in_0 ? 8'h2a : _GEN_148; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_150 = 8'h96 == io_state_in_0 ? 8'h90 : _GEN_149; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_151 = 8'h97 == io_state_in_0 ? 8'h88 : _GEN_150; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_152 = 8'h98 == io_state_in_0 ? 8'h46 : _GEN_151; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_153 = 8'h99 == io_state_in_0 ? 8'hee : _GEN_152; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_154 = 8'h9a == io_state_in_0 ? 8'hb8 : _GEN_153; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_155 = 8'h9b == io_state_in_0 ? 8'h14 : _GEN_154; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_156 = 8'h9c == io_state_in_0 ? 8'hde : _GEN_155; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_157 = 8'h9d == io_state_in_0 ? 8'h5e : _GEN_156; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_158 = 8'h9e == io_state_in_0 ? 8'hb : _GEN_157; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_159 = 8'h9f == io_state_in_0 ? 8'hdb : _GEN_158; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_160 = 8'ha0 == io_state_in_0 ? 8'he0 : _GEN_159; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_161 = 8'ha1 == io_state_in_0 ? 8'h32 : _GEN_160; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_162 = 8'ha2 == io_state_in_0 ? 8'h3a : _GEN_161; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_163 = 8'ha3 == io_state_in_0 ? 8'ha : _GEN_162; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_164 = 8'ha4 == io_state_in_0 ? 8'h49 : _GEN_163; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_165 = 8'ha5 == io_state_in_0 ? 8'h6 : _GEN_164; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_166 = 8'ha6 == io_state_in_0 ? 8'h24 : _GEN_165; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_167 = 8'ha7 == io_state_in_0 ? 8'h5c : _GEN_166; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_168 = 8'ha8 == io_state_in_0 ? 8'hc2 : _GEN_167; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_169 = 8'ha9 == io_state_in_0 ? 8'hd3 : _GEN_168; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_170 = 8'haa == io_state_in_0 ? 8'hac : _GEN_169; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_171 = 8'hab == io_state_in_0 ? 8'h62 : _GEN_170; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_172 = 8'hac == io_state_in_0 ? 8'h91 : _GEN_171; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_173 = 8'had == io_state_in_0 ? 8'h95 : _GEN_172; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_174 = 8'hae == io_state_in_0 ? 8'he4 : _GEN_173; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_175 = 8'haf == io_state_in_0 ? 8'h79 : _GEN_174; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_176 = 8'hb0 == io_state_in_0 ? 8'he7 : _GEN_175; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_177 = 8'hb1 == io_state_in_0 ? 8'hc8 : _GEN_176; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_178 = 8'hb2 == io_state_in_0 ? 8'h37 : _GEN_177; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_179 = 8'hb3 == io_state_in_0 ? 8'h6d : _GEN_178; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_180 = 8'hb4 == io_state_in_0 ? 8'h8d : _GEN_179; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_181 = 8'hb5 == io_state_in_0 ? 8'hd5 : _GEN_180; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_182 = 8'hb6 == io_state_in_0 ? 8'h4e : _GEN_181; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_183 = 8'hb7 == io_state_in_0 ? 8'ha9 : _GEN_182; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_184 = 8'hb8 == io_state_in_0 ? 8'h6c : _GEN_183; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_185 = 8'hb9 == io_state_in_0 ? 8'h56 : _GEN_184; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_186 = 8'hba == io_state_in_0 ? 8'hf4 : _GEN_185; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_187 = 8'hbb == io_state_in_0 ? 8'hea : _GEN_186; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_188 = 8'hbc == io_state_in_0 ? 8'h65 : _GEN_187; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_189 = 8'hbd == io_state_in_0 ? 8'h7a : _GEN_188; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_190 = 8'hbe == io_state_in_0 ? 8'hae : _GEN_189; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_191 = 8'hbf == io_state_in_0 ? 8'h8 : _GEN_190; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_192 = 8'hc0 == io_state_in_0 ? 8'hba : _GEN_191; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_193 = 8'hc1 == io_state_in_0 ? 8'h78 : _GEN_192; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_194 = 8'hc2 == io_state_in_0 ? 8'h25 : _GEN_193; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_195 = 8'hc3 == io_state_in_0 ? 8'h2e : _GEN_194; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_196 = 8'hc4 == io_state_in_0 ? 8'h1c : _GEN_195; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_197 = 8'hc5 == io_state_in_0 ? 8'ha6 : _GEN_196; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_198 = 8'hc6 == io_state_in_0 ? 8'hb4 : _GEN_197; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_199 = 8'hc7 == io_state_in_0 ? 8'hc6 : _GEN_198; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_200 = 8'hc8 == io_state_in_0 ? 8'he8 : _GEN_199; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_201 = 8'hc9 == io_state_in_0 ? 8'hdd : _GEN_200; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_202 = 8'hca == io_state_in_0 ? 8'h74 : _GEN_201; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_203 = 8'hcb == io_state_in_0 ? 8'h1f : _GEN_202; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_204 = 8'hcc == io_state_in_0 ? 8'h4b : _GEN_203; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_205 = 8'hcd == io_state_in_0 ? 8'hbd : _GEN_204; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_206 = 8'hce == io_state_in_0 ? 8'h8b : _GEN_205; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_207 = 8'hcf == io_state_in_0 ? 8'h8a : _GEN_206; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_208 = 8'hd0 == io_state_in_0 ? 8'h70 : _GEN_207; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_209 = 8'hd1 == io_state_in_0 ? 8'h3e : _GEN_208; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_210 = 8'hd2 == io_state_in_0 ? 8'hb5 : _GEN_209; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_211 = 8'hd3 == io_state_in_0 ? 8'h66 : _GEN_210; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_212 = 8'hd4 == io_state_in_0 ? 8'h48 : _GEN_211; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_213 = 8'hd5 == io_state_in_0 ? 8'h3 : _GEN_212; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_214 = 8'hd6 == io_state_in_0 ? 8'hf6 : _GEN_213; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_215 = 8'hd7 == io_state_in_0 ? 8'he : _GEN_214; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_216 = 8'hd8 == io_state_in_0 ? 8'h61 : _GEN_215; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_217 = 8'hd9 == io_state_in_0 ? 8'h35 : _GEN_216; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_218 = 8'hda == io_state_in_0 ? 8'h57 : _GEN_217; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_219 = 8'hdb == io_state_in_0 ? 8'hb9 : _GEN_218; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_220 = 8'hdc == io_state_in_0 ? 8'h86 : _GEN_219; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_221 = 8'hdd == io_state_in_0 ? 8'hc1 : _GEN_220; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_222 = 8'hde == io_state_in_0 ? 8'h1d : _GEN_221; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_223 = 8'hdf == io_state_in_0 ? 8'h9e : _GEN_222; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_224 = 8'he0 == io_state_in_0 ? 8'he1 : _GEN_223; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_225 = 8'he1 == io_state_in_0 ? 8'hf8 : _GEN_224; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_226 = 8'he2 == io_state_in_0 ? 8'h98 : _GEN_225; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_227 = 8'he3 == io_state_in_0 ? 8'h11 : _GEN_226; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_228 = 8'he4 == io_state_in_0 ? 8'h69 : _GEN_227; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_229 = 8'he5 == io_state_in_0 ? 8'hd9 : _GEN_228; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_230 = 8'he6 == io_state_in_0 ? 8'h8e : _GEN_229; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_231 = 8'he7 == io_state_in_0 ? 8'h94 : _GEN_230; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_232 = 8'he8 == io_state_in_0 ? 8'h9b : _GEN_231; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_233 = 8'he9 == io_state_in_0 ? 8'h1e : _GEN_232; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_234 = 8'hea == io_state_in_0 ? 8'h87 : _GEN_233; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_235 = 8'heb == io_state_in_0 ? 8'he9 : _GEN_234; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_236 = 8'hec == io_state_in_0 ? 8'hce : _GEN_235; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_237 = 8'hed == io_state_in_0 ? 8'h55 : _GEN_236; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_238 = 8'hee == io_state_in_0 ? 8'h28 : _GEN_237; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_239 = 8'hef == io_state_in_0 ? 8'hdf : _GEN_238; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_240 = 8'hf0 == io_state_in_0 ? 8'h8c : _GEN_239; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_241 = 8'hf1 == io_state_in_0 ? 8'ha1 : _GEN_240; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_242 = 8'hf2 == io_state_in_0 ? 8'h89 : _GEN_241; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_243 = 8'hf3 == io_state_in_0 ? 8'hd : _GEN_242; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_244 = 8'hf4 == io_state_in_0 ? 8'hbf : _GEN_243; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_245 = 8'hf5 == io_state_in_0 ? 8'he6 : _GEN_244; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_246 = 8'hf6 == io_state_in_0 ? 8'h42 : _GEN_245; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_247 = 8'hf7 == io_state_in_0 ? 8'h68 : _GEN_246; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_248 = 8'hf8 == io_state_in_0 ? 8'h41 : _GEN_247; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_249 = 8'hf9 == io_state_in_0 ? 8'h99 : _GEN_248; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_250 = 8'hfa == io_state_in_0 ? 8'h2d : _GEN_249; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_251 = 8'hfb == io_state_in_0 ? 8'hf : _GEN_250; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_252 = 8'hfc == io_state_in_0 ? 8'hb0 : _GEN_251; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_253 = 8'hfd == io_state_in_0 ? 8'h54 : _GEN_252; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_254 = 8'hfe == io_state_in_0 ? 8'hbb : _GEN_253; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_257 = 8'h1 == io_state_in_1 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_258 = 8'h2 == io_state_in_1 ? 8'h77 : _GEN_257; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_259 = 8'h3 == io_state_in_1 ? 8'h7b : _GEN_258; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_260 = 8'h4 == io_state_in_1 ? 8'hf2 : _GEN_259; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_261 = 8'h5 == io_state_in_1 ? 8'h6b : _GEN_260; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_262 = 8'h6 == io_state_in_1 ? 8'h6f : _GEN_261; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_263 = 8'h7 == io_state_in_1 ? 8'hc5 : _GEN_262; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_264 = 8'h8 == io_state_in_1 ? 8'h30 : _GEN_263; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_265 = 8'h9 == io_state_in_1 ? 8'h1 : _GEN_264; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_266 = 8'ha == io_state_in_1 ? 8'h67 : _GEN_265; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_267 = 8'hb == io_state_in_1 ? 8'h2b : _GEN_266; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_268 = 8'hc == io_state_in_1 ? 8'hfe : _GEN_267; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_269 = 8'hd == io_state_in_1 ? 8'hd7 : _GEN_268; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_270 = 8'he == io_state_in_1 ? 8'hab : _GEN_269; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_271 = 8'hf == io_state_in_1 ? 8'h76 : _GEN_270; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_272 = 8'h10 == io_state_in_1 ? 8'hca : _GEN_271; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_273 = 8'h11 == io_state_in_1 ? 8'h82 : _GEN_272; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_274 = 8'h12 == io_state_in_1 ? 8'hc9 : _GEN_273; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_275 = 8'h13 == io_state_in_1 ? 8'h7d : _GEN_274; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_276 = 8'h14 == io_state_in_1 ? 8'hfa : _GEN_275; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_277 = 8'h15 == io_state_in_1 ? 8'h59 : _GEN_276; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_278 = 8'h16 == io_state_in_1 ? 8'h47 : _GEN_277; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_279 = 8'h17 == io_state_in_1 ? 8'hf0 : _GEN_278; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_280 = 8'h18 == io_state_in_1 ? 8'had : _GEN_279; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_281 = 8'h19 == io_state_in_1 ? 8'hd4 : _GEN_280; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_282 = 8'h1a == io_state_in_1 ? 8'ha2 : _GEN_281; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_283 = 8'h1b == io_state_in_1 ? 8'haf : _GEN_282; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_284 = 8'h1c == io_state_in_1 ? 8'h9c : _GEN_283; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_285 = 8'h1d == io_state_in_1 ? 8'ha4 : _GEN_284; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_286 = 8'h1e == io_state_in_1 ? 8'h72 : _GEN_285; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_287 = 8'h1f == io_state_in_1 ? 8'hc0 : _GEN_286; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_288 = 8'h20 == io_state_in_1 ? 8'hb7 : _GEN_287; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_289 = 8'h21 == io_state_in_1 ? 8'hfd : _GEN_288; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_290 = 8'h22 == io_state_in_1 ? 8'h93 : _GEN_289; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_291 = 8'h23 == io_state_in_1 ? 8'h26 : _GEN_290; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_292 = 8'h24 == io_state_in_1 ? 8'h36 : _GEN_291; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_293 = 8'h25 == io_state_in_1 ? 8'h3f : _GEN_292; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_294 = 8'h26 == io_state_in_1 ? 8'hf7 : _GEN_293; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_295 = 8'h27 == io_state_in_1 ? 8'hcc : _GEN_294; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_296 = 8'h28 == io_state_in_1 ? 8'h34 : _GEN_295; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_297 = 8'h29 == io_state_in_1 ? 8'ha5 : _GEN_296; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_298 = 8'h2a == io_state_in_1 ? 8'he5 : _GEN_297; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_299 = 8'h2b == io_state_in_1 ? 8'hf1 : _GEN_298; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_300 = 8'h2c == io_state_in_1 ? 8'h71 : _GEN_299; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_301 = 8'h2d == io_state_in_1 ? 8'hd8 : _GEN_300; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_302 = 8'h2e == io_state_in_1 ? 8'h31 : _GEN_301; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_303 = 8'h2f == io_state_in_1 ? 8'h15 : _GEN_302; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_304 = 8'h30 == io_state_in_1 ? 8'h4 : _GEN_303; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_305 = 8'h31 == io_state_in_1 ? 8'hc7 : _GEN_304; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_306 = 8'h32 == io_state_in_1 ? 8'h23 : _GEN_305; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_307 = 8'h33 == io_state_in_1 ? 8'hc3 : _GEN_306; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_308 = 8'h34 == io_state_in_1 ? 8'h18 : _GEN_307; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_309 = 8'h35 == io_state_in_1 ? 8'h96 : _GEN_308; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_310 = 8'h36 == io_state_in_1 ? 8'h5 : _GEN_309; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_311 = 8'h37 == io_state_in_1 ? 8'h9a : _GEN_310; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_312 = 8'h38 == io_state_in_1 ? 8'h7 : _GEN_311; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_313 = 8'h39 == io_state_in_1 ? 8'h12 : _GEN_312; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_314 = 8'h3a == io_state_in_1 ? 8'h80 : _GEN_313; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_315 = 8'h3b == io_state_in_1 ? 8'he2 : _GEN_314; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_316 = 8'h3c == io_state_in_1 ? 8'heb : _GEN_315; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_317 = 8'h3d == io_state_in_1 ? 8'h27 : _GEN_316; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_318 = 8'h3e == io_state_in_1 ? 8'hb2 : _GEN_317; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_319 = 8'h3f == io_state_in_1 ? 8'h75 : _GEN_318; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_320 = 8'h40 == io_state_in_1 ? 8'h9 : _GEN_319; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_321 = 8'h41 == io_state_in_1 ? 8'h83 : _GEN_320; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_322 = 8'h42 == io_state_in_1 ? 8'h2c : _GEN_321; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_323 = 8'h43 == io_state_in_1 ? 8'h1a : _GEN_322; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_324 = 8'h44 == io_state_in_1 ? 8'h1b : _GEN_323; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_325 = 8'h45 == io_state_in_1 ? 8'h6e : _GEN_324; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_326 = 8'h46 == io_state_in_1 ? 8'h5a : _GEN_325; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_327 = 8'h47 == io_state_in_1 ? 8'ha0 : _GEN_326; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_328 = 8'h48 == io_state_in_1 ? 8'h52 : _GEN_327; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_329 = 8'h49 == io_state_in_1 ? 8'h3b : _GEN_328; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_330 = 8'h4a == io_state_in_1 ? 8'hd6 : _GEN_329; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_331 = 8'h4b == io_state_in_1 ? 8'hb3 : _GEN_330; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_332 = 8'h4c == io_state_in_1 ? 8'h29 : _GEN_331; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_333 = 8'h4d == io_state_in_1 ? 8'he3 : _GEN_332; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_334 = 8'h4e == io_state_in_1 ? 8'h2f : _GEN_333; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_335 = 8'h4f == io_state_in_1 ? 8'h84 : _GEN_334; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_336 = 8'h50 == io_state_in_1 ? 8'h53 : _GEN_335; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_337 = 8'h51 == io_state_in_1 ? 8'hd1 : _GEN_336; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_338 = 8'h52 == io_state_in_1 ? 8'h0 : _GEN_337; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_339 = 8'h53 == io_state_in_1 ? 8'hed : _GEN_338; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_340 = 8'h54 == io_state_in_1 ? 8'h20 : _GEN_339; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_341 = 8'h55 == io_state_in_1 ? 8'hfc : _GEN_340; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_342 = 8'h56 == io_state_in_1 ? 8'hb1 : _GEN_341; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_343 = 8'h57 == io_state_in_1 ? 8'h5b : _GEN_342; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_344 = 8'h58 == io_state_in_1 ? 8'h6a : _GEN_343; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_345 = 8'h59 == io_state_in_1 ? 8'hcb : _GEN_344; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_346 = 8'h5a == io_state_in_1 ? 8'hbe : _GEN_345; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_347 = 8'h5b == io_state_in_1 ? 8'h39 : _GEN_346; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_348 = 8'h5c == io_state_in_1 ? 8'h4a : _GEN_347; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_349 = 8'h5d == io_state_in_1 ? 8'h4c : _GEN_348; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_350 = 8'h5e == io_state_in_1 ? 8'h58 : _GEN_349; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_351 = 8'h5f == io_state_in_1 ? 8'hcf : _GEN_350; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_352 = 8'h60 == io_state_in_1 ? 8'hd0 : _GEN_351; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_353 = 8'h61 == io_state_in_1 ? 8'hef : _GEN_352; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_354 = 8'h62 == io_state_in_1 ? 8'haa : _GEN_353; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_355 = 8'h63 == io_state_in_1 ? 8'hfb : _GEN_354; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_356 = 8'h64 == io_state_in_1 ? 8'h43 : _GEN_355; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_357 = 8'h65 == io_state_in_1 ? 8'h4d : _GEN_356; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_358 = 8'h66 == io_state_in_1 ? 8'h33 : _GEN_357; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_359 = 8'h67 == io_state_in_1 ? 8'h85 : _GEN_358; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_360 = 8'h68 == io_state_in_1 ? 8'h45 : _GEN_359; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_361 = 8'h69 == io_state_in_1 ? 8'hf9 : _GEN_360; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_362 = 8'h6a == io_state_in_1 ? 8'h2 : _GEN_361; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_363 = 8'h6b == io_state_in_1 ? 8'h7f : _GEN_362; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_364 = 8'h6c == io_state_in_1 ? 8'h50 : _GEN_363; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_365 = 8'h6d == io_state_in_1 ? 8'h3c : _GEN_364; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_366 = 8'h6e == io_state_in_1 ? 8'h9f : _GEN_365; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_367 = 8'h6f == io_state_in_1 ? 8'ha8 : _GEN_366; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_368 = 8'h70 == io_state_in_1 ? 8'h51 : _GEN_367; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_369 = 8'h71 == io_state_in_1 ? 8'ha3 : _GEN_368; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_370 = 8'h72 == io_state_in_1 ? 8'h40 : _GEN_369; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_371 = 8'h73 == io_state_in_1 ? 8'h8f : _GEN_370; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_372 = 8'h74 == io_state_in_1 ? 8'h92 : _GEN_371; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_373 = 8'h75 == io_state_in_1 ? 8'h9d : _GEN_372; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_374 = 8'h76 == io_state_in_1 ? 8'h38 : _GEN_373; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_375 = 8'h77 == io_state_in_1 ? 8'hf5 : _GEN_374; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_376 = 8'h78 == io_state_in_1 ? 8'hbc : _GEN_375; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_377 = 8'h79 == io_state_in_1 ? 8'hb6 : _GEN_376; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_378 = 8'h7a == io_state_in_1 ? 8'hda : _GEN_377; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_379 = 8'h7b == io_state_in_1 ? 8'h21 : _GEN_378; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_380 = 8'h7c == io_state_in_1 ? 8'h10 : _GEN_379; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_381 = 8'h7d == io_state_in_1 ? 8'hff : _GEN_380; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_382 = 8'h7e == io_state_in_1 ? 8'hf3 : _GEN_381; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_383 = 8'h7f == io_state_in_1 ? 8'hd2 : _GEN_382; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_384 = 8'h80 == io_state_in_1 ? 8'hcd : _GEN_383; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_385 = 8'h81 == io_state_in_1 ? 8'hc : _GEN_384; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_386 = 8'h82 == io_state_in_1 ? 8'h13 : _GEN_385; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_387 = 8'h83 == io_state_in_1 ? 8'hec : _GEN_386; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_388 = 8'h84 == io_state_in_1 ? 8'h5f : _GEN_387; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_389 = 8'h85 == io_state_in_1 ? 8'h97 : _GEN_388; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_390 = 8'h86 == io_state_in_1 ? 8'h44 : _GEN_389; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_391 = 8'h87 == io_state_in_1 ? 8'h17 : _GEN_390; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_392 = 8'h88 == io_state_in_1 ? 8'hc4 : _GEN_391; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_393 = 8'h89 == io_state_in_1 ? 8'ha7 : _GEN_392; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_394 = 8'h8a == io_state_in_1 ? 8'h7e : _GEN_393; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_395 = 8'h8b == io_state_in_1 ? 8'h3d : _GEN_394; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_396 = 8'h8c == io_state_in_1 ? 8'h64 : _GEN_395; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_397 = 8'h8d == io_state_in_1 ? 8'h5d : _GEN_396; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_398 = 8'h8e == io_state_in_1 ? 8'h19 : _GEN_397; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_399 = 8'h8f == io_state_in_1 ? 8'h73 : _GEN_398; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_400 = 8'h90 == io_state_in_1 ? 8'h60 : _GEN_399; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_401 = 8'h91 == io_state_in_1 ? 8'h81 : _GEN_400; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_402 = 8'h92 == io_state_in_1 ? 8'h4f : _GEN_401; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_403 = 8'h93 == io_state_in_1 ? 8'hdc : _GEN_402; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_404 = 8'h94 == io_state_in_1 ? 8'h22 : _GEN_403; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_405 = 8'h95 == io_state_in_1 ? 8'h2a : _GEN_404; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_406 = 8'h96 == io_state_in_1 ? 8'h90 : _GEN_405; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_407 = 8'h97 == io_state_in_1 ? 8'h88 : _GEN_406; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_408 = 8'h98 == io_state_in_1 ? 8'h46 : _GEN_407; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_409 = 8'h99 == io_state_in_1 ? 8'hee : _GEN_408; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_410 = 8'h9a == io_state_in_1 ? 8'hb8 : _GEN_409; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_411 = 8'h9b == io_state_in_1 ? 8'h14 : _GEN_410; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_412 = 8'h9c == io_state_in_1 ? 8'hde : _GEN_411; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_413 = 8'h9d == io_state_in_1 ? 8'h5e : _GEN_412; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_414 = 8'h9e == io_state_in_1 ? 8'hb : _GEN_413; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_415 = 8'h9f == io_state_in_1 ? 8'hdb : _GEN_414; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_416 = 8'ha0 == io_state_in_1 ? 8'he0 : _GEN_415; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_417 = 8'ha1 == io_state_in_1 ? 8'h32 : _GEN_416; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_418 = 8'ha2 == io_state_in_1 ? 8'h3a : _GEN_417; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_419 = 8'ha3 == io_state_in_1 ? 8'ha : _GEN_418; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_420 = 8'ha4 == io_state_in_1 ? 8'h49 : _GEN_419; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_421 = 8'ha5 == io_state_in_1 ? 8'h6 : _GEN_420; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_422 = 8'ha6 == io_state_in_1 ? 8'h24 : _GEN_421; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_423 = 8'ha7 == io_state_in_1 ? 8'h5c : _GEN_422; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_424 = 8'ha8 == io_state_in_1 ? 8'hc2 : _GEN_423; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_425 = 8'ha9 == io_state_in_1 ? 8'hd3 : _GEN_424; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_426 = 8'haa == io_state_in_1 ? 8'hac : _GEN_425; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_427 = 8'hab == io_state_in_1 ? 8'h62 : _GEN_426; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_428 = 8'hac == io_state_in_1 ? 8'h91 : _GEN_427; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_429 = 8'had == io_state_in_1 ? 8'h95 : _GEN_428; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_430 = 8'hae == io_state_in_1 ? 8'he4 : _GEN_429; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_431 = 8'haf == io_state_in_1 ? 8'h79 : _GEN_430; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_432 = 8'hb0 == io_state_in_1 ? 8'he7 : _GEN_431; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_433 = 8'hb1 == io_state_in_1 ? 8'hc8 : _GEN_432; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_434 = 8'hb2 == io_state_in_1 ? 8'h37 : _GEN_433; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_435 = 8'hb3 == io_state_in_1 ? 8'h6d : _GEN_434; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_436 = 8'hb4 == io_state_in_1 ? 8'h8d : _GEN_435; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_437 = 8'hb5 == io_state_in_1 ? 8'hd5 : _GEN_436; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_438 = 8'hb6 == io_state_in_1 ? 8'h4e : _GEN_437; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_439 = 8'hb7 == io_state_in_1 ? 8'ha9 : _GEN_438; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_440 = 8'hb8 == io_state_in_1 ? 8'h6c : _GEN_439; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_441 = 8'hb9 == io_state_in_1 ? 8'h56 : _GEN_440; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_442 = 8'hba == io_state_in_1 ? 8'hf4 : _GEN_441; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_443 = 8'hbb == io_state_in_1 ? 8'hea : _GEN_442; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_444 = 8'hbc == io_state_in_1 ? 8'h65 : _GEN_443; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_445 = 8'hbd == io_state_in_1 ? 8'h7a : _GEN_444; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_446 = 8'hbe == io_state_in_1 ? 8'hae : _GEN_445; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_447 = 8'hbf == io_state_in_1 ? 8'h8 : _GEN_446; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_448 = 8'hc0 == io_state_in_1 ? 8'hba : _GEN_447; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_449 = 8'hc1 == io_state_in_1 ? 8'h78 : _GEN_448; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_450 = 8'hc2 == io_state_in_1 ? 8'h25 : _GEN_449; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_451 = 8'hc3 == io_state_in_1 ? 8'h2e : _GEN_450; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_452 = 8'hc4 == io_state_in_1 ? 8'h1c : _GEN_451; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_453 = 8'hc5 == io_state_in_1 ? 8'ha6 : _GEN_452; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_454 = 8'hc6 == io_state_in_1 ? 8'hb4 : _GEN_453; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_455 = 8'hc7 == io_state_in_1 ? 8'hc6 : _GEN_454; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_456 = 8'hc8 == io_state_in_1 ? 8'he8 : _GEN_455; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_457 = 8'hc9 == io_state_in_1 ? 8'hdd : _GEN_456; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_458 = 8'hca == io_state_in_1 ? 8'h74 : _GEN_457; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_459 = 8'hcb == io_state_in_1 ? 8'h1f : _GEN_458; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_460 = 8'hcc == io_state_in_1 ? 8'h4b : _GEN_459; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_461 = 8'hcd == io_state_in_1 ? 8'hbd : _GEN_460; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_462 = 8'hce == io_state_in_1 ? 8'h8b : _GEN_461; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_463 = 8'hcf == io_state_in_1 ? 8'h8a : _GEN_462; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_464 = 8'hd0 == io_state_in_1 ? 8'h70 : _GEN_463; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_465 = 8'hd1 == io_state_in_1 ? 8'h3e : _GEN_464; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_466 = 8'hd2 == io_state_in_1 ? 8'hb5 : _GEN_465; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_467 = 8'hd3 == io_state_in_1 ? 8'h66 : _GEN_466; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_468 = 8'hd4 == io_state_in_1 ? 8'h48 : _GEN_467; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_469 = 8'hd5 == io_state_in_1 ? 8'h3 : _GEN_468; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_470 = 8'hd6 == io_state_in_1 ? 8'hf6 : _GEN_469; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_471 = 8'hd7 == io_state_in_1 ? 8'he : _GEN_470; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_472 = 8'hd8 == io_state_in_1 ? 8'h61 : _GEN_471; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_473 = 8'hd9 == io_state_in_1 ? 8'h35 : _GEN_472; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_474 = 8'hda == io_state_in_1 ? 8'h57 : _GEN_473; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_475 = 8'hdb == io_state_in_1 ? 8'hb9 : _GEN_474; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_476 = 8'hdc == io_state_in_1 ? 8'h86 : _GEN_475; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_477 = 8'hdd == io_state_in_1 ? 8'hc1 : _GEN_476; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_478 = 8'hde == io_state_in_1 ? 8'h1d : _GEN_477; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_479 = 8'hdf == io_state_in_1 ? 8'h9e : _GEN_478; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_480 = 8'he0 == io_state_in_1 ? 8'he1 : _GEN_479; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_481 = 8'he1 == io_state_in_1 ? 8'hf8 : _GEN_480; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_482 = 8'he2 == io_state_in_1 ? 8'h98 : _GEN_481; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_483 = 8'he3 == io_state_in_1 ? 8'h11 : _GEN_482; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_484 = 8'he4 == io_state_in_1 ? 8'h69 : _GEN_483; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_485 = 8'he5 == io_state_in_1 ? 8'hd9 : _GEN_484; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_486 = 8'he6 == io_state_in_1 ? 8'h8e : _GEN_485; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_487 = 8'he7 == io_state_in_1 ? 8'h94 : _GEN_486; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_488 = 8'he8 == io_state_in_1 ? 8'h9b : _GEN_487; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_489 = 8'he9 == io_state_in_1 ? 8'h1e : _GEN_488; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_490 = 8'hea == io_state_in_1 ? 8'h87 : _GEN_489; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_491 = 8'heb == io_state_in_1 ? 8'he9 : _GEN_490; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_492 = 8'hec == io_state_in_1 ? 8'hce : _GEN_491; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_493 = 8'hed == io_state_in_1 ? 8'h55 : _GEN_492; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_494 = 8'hee == io_state_in_1 ? 8'h28 : _GEN_493; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_495 = 8'hef == io_state_in_1 ? 8'hdf : _GEN_494; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_496 = 8'hf0 == io_state_in_1 ? 8'h8c : _GEN_495; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_497 = 8'hf1 == io_state_in_1 ? 8'ha1 : _GEN_496; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_498 = 8'hf2 == io_state_in_1 ? 8'h89 : _GEN_497; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_499 = 8'hf3 == io_state_in_1 ? 8'hd : _GEN_498; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_500 = 8'hf4 == io_state_in_1 ? 8'hbf : _GEN_499; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_501 = 8'hf5 == io_state_in_1 ? 8'he6 : _GEN_500; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_502 = 8'hf6 == io_state_in_1 ? 8'h42 : _GEN_501; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_503 = 8'hf7 == io_state_in_1 ? 8'h68 : _GEN_502; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_504 = 8'hf8 == io_state_in_1 ? 8'h41 : _GEN_503; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_505 = 8'hf9 == io_state_in_1 ? 8'h99 : _GEN_504; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_506 = 8'hfa == io_state_in_1 ? 8'h2d : _GEN_505; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_507 = 8'hfb == io_state_in_1 ? 8'hf : _GEN_506; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_508 = 8'hfc == io_state_in_1 ? 8'hb0 : _GEN_507; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_509 = 8'hfd == io_state_in_1 ? 8'h54 : _GEN_508; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_510 = 8'hfe == io_state_in_1 ? 8'hbb : _GEN_509; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_513 = 8'h1 == io_state_in_2 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_514 = 8'h2 == io_state_in_2 ? 8'h77 : _GEN_513; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_515 = 8'h3 == io_state_in_2 ? 8'h7b : _GEN_514; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_516 = 8'h4 == io_state_in_2 ? 8'hf2 : _GEN_515; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_517 = 8'h5 == io_state_in_2 ? 8'h6b : _GEN_516; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_518 = 8'h6 == io_state_in_2 ? 8'h6f : _GEN_517; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_519 = 8'h7 == io_state_in_2 ? 8'hc5 : _GEN_518; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_520 = 8'h8 == io_state_in_2 ? 8'h30 : _GEN_519; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_521 = 8'h9 == io_state_in_2 ? 8'h1 : _GEN_520; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_522 = 8'ha == io_state_in_2 ? 8'h67 : _GEN_521; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_523 = 8'hb == io_state_in_2 ? 8'h2b : _GEN_522; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_524 = 8'hc == io_state_in_2 ? 8'hfe : _GEN_523; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_525 = 8'hd == io_state_in_2 ? 8'hd7 : _GEN_524; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_526 = 8'he == io_state_in_2 ? 8'hab : _GEN_525; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_527 = 8'hf == io_state_in_2 ? 8'h76 : _GEN_526; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_528 = 8'h10 == io_state_in_2 ? 8'hca : _GEN_527; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_529 = 8'h11 == io_state_in_2 ? 8'h82 : _GEN_528; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_530 = 8'h12 == io_state_in_2 ? 8'hc9 : _GEN_529; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_531 = 8'h13 == io_state_in_2 ? 8'h7d : _GEN_530; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_532 = 8'h14 == io_state_in_2 ? 8'hfa : _GEN_531; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_533 = 8'h15 == io_state_in_2 ? 8'h59 : _GEN_532; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_534 = 8'h16 == io_state_in_2 ? 8'h47 : _GEN_533; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_535 = 8'h17 == io_state_in_2 ? 8'hf0 : _GEN_534; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_536 = 8'h18 == io_state_in_2 ? 8'had : _GEN_535; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_537 = 8'h19 == io_state_in_2 ? 8'hd4 : _GEN_536; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_538 = 8'h1a == io_state_in_2 ? 8'ha2 : _GEN_537; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_539 = 8'h1b == io_state_in_2 ? 8'haf : _GEN_538; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_540 = 8'h1c == io_state_in_2 ? 8'h9c : _GEN_539; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_541 = 8'h1d == io_state_in_2 ? 8'ha4 : _GEN_540; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_542 = 8'h1e == io_state_in_2 ? 8'h72 : _GEN_541; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_543 = 8'h1f == io_state_in_2 ? 8'hc0 : _GEN_542; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_544 = 8'h20 == io_state_in_2 ? 8'hb7 : _GEN_543; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_545 = 8'h21 == io_state_in_2 ? 8'hfd : _GEN_544; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_546 = 8'h22 == io_state_in_2 ? 8'h93 : _GEN_545; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_547 = 8'h23 == io_state_in_2 ? 8'h26 : _GEN_546; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_548 = 8'h24 == io_state_in_2 ? 8'h36 : _GEN_547; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_549 = 8'h25 == io_state_in_2 ? 8'h3f : _GEN_548; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_550 = 8'h26 == io_state_in_2 ? 8'hf7 : _GEN_549; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_551 = 8'h27 == io_state_in_2 ? 8'hcc : _GEN_550; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_552 = 8'h28 == io_state_in_2 ? 8'h34 : _GEN_551; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_553 = 8'h29 == io_state_in_2 ? 8'ha5 : _GEN_552; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_554 = 8'h2a == io_state_in_2 ? 8'he5 : _GEN_553; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_555 = 8'h2b == io_state_in_2 ? 8'hf1 : _GEN_554; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_556 = 8'h2c == io_state_in_2 ? 8'h71 : _GEN_555; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_557 = 8'h2d == io_state_in_2 ? 8'hd8 : _GEN_556; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_558 = 8'h2e == io_state_in_2 ? 8'h31 : _GEN_557; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_559 = 8'h2f == io_state_in_2 ? 8'h15 : _GEN_558; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_560 = 8'h30 == io_state_in_2 ? 8'h4 : _GEN_559; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_561 = 8'h31 == io_state_in_2 ? 8'hc7 : _GEN_560; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_562 = 8'h32 == io_state_in_2 ? 8'h23 : _GEN_561; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_563 = 8'h33 == io_state_in_2 ? 8'hc3 : _GEN_562; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_564 = 8'h34 == io_state_in_2 ? 8'h18 : _GEN_563; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_565 = 8'h35 == io_state_in_2 ? 8'h96 : _GEN_564; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_566 = 8'h36 == io_state_in_2 ? 8'h5 : _GEN_565; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_567 = 8'h37 == io_state_in_2 ? 8'h9a : _GEN_566; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_568 = 8'h38 == io_state_in_2 ? 8'h7 : _GEN_567; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_569 = 8'h39 == io_state_in_2 ? 8'h12 : _GEN_568; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_570 = 8'h3a == io_state_in_2 ? 8'h80 : _GEN_569; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_571 = 8'h3b == io_state_in_2 ? 8'he2 : _GEN_570; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_572 = 8'h3c == io_state_in_2 ? 8'heb : _GEN_571; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_573 = 8'h3d == io_state_in_2 ? 8'h27 : _GEN_572; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_574 = 8'h3e == io_state_in_2 ? 8'hb2 : _GEN_573; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_575 = 8'h3f == io_state_in_2 ? 8'h75 : _GEN_574; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_576 = 8'h40 == io_state_in_2 ? 8'h9 : _GEN_575; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_577 = 8'h41 == io_state_in_2 ? 8'h83 : _GEN_576; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_578 = 8'h42 == io_state_in_2 ? 8'h2c : _GEN_577; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_579 = 8'h43 == io_state_in_2 ? 8'h1a : _GEN_578; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_580 = 8'h44 == io_state_in_2 ? 8'h1b : _GEN_579; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_581 = 8'h45 == io_state_in_2 ? 8'h6e : _GEN_580; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_582 = 8'h46 == io_state_in_2 ? 8'h5a : _GEN_581; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_583 = 8'h47 == io_state_in_2 ? 8'ha0 : _GEN_582; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_584 = 8'h48 == io_state_in_2 ? 8'h52 : _GEN_583; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_585 = 8'h49 == io_state_in_2 ? 8'h3b : _GEN_584; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_586 = 8'h4a == io_state_in_2 ? 8'hd6 : _GEN_585; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_587 = 8'h4b == io_state_in_2 ? 8'hb3 : _GEN_586; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_588 = 8'h4c == io_state_in_2 ? 8'h29 : _GEN_587; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_589 = 8'h4d == io_state_in_2 ? 8'he3 : _GEN_588; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_590 = 8'h4e == io_state_in_2 ? 8'h2f : _GEN_589; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_591 = 8'h4f == io_state_in_2 ? 8'h84 : _GEN_590; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_592 = 8'h50 == io_state_in_2 ? 8'h53 : _GEN_591; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_593 = 8'h51 == io_state_in_2 ? 8'hd1 : _GEN_592; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_594 = 8'h52 == io_state_in_2 ? 8'h0 : _GEN_593; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_595 = 8'h53 == io_state_in_2 ? 8'hed : _GEN_594; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_596 = 8'h54 == io_state_in_2 ? 8'h20 : _GEN_595; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_597 = 8'h55 == io_state_in_2 ? 8'hfc : _GEN_596; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_598 = 8'h56 == io_state_in_2 ? 8'hb1 : _GEN_597; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_599 = 8'h57 == io_state_in_2 ? 8'h5b : _GEN_598; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_600 = 8'h58 == io_state_in_2 ? 8'h6a : _GEN_599; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_601 = 8'h59 == io_state_in_2 ? 8'hcb : _GEN_600; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_602 = 8'h5a == io_state_in_2 ? 8'hbe : _GEN_601; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_603 = 8'h5b == io_state_in_2 ? 8'h39 : _GEN_602; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_604 = 8'h5c == io_state_in_2 ? 8'h4a : _GEN_603; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_605 = 8'h5d == io_state_in_2 ? 8'h4c : _GEN_604; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_606 = 8'h5e == io_state_in_2 ? 8'h58 : _GEN_605; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_607 = 8'h5f == io_state_in_2 ? 8'hcf : _GEN_606; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_608 = 8'h60 == io_state_in_2 ? 8'hd0 : _GEN_607; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_609 = 8'h61 == io_state_in_2 ? 8'hef : _GEN_608; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_610 = 8'h62 == io_state_in_2 ? 8'haa : _GEN_609; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_611 = 8'h63 == io_state_in_2 ? 8'hfb : _GEN_610; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_612 = 8'h64 == io_state_in_2 ? 8'h43 : _GEN_611; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_613 = 8'h65 == io_state_in_2 ? 8'h4d : _GEN_612; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_614 = 8'h66 == io_state_in_2 ? 8'h33 : _GEN_613; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_615 = 8'h67 == io_state_in_2 ? 8'h85 : _GEN_614; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_616 = 8'h68 == io_state_in_2 ? 8'h45 : _GEN_615; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_617 = 8'h69 == io_state_in_2 ? 8'hf9 : _GEN_616; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_618 = 8'h6a == io_state_in_2 ? 8'h2 : _GEN_617; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_619 = 8'h6b == io_state_in_2 ? 8'h7f : _GEN_618; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_620 = 8'h6c == io_state_in_2 ? 8'h50 : _GEN_619; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_621 = 8'h6d == io_state_in_2 ? 8'h3c : _GEN_620; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_622 = 8'h6e == io_state_in_2 ? 8'h9f : _GEN_621; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_623 = 8'h6f == io_state_in_2 ? 8'ha8 : _GEN_622; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_624 = 8'h70 == io_state_in_2 ? 8'h51 : _GEN_623; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_625 = 8'h71 == io_state_in_2 ? 8'ha3 : _GEN_624; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_626 = 8'h72 == io_state_in_2 ? 8'h40 : _GEN_625; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_627 = 8'h73 == io_state_in_2 ? 8'h8f : _GEN_626; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_628 = 8'h74 == io_state_in_2 ? 8'h92 : _GEN_627; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_629 = 8'h75 == io_state_in_2 ? 8'h9d : _GEN_628; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_630 = 8'h76 == io_state_in_2 ? 8'h38 : _GEN_629; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_631 = 8'h77 == io_state_in_2 ? 8'hf5 : _GEN_630; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_632 = 8'h78 == io_state_in_2 ? 8'hbc : _GEN_631; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_633 = 8'h79 == io_state_in_2 ? 8'hb6 : _GEN_632; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_634 = 8'h7a == io_state_in_2 ? 8'hda : _GEN_633; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_635 = 8'h7b == io_state_in_2 ? 8'h21 : _GEN_634; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_636 = 8'h7c == io_state_in_2 ? 8'h10 : _GEN_635; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_637 = 8'h7d == io_state_in_2 ? 8'hff : _GEN_636; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_638 = 8'h7e == io_state_in_2 ? 8'hf3 : _GEN_637; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_639 = 8'h7f == io_state_in_2 ? 8'hd2 : _GEN_638; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_640 = 8'h80 == io_state_in_2 ? 8'hcd : _GEN_639; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_641 = 8'h81 == io_state_in_2 ? 8'hc : _GEN_640; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_642 = 8'h82 == io_state_in_2 ? 8'h13 : _GEN_641; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_643 = 8'h83 == io_state_in_2 ? 8'hec : _GEN_642; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_644 = 8'h84 == io_state_in_2 ? 8'h5f : _GEN_643; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_645 = 8'h85 == io_state_in_2 ? 8'h97 : _GEN_644; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_646 = 8'h86 == io_state_in_2 ? 8'h44 : _GEN_645; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_647 = 8'h87 == io_state_in_2 ? 8'h17 : _GEN_646; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_648 = 8'h88 == io_state_in_2 ? 8'hc4 : _GEN_647; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_649 = 8'h89 == io_state_in_2 ? 8'ha7 : _GEN_648; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_650 = 8'h8a == io_state_in_2 ? 8'h7e : _GEN_649; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_651 = 8'h8b == io_state_in_2 ? 8'h3d : _GEN_650; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_652 = 8'h8c == io_state_in_2 ? 8'h64 : _GEN_651; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_653 = 8'h8d == io_state_in_2 ? 8'h5d : _GEN_652; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_654 = 8'h8e == io_state_in_2 ? 8'h19 : _GEN_653; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_655 = 8'h8f == io_state_in_2 ? 8'h73 : _GEN_654; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_656 = 8'h90 == io_state_in_2 ? 8'h60 : _GEN_655; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_657 = 8'h91 == io_state_in_2 ? 8'h81 : _GEN_656; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_658 = 8'h92 == io_state_in_2 ? 8'h4f : _GEN_657; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_659 = 8'h93 == io_state_in_2 ? 8'hdc : _GEN_658; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_660 = 8'h94 == io_state_in_2 ? 8'h22 : _GEN_659; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_661 = 8'h95 == io_state_in_2 ? 8'h2a : _GEN_660; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_662 = 8'h96 == io_state_in_2 ? 8'h90 : _GEN_661; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_663 = 8'h97 == io_state_in_2 ? 8'h88 : _GEN_662; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_664 = 8'h98 == io_state_in_2 ? 8'h46 : _GEN_663; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_665 = 8'h99 == io_state_in_2 ? 8'hee : _GEN_664; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_666 = 8'h9a == io_state_in_2 ? 8'hb8 : _GEN_665; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_667 = 8'h9b == io_state_in_2 ? 8'h14 : _GEN_666; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_668 = 8'h9c == io_state_in_2 ? 8'hde : _GEN_667; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_669 = 8'h9d == io_state_in_2 ? 8'h5e : _GEN_668; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_670 = 8'h9e == io_state_in_2 ? 8'hb : _GEN_669; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_671 = 8'h9f == io_state_in_2 ? 8'hdb : _GEN_670; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_672 = 8'ha0 == io_state_in_2 ? 8'he0 : _GEN_671; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_673 = 8'ha1 == io_state_in_2 ? 8'h32 : _GEN_672; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_674 = 8'ha2 == io_state_in_2 ? 8'h3a : _GEN_673; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_675 = 8'ha3 == io_state_in_2 ? 8'ha : _GEN_674; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_676 = 8'ha4 == io_state_in_2 ? 8'h49 : _GEN_675; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_677 = 8'ha5 == io_state_in_2 ? 8'h6 : _GEN_676; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_678 = 8'ha6 == io_state_in_2 ? 8'h24 : _GEN_677; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_679 = 8'ha7 == io_state_in_2 ? 8'h5c : _GEN_678; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_680 = 8'ha8 == io_state_in_2 ? 8'hc2 : _GEN_679; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_681 = 8'ha9 == io_state_in_2 ? 8'hd3 : _GEN_680; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_682 = 8'haa == io_state_in_2 ? 8'hac : _GEN_681; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_683 = 8'hab == io_state_in_2 ? 8'h62 : _GEN_682; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_684 = 8'hac == io_state_in_2 ? 8'h91 : _GEN_683; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_685 = 8'had == io_state_in_2 ? 8'h95 : _GEN_684; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_686 = 8'hae == io_state_in_2 ? 8'he4 : _GEN_685; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_687 = 8'haf == io_state_in_2 ? 8'h79 : _GEN_686; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_688 = 8'hb0 == io_state_in_2 ? 8'he7 : _GEN_687; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_689 = 8'hb1 == io_state_in_2 ? 8'hc8 : _GEN_688; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_690 = 8'hb2 == io_state_in_2 ? 8'h37 : _GEN_689; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_691 = 8'hb3 == io_state_in_2 ? 8'h6d : _GEN_690; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_692 = 8'hb4 == io_state_in_2 ? 8'h8d : _GEN_691; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_693 = 8'hb5 == io_state_in_2 ? 8'hd5 : _GEN_692; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_694 = 8'hb6 == io_state_in_2 ? 8'h4e : _GEN_693; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_695 = 8'hb7 == io_state_in_2 ? 8'ha9 : _GEN_694; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_696 = 8'hb8 == io_state_in_2 ? 8'h6c : _GEN_695; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_697 = 8'hb9 == io_state_in_2 ? 8'h56 : _GEN_696; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_698 = 8'hba == io_state_in_2 ? 8'hf4 : _GEN_697; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_699 = 8'hbb == io_state_in_2 ? 8'hea : _GEN_698; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_700 = 8'hbc == io_state_in_2 ? 8'h65 : _GEN_699; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_701 = 8'hbd == io_state_in_2 ? 8'h7a : _GEN_700; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_702 = 8'hbe == io_state_in_2 ? 8'hae : _GEN_701; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_703 = 8'hbf == io_state_in_2 ? 8'h8 : _GEN_702; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_704 = 8'hc0 == io_state_in_2 ? 8'hba : _GEN_703; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_705 = 8'hc1 == io_state_in_2 ? 8'h78 : _GEN_704; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_706 = 8'hc2 == io_state_in_2 ? 8'h25 : _GEN_705; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_707 = 8'hc3 == io_state_in_2 ? 8'h2e : _GEN_706; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_708 = 8'hc4 == io_state_in_2 ? 8'h1c : _GEN_707; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_709 = 8'hc5 == io_state_in_2 ? 8'ha6 : _GEN_708; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_710 = 8'hc6 == io_state_in_2 ? 8'hb4 : _GEN_709; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_711 = 8'hc7 == io_state_in_2 ? 8'hc6 : _GEN_710; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_712 = 8'hc8 == io_state_in_2 ? 8'he8 : _GEN_711; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_713 = 8'hc9 == io_state_in_2 ? 8'hdd : _GEN_712; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_714 = 8'hca == io_state_in_2 ? 8'h74 : _GEN_713; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_715 = 8'hcb == io_state_in_2 ? 8'h1f : _GEN_714; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_716 = 8'hcc == io_state_in_2 ? 8'h4b : _GEN_715; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_717 = 8'hcd == io_state_in_2 ? 8'hbd : _GEN_716; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_718 = 8'hce == io_state_in_2 ? 8'h8b : _GEN_717; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_719 = 8'hcf == io_state_in_2 ? 8'h8a : _GEN_718; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_720 = 8'hd0 == io_state_in_2 ? 8'h70 : _GEN_719; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_721 = 8'hd1 == io_state_in_2 ? 8'h3e : _GEN_720; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_722 = 8'hd2 == io_state_in_2 ? 8'hb5 : _GEN_721; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_723 = 8'hd3 == io_state_in_2 ? 8'h66 : _GEN_722; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_724 = 8'hd4 == io_state_in_2 ? 8'h48 : _GEN_723; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_725 = 8'hd5 == io_state_in_2 ? 8'h3 : _GEN_724; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_726 = 8'hd6 == io_state_in_2 ? 8'hf6 : _GEN_725; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_727 = 8'hd7 == io_state_in_2 ? 8'he : _GEN_726; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_728 = 8'hd8 == io_state_in_2 ? 8'h61 : _GEN_727; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_729 = 8'hd9 == io_state_in_2 ? 8'h35 : _GEN_728; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_730 = 8'hda == io_state_in_2 ? 8'h57 : _GEN_729; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_731 = 8'hdb == io_state_in_2 ? 8'hb9 : _GEN_730; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_732 = 8'hdc == io_state_in_2 ? 8'h86 : _GEN_731; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_733 = 8'hdd == io_state_in_2 ? 8'hc1 : _GEN_732; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_734 = 8'hde == io_state_in_2 ? 8'h1d : _GEN_733; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_735 = 8'hdf == io_state_in_2 ? 8'h9e : _GEN_734; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_736 = 8'he0 == io_state_in_2 ? 8'he1 : _GEN_735; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_737 = 8'he1 == io_state_in_2 ? 8'hf8 : _GEN_736; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_738 = 8'he2 == io_state_in_2 ? 8'h98 : _GEN_737; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_739 = 8'he3 == io_state_in_2 ? 8'h11 : _GEN_738; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_740 = 8'he4 == io_state_in_2 ? 8'h69 : _GEN_739; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_741 = 8'he5 == io_state_in_2 ? 8'hd9 : _GEN_740; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_742 = 8'he6 == io_state_in_2 ? 8'h8e : _GEN_741; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_743 = 8'he7 == io_state_in_2 ? 8'h94 : _GEN_742; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_744 = 8'he8 == io_state_in_2 ? 8'h9b : _GEN_743; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_745 = 8'he9 == io_state_in_2 ? 8'h1e : _GEN_744; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_746 = 8'hea == io_state_in_2 ? 8'h87 : _GEN_745; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_747 = 8'heb == io_state_in_2 ? 8'he9 : _GEN_746; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_748 = 8'hec == io_state_in_2 ? 8'hce : _GEN_747; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_749 = 8'hed == io_state_in_2 ? 8'h55 : _GEN_748; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_750 = 8'hee == io_state_in_2 ? 8'h28 : _GEN_749; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_751 = 8'hef == io_state_in_2 ? 8'hdf : _GEN_750; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_752 = 8'hf0 == io_state_in_2 ? 8'h8c : _GEN_751; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_753 = 8'hf1 == io_state_in_2 ? 8'ha1 : _GEN_752; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_754 = 8'hf2 == io_state_in_2 ? 8'h89 : _GEN_753; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_755 = 8'hf3 == io_state_in_2 ? 8'hd : _GEN_754; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_756 = 8'hf4 == io_state_in_2 ? 8'hbf : _GEN_755; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_757 = 8'hf5 == io_state_in_2 ? 8'he6 : _GEN_756; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_758 = 8'hf6 == io_state_in_2 ? 8'h42 : _GEN_757; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_759 = 8'hf7 == io_state_in_2 ? 8'h68 : _GEN_758; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_760 = 8'hf8 == io_state_in_2 ? 8'h41 : _GEN_759; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_761 = 8'hf9 == io_state_in_2 ? 8'h99 : _GEN_760; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_762 = 8'hfa == io_state_in_2 ? 8'h2d : _GEN_761; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_763 = 8'hfb == io_state_in_2 ? 8'hf : _GEN_762; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_764 = 8'hfc == io_state_in_2 ? 8'hb0 : _GEN_763; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_765 = 8'hfd == io_state_in_2 ? 8'h54 : _GEN_764; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_766 = 8'hfe == io_state_in_2 ? 8'hbb : _GEN_765; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_769 = 8'h1 == io_state_in_3 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_770 = 8'h2 == io_state_in_3 ? 8'h77 : _GEN_769; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_771 = 8'h3 == io_state_in_3 ? 8'h7b : _GEN_770; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_772 = 8'h4 == io_state_in_3 ? 8'hf2 : _GEN_771; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_773 = 8'h5 == io_state_in_3 ? 8'h6b : _GEN_772; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_774 = 8'h6 == io_state_in_3 ? 8'h6f : _GEN_773; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_775 = 8'h7 == io_state_in_3 ? 8'hc5 : _GEN_774; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_776 = 8'h8 == io_state_in_3 ? 8'h30 : _GEN_775; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_777 = 8'h9 == io_state_in_3 ? 8'h1 : _GEN_776; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_778 = 8'ha == io_state_in_3 ? 8'h67 : _GEN_777; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_779 = 8'hb == io_state_in_3 ? 8'h2b : _GEN_778; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_780 = 8'hc == io_state_in_3 ? 8'hfe : _GEN_779; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_781 = 8'hd == io_state_in_3 ? 8'hd7 : _GEN_780; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_782 = 8'he == io_state_in_3 ? 8'hab : _GEN_781; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_783 = 8'hf == io_state_in_3 ? 8'h76 : _GEN_782; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_784 = 8'h10 == io_state_in_3 ? 8'hca : _GEN_783; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_785 = 8'h11 == io_state_in_3 ? 8'h82 : _GEN_784; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_786 = 8'h12 == io_state_in_3 ? 8'hc9 : _GEN_785; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_787 = 8'h13 == io_state_in_3 ? 8'h7d : _GEN_786; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_788 = 8'h14 == io_state_in_3 ? 8'hfa : _GEN_787; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_789 = 8'h15 == io_state_in_3 ? 8'h59 : _GEN_788; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_790 = 8'h16 == io_state_in_3 ? 8'h47 : _GEN_789; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_791 = 8'h17 == io_state_in_3 ? 8'hf0 : _GEN_790; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_792 = 8'h18 == io_state_in_3 ? 8'had : _GEN_791; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_793 = 8'h19 == io_state_in_3 ? 8'hd4 : _GEN_792; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_794 = 8'h1a == io_state_in_3 ? 8'ha2 : _GEN_793; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_795 = 8'h1b == io_state_in_3 ? 8'haf : _GEN_794; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_796 = 8'h1c == io_state_in_3 ? 8'h9c : _GEN_795; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_797 = 8'h1d == io_state_in_3 ? 8'ha4 : _GEN_796; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_798 = 8'h1e == io_state_in_3 ? 8'h72 : _GEN_797; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_799 = 8'h1f == io_state_in_3 ? 8'hc0 : _GEN_798; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_800 = 8'h20 == io_state_in_3 ? 8'hb7 : _GEN_799; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_801 = 8'h21 == io_state_in_3 ? 8'hfd : _GEN_800; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_802 = 8'h22 == io_state_in_3 ? 8'h93 : _GEN_801; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_803 = 8'h23 == io_state_in_3 ? 8'h26 : _GEN_802; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_804 = 8'h24 == io_state_in_3 ? 8'h36 : _GEN_803; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_805 = 8'h25 == io_state_in_3 ? 8'h3f : _GEN_804; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_806 = 8'h26 == io_state_in_3 ? 8'hf7 : _GEN_805; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_807 = 8'h27 == io_state_in_3 ? 8'hcc : _GEN_806; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_808 = 8'h28 == io_state_in_3 ? 8'h34 : _GEN_807; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_809 = 8'h29 == io_state_in_3 ? 8'ha5 : _GEN_808; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_810 = 8'h2a == io_state_in_3 ? 8'he5 : _GEN_809; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_811 = 8'h2b == io_state_in_3 ? 8'hf1 : _GEN_810; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_812 = 8'h2c == io_state_in_3 ? 8'h71 : _GEN_811; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_813 = 8'h2d == io_state_in_3 ? 8'hd8 : _GEN_812; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_814 = 8'h2e == io_state_in_3 ? 8'h31 : _GEN_813; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_815 = 8'h2f == io_state_in_3 ? 8'h15 : _GEN_814; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_816 = 8'h30 == io_state_in_3 ? 8'h4 : _GEN_815; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_817 = 8'h31 == io_state_in_3 ? 8'hc7 : _GEN_816; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_818 = 8'h32 == io_state_in_3 ? 8'h23 : _GEN_817; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_819 = 8'h33 == io_state_in_3 ? 8'hc3 : _GEN_818; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_820 = 8'h34 == io_state_in_3 ? 8'h18 : _GEN_819; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_821 = 8'h35 == io_state_in_3 ? 8'h96 : _GEN_820; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_822 = 8'h36 == io_state_in_3 ? 8'h5 : _GEN_821; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_823 = 8'h37 == io_state_in_3 ? 8'h9a : _GEN_822; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_824 = 8'h38 == io_state_in_3 ? 8'h7 : _GEN_823; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_825 = 8'h39 == io_state_in_3 ? 8'h12 : _GEN_824; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_826 = 8'h3a == io_state_in_3 ? 8'h80 : _GEN_825; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_827 = 8'h3b == io_state_in_3 ? 8'he2 : _GEN_826; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_828 = 8'h3c == io_state_in_3 ? 8'heb : _GEN_827; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_829 = 8'h3d == io_state_in_3 ? 8'h27 : _GEN_828; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_830 = 8'h3e == io_state_in_3 ? 8'hb2 : _GEN_829; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_831 = 8'h3f == io_state_in_3 ? 8'h75 : _GEN_830; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_832 = 8'h40 == io_state_in_3 ? 8'h9 : _GEN_831; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_833 = 8'h41 == io_state_in_3 ? 8'h83 : _GEN_832; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_834 = 8'h42 == io_state_in_3 ? 8'h2c : _GEN_833; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_835 = 8'h43 == io_state_in_3 ? 8'h1a : _GEN_834; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_836 = 8'h44 == io_state_in_3 ? 8'h1b : _GEN_835; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_837 = 8'h45 == io_state_in_3 ? 8'h6e : _GEN_836; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_838 = 8'h46 == io_state_in_3 ? 8'h5a : _GEN_837; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_839 = 8'h47 == io_state_in_3 ? 8'ha0 : _GEN_838; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_840 = 8'h48 == io_state_in_3 ? 8'h52 : _GEN_839; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_841 = 8'h49 == io_state_in_3 ? 8'h3b : _GEN_840; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_842 = 8'h4a == io_state_in_3 ? 8'hd6 : _GEN_841; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_843 = 8'h4b == io_state_in_3 ? 8'hb3 : _GEN_842; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_844 = 8'h4c == io_state_in_3 ? 8'h29 : _GEN_843; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_845 = 8'h4d == io_state_in_3 ? 8'he3 : _GEN_844; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_846 = 8'h4e == io_state_in_3 ? 8'h2f : _GEN_845; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_847 = 8'h4f == io_state_in_3 ? 8'h84 : _GEN_846; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_848 = 8'h50 == io_state_in_3 ? 8'h53 : _GEN_847; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_849 = 8'h51 == io_state_in_3 ? 8'hd1 : _GEN_848; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_850 = 8'h52 == io_state_in_3 ? 8'h0 : _GEN_849; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_851 = 8'h53 == io_state_in_3 ? 8'hed : _GEN_850; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_852 = 8'h54 == io_state_in_3 ? 8'h20 : _GEN_851; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_853 = 8'h55 == io_state_in_3 ? 8'hfc : _GEN_852; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_854 = 8'h56 == io_state_in_3 ? 8'hb1 : _GEN_853; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_855 = 8'h57 == io_state_in_3 ? 8'h5b : _GEN_854; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_856 = 8'h58 == io_state_in_3 ? 8'h6a : _GEN_855; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_857 = 8'h59 == io_state_in_3 ? 8'hcb : _GEN_856; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_858 = 8'h5a == io_state_in_3 ? 8'hbe : _GEN_857; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_859 = 8'h5b == io_state_in_3 ? 8'h39 : _GEN_858; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_860 = 8'h5c == io_state_in_3 ? 8'h4a : _GEN_859; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_861 = 8'h5d == io_state_in_3 ? 8'h4c : _GEN_860; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_862 = 8'h5e == io_state_in_3 ? 8'h58 : _GEN_861; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_863 = 8'h5f == io_state_in_3 ? 8'hcf : _GEN_862; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_864 = 8'h60 == io_state_in_3 ? 8'hd0 : _GEN_863; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_865 = 8'h61 == io_state_in_3 ? 8'hef : _GEN_864; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_866 = 8'h62 == io_state_in_3 ? 8'haa : _GEN_865; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_867 = 8'h63 == io_state_in_3 ? 8'hfb : _GEN_866; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_868 = 8'h64 == io_state_in_3 ? 8'h43 : _GEN_867; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_869 = 8'h65 == io_state_in_3 ? 8'h4d : _GEN_868; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_870 = 8'h66 == io_state_in_3 ? 8'h33 : _GEN_869; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_871 = 8'h67 == io_state_in_3 ? 8'h85 : _GEN_870; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_872 = 8'h68 == io_state_in_3 ? 8'h45 : _GEN_871; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_873 = 8'h69 == io_state_in_3 ? 8'hf9 : _GEN_872; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_874 = 8'h6a == io_state_in_3 ? 8'h2 : _GEN_873; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_875 = 8'h6b == io_state_in_3 ? 8'h7f : _GEN_874; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_876 = 8'h6c == io_state_in_3 ? 8'h50 : _GEN_875; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_877 = 8'h6d == io_state_in_3 ? 8'h3c : _GEN_876; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_878 = 8'h6e == io_state_in_3 ? 8'h9f : _GEN_877; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_879 = 8'h6f == io_state_in_3 ? 8'ha8 : _GEN_878; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_880 = 8'h70 == io_state_in_3 ? 8'h51 : _GEN_879; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_881 = 8'h71 == io_state_in_3 ? 8'ha3 : _GEN_880; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_882 = 8'h72 == io_state_in_3 ? 8'h40 : _GEN_881; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_883 = 8'h73 == io_state_in_3 ? 8'h8f : _GEN_882; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_884 = 8'h74 == io_state_in_3 ? 8'h92 : _GEN_883; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_885 = 8'h75 == io_state_in_3 ? 8'h9d : _GEN_884; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_886 = 8'h76 == io_state_in_3 ? 8'h38 : _GEN_885; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_887 = 8'h77 == io_state_in_3 ? 8'hf5 : _GEN_886; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_888 = 8'h78 == io_state_in_3 ? 8'hbc : _GEN_887; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_889 = 8'h79 == io_state_in_3 ? 8'hb6 : _GEN_888; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_890 = 8'h7a == io_state_in_3 ? 8'hda : _GEN_889; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_891 = 8'h7b == io_state_in_3 ? 8'h21 : _GEN_890; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_892 = 8'h7c == io_state_in_3 ? 8'h10 : _GEN_891; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_893 = 8'h7d == io_state_in_3 ? 8'hff : _GEN_892; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_894 = 8'h7e == io_state_in_3 ? 8'hf3 : _GEN_893; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_895 = 8'h7f == io_state_in_3 ? 8'hd2 : _GEN_894; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_896 = 8'h80 == io_state_in_3 ? 8'hcd : _GEN_895; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_897 = 8'h81 == io_state_in_3 ? 8'hc : _GEN_896; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_898 = 8'h82 == io_state_in_3 ? 8'h13 : _GEN_897; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_899 = 8'h83 == io_state_in_3 ? 8'hec : _GEN_898; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_900 = 8'h84 == io_state_in_3 ? 8'h5f : _GEN_899; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_901 = 8'h85 == io_state_in_3 ? 8'h97 : _GEN_900; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_902 = 8'h86 == io_state_in_3 ? 8'h44 : _GEN_901; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_903 = 8'h87 == io_state_in_3 ? 8'h17 : _GEN_902; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_904 = 8'h88 == io_state_in_3 ? 8'hc4 : _GEN_903; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_905 = 8'h89 == io_state_in_3 ? 8'ha7 : _GEN_904; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_906 = 8'h8a == io_state_in_3 ? 8'h7e : _GEN_905; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_907 = 8'h8b == io_state_in_3 ? 8'h3d : _GEN_906; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_908 = 8'h8c == io_state_in_3 ? 8'h64 : _GEN_907; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_909 = 8'h8d == io_state_in_3 ? 8'h5d : _GEN_908; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_910 = 8'h8e == io_state_in_3 ? 8'h19 : _GEN_909; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_911 = 8'h8f == io_state_in_3 ? 8'h73 : _GEN_910; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_912 = 8'h90 == io_state_in_3 ? 8'h60 : _GEN_911; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_913 = 8'h91 == io_state_in_3 ? 8'h81 : _GEN_912; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_914 = 8'h92 == io_state_in_3 ? 8'h4f : _GEN_913; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_915 = 8'h93 == io_state_in_3 ? 8'hdc : _GEN_914; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_916 = 8'h94 == io_state_in_3 ? 8'h22 : _GEN_915; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_917 = 8'h95 == io_state_in_3 ? 8'h2a : _GEN_916; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_918 = 8'h96 == io_state_in_3 ? 8'h90 : _GEN_917; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_919 = 8'h97 == io_state_in_3 ? 8'h88 : _GEN_918; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_920 = 8'h98 == io_state_in_3 ? 8'h46 : _GEN_919; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_921 = 8'h99 == io_state_in_3 ? 8'hee : _GEN_920; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_922 = 8'h9a == io_state_in_3 ? 8'hb8 : _GEN_921; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_923 = 8'h9b == io_state_in_3 ? 8'h14 : _GEN_922; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_924 = 8'h9c == io_state_in_3 ? 8'hde : _GEN_923; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_925 = 8'h9d == io_state_in_3 ? 8'h5e : _GEN_924; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_926 = 8'h9e == io_state_in_3 ? 8'hb : _GEN_925; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_927 = 8'h9f == io_state_in_3 ? 8'hdb : _GEN_926; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_928 = 8'ha0 == io_state_in_3 ? 8'he0 : _GEN_927; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_929 = 8'ha1 == io_state_in_3 ? 8'h32 : _GEN_928; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_930 = 8'ha2 == io_state_in_3 ? 8'h3a : _GEN_929; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_931 = 8'ha3 == io_state_in_3 ? 8'ha : _GEN_930; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_932 = 8'ha4 == io_state_in_3 ? 8'h49 : _GEN_931; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_933 = 8'ha5 == io_state_in_3 ? 8'h6 : _GEN_932; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_934 = 8'ha6 == io_state_in_3 ? 8'h24 : _GEN_933; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_935 = 8'ha7 == io_state_in_3 ? 8'h5c : _GEN_934; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_936 = 8'ha8 == io_state_in_3 ? 8'hc2 : _GEN_935; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_937 = 8'ha9 == io_state_in_3 ? 8'hd3 : _GEN_936; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_938 = 8'haa == io_state_in_3 ? 8'hac : _GEN_937; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_939 = 8'hab == io_state_in_3 ? 8'h62 : _GEN_938; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_940 = 8'hac == io_state_in_3 ? 8'h91 : _GEN_939; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_941 = 8'had == io_state_in_3 ? 8'h95 : _GEN_940; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_942 = 8'hae == io_state_in_3 ? 8'he4 : _GEN_941; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_943 = 8'haf == io_state_in_3 ? 8'h79 : _GEN_942; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_944 = 8'hb0 == io_state_in_3 ? 8'he7 : _GEN_943; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_945 = 8'hb1 == io_state_in_3 ? 8'hc8 : _GEN_944; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_946 = 8'hb2 == io_state_in_3 ? 8'h37 : _GEN_945; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_947 = 8'hb3 == io_state_in_3 ? 8'h6d : _GEN_946; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_948 = 8'hb4 == io_state_in_3 ? 8'h8d : _GEN_947; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_949 = 8'hb5 == io_state_in_3 ? 8'hd5 : _GEN_948; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_950 = 8'hb6 == io_state_in_3 ? 8'h4e : _GEN_949; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_951 = 8'hb7 == io_state_in_3 ? 8'ha9 : _GEN_950; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_952 = 8'hb8 == io_state_in_3 ? 8'h6c : _GEN_951; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_953 = 8'hb9 == io_state_in_3 ? 8'h56 : _GEN_952; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_954 = 8'hba == io_state_in_3 ? 8'hf4 : _GEN_953; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_955 = 8'hbb == io_state_in_3 ? 8'hea : _GEN_954; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_956 = 8'hbc == io_state_in_3 ? 8'h65 : _GEN_955; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_957 = 8'hbd == io_state_in_3 ? 8'h7a : _GEN_956; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_958 = 8'hbe == io_state_in_3 ? 8'hae : _GEN_957; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_959 = 8'hbf == io_state_in_3 ? 8'h8 : _GEN_958; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_960 = 8'hc0 == io_state_in_3 ? 8'hba : _GEN_959; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_961 = 8'hc1 == io_state_in_3 ? 8'h78 : _GEN_960; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_962 = 8'hc2 == io_state_in_3 ? 8'h25 : _GEN_961; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_963 = 8'hc3 == io_state_in_3 ? 8'h2e : _GEN_962; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_964 = 8'hc4 == io_state_in_3 ? 8'h1c : _GEN_963; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_965 = 8'hc5 == io_state_in_3 ? 8'ha6 : _GEN_964; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_966 = 8'hc6 == io_state_in_3 ? 8'hb4 : _GEN_965; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_967 = 8'hc7 == io_state_in_3 ? 8'hc6 : _GEN_966; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_968 = 8'hc8 == io_state_in_3 ? 8'he8 : _GEN_967; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_969 = 8'hc9 == io_state_in_3 ? 8'hdd : _GEN_968; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_970 = 8'hca == io_state_in_3 ? 8'h74 : _GEN_969; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_971 = 8'hcb == io_state_in_3 ? 8'h1f : _GEN_970; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_972 = 8'hcc == io_state_in_3 ? 8'h4b : _GEN_971; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_973 = 8'hcd == io_state_in_3 ? 8'hbd : _GEN_972; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_974 = 8'hce == io_state_in_3 ? 8'h8b : _GEN_973; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_975 = 8'hcf == io_state_in_3 ? 8'h8a : _GEN_974; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_976 = 8'hd0 == io_state_in_3 ? 8'h70 : _GEN_975; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_977 = 8'hd1 == io_state_in_3 ? 8'h3e : _GEN_976; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_978 = 8'hd2 == io_state_in_3 ? 8'hb5 : _GEN_977; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_979 = 8'hd3 == io_state_in_3 ? 8'h66 : _GEN_978; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_980 = 8'hd4 == io_state_in_3 ? 8'h48 : _GEN_979; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_981 = 8'hd5 == io_state_in_3 ? 8'h3 : _GEN_980; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_982 = 8'hd6 == io_state_in_3 ? 8'hf6 : _GEN_981; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_983 = 8'hd7 == io_state_in_3 ? 8'he : _GEN_982; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_984 = 8'hd8 == io_state_in_3 ? 8'h61 : _GEN_983; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_985 = 8'hd9 == io_state_in_3 ? 8'h35 : _GEN_984; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_986 = 8'hda == io_state_in_3 ? 8'h57 : _GEN_985; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_987 = 8'hdb == io_state_in_3 ? 8'hb9 : _GEN_986; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_988 = 8'hdc == io_state_in_3 ? 8'h86 : _GEN_987; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_989 = 8'hdd == io_state_in_3 ? 8'hc1 : _GEN_988; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_990 = 8'hde == io_state_in_3 ? 8'h1d : _GEN_989; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_991 = 8'hdf == io_state_in_3 ? 8'h9e : _GEN_990; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_992 = 8'he0 == io_state_in_3 ? 8'he1 : _GEN_991; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_993 = 8'he1 == io_state_in_3 ? 8'hf8 : _GEN_992; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_994 = 8'he2 == io_state_in_3 ? 8'h98 : _GEN_993; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_995 = 8'he3 == io_state_in_3 ? 8'h11 : _GEN_994; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_996 = 8'he4 == io_state_in_3 ? 8'h69 : _GEN_995; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_997 = 8'he5 == io_state_in_3 ? 8'hd9 : _GEN_996; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_998 = 8'he6 == io_state_in_3 ? 8'h8e : _GEN_997; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_999 = 8'he7 == io_state_in_3 ? 8'h94 : _GEN_998; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1000 = 8'he8 == io_state_in_3 ? 8'h9b : _GEN_999; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1001 = 8'he9 == io_state_in_3 ? 8'h1e : _GEN_1000; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1002 = 8'hea == io_state_in_3 ? 8'h87 : _GEN_1001; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1003 = 8'heb == io_state_in_3 ? 8'he9 : _GEN_1002; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1004 = 8'hec == io_state_in_3 ? 8'hce : _GEN_1003; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1005 = 8'hed == io_state_in_3 ? 8'h55 : _GEN_1004; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1006 = 8'hee == io_state_in_3 ? 8'h28 : _GEN_1005; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1007 = 8'hef == io_state_in_3 ? 8'hdf : _GEN_1006; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1008 = 8'hf0 == io_state_in_3 ? 8'h8c : _GEN_1007; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1009 = 8'hf1 == io_state_in_3 ? 8'ha1 : _GEN_1008; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1010 = 8'hf2 == io_state_in_3 ? 8'h89 : _GEN_1009; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1011 = 8'hf3 == io_state_in_3 ? 8'hd : _GEN_1010; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1012 = 8'hf4 == io_state_in_3 ? 8'hbf : _GEN_1011; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1013 = 8'hf5 == io_state_in_3 ? 8'he6 : _GEN_1012; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1014 = 8'hf6 == io_state_in_3 ? 8'h42 : _GEN_1013; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1015 = 8'hf7 == io_state_in_3 ? 8'h68 : _GEN_1014; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1016 = 8'hf8 == io_state_in_3 ? 8'h41 : _GEN_1015; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1017 = 8'hf9 == io_state_in_3 ? 8'h99 : _GEN_1016; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1018 = 8'hfa == io_state_in_3 ? 8'h2d : _GEN_1017; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1019 = 8'hfb == io_state_in_3 ? 8'hf : _GEN_1018; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1020 = 8'hfc == io_state_in_3 ? 8'hb0 : _GEN_1019; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1021 = 8'hfd == io_state_in_3 ? 8'h54 : _GEN_1020; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1022 = 8'hfe == io_state_in_3 ? 8'hbb : _GEN_1021; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1025 = 8'h1 == io_state_in_4 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1026 = 8'h2 == io_state_in_4 ? 8'h77 : _GEN_1025; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1027 = 8'h3 == io_state_in_4 ? 8'h7b : _GEN_1026; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1028 = 8'h4 == io_state_in_4 ? 8'hf2 : _GEN_1027; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1029 = 8'h5 == io_state_in_4 ? 8'h6b : _GEN_1028; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1030 = 8'h6 == io_state_in_4 ? 8'h6f : _GEN_1029; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1031 = 8'h7 == io_state_in_4 ? 8'hc5 : _GEN_1030; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1032 = 8'h8 == io_state_in_4 ? 8'h30 : _GEN_1031; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1033 = 8'h9 == io_state_in_4 ? 8'h1 : _GEN_1032; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1034 = 8'ha == io_state_in_4 ? 8'h67 : _GEN_1033; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1035 = 8'hb == io_state_in_4 ? 8'h2b : _GEN_1034; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1036 = 8'hc == io_state_in_4 ? 8'hfe : _GEN_1035; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1037 = 8'hd == io_state_in_4 ? 8'hd7 : _GEN_1036; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1038 = 8'he == io_state_in_4 ? 8'hab : _GEN_1037; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1039 = 8'hf == io_state_in_4 ? 8'h76 : _GEN_1038; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1040 = 8'h10 == io_state_in_4 ? 8'hca : _GEN_1039; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1041 = 8'h11 == io_state_in_4 ? 8'h82 : _GEN_1040; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1042 = 8'h12 == io_state_in_4 ? 8'hc9 : _GEN_1041; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1043 = 8'h13 == io_state_in_4 ? 8'h7d : _GEN_1042; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1044 = 8'h14 == io_state_in_4 ? 8'hfa : _GEN_1043; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1045 = 8'h15 == io_state_in_4 ? 8'h59 : _GEN_1044; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1046 = 8'h16 == io_state_in_4 ? 8'h47 : _GEN_1045; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1047 = 8'h17 == io_state_in_4 ? 8'hf0 : _GEN_1046; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1048 = 8'h18 == io_state_in_4 ? 8'had : _GEN_1047; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1049 = 8'h19 == io_state_in_4 ? 8'hd4 : _GEN_1048; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1050 = 8'h1a == io_state_in_4 ? 8'ha2 : _GEN_1049; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1051 = 8'h1b == io_state_in_4 ? 8'haf : _GEN_1050; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1052 = 8'h1c == io_state_in_4 ? 8'h9c : _GEN_1051; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1053 = 8'h1d == io_state_in_4 ? 8'ha4 : _GEN_1052; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1054 = 8'h1e == io_state_in_4 ? 8'h72 : _GEN_1053; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1055 = 8'h1f == io_state_in_4 ? 8'hc0 : _GEN_1054; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1056 = 8'h20 == io_state_in_4 ? 8'hb7 : _GEN_1055; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1057 = 8'h21 == io_state_in_4 ? 8'hfd : _GEN_1056; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1058 = 8'h22 == io_state_in_4 ? 8'h93 : _GEN_1057; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1059 = 8'h23 == io_state_in_4 ? 8'h26 : _GEN_1058; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1060 = 8'h24 == io_state_in_4 ? 8'h36 : _GEN_1059; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1061 = 8'h25 == io_state_in_4 ? 8'h3f : _GEN_1060; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1062 = 8'h26 == io_state_in_4 ? 8'hf7 : _GEN_1061; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1063 = 8'h27 == io_state_in_4 ? 8'hcc : _GEN_1062; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1064 = 8'h28 == io_state_in_4 ? 8'h34 : _GEN_1063; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1065 = 8'h29 == io_state_in_4 ? 8'ha5 : _GEN_1064; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1066 = 8'h2a == io_state_in_4 ? 8'he5 : _GEN_1065; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1067 = 8'h2b == io_state_in_4 ? 8'hf1 : _GEN_1066; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1068 = 8'h2c == io_state_in_4 ? 8'h71 : _GEN_1067; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1069 = 8'h2d == io_state_in_4 ? 8'hd8 : _GEN_1068; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1070 = 8'h2e == io_state_in_4 ? 8'h31 : _GEN_1069; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1071 = 8'h2f == io_state_in_4 ? 8'h15 : _GEN_1070; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1072 = 8'h30 == io_state_in_4 ? 8'h4 : _GEN_1071; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1073 = 8'h31 == io_state_in_4 ? 8'hc7 : _GEN_1072; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1074 = 8'h32 == io_state_in_4 ? 8'h23 : _GEN_1073; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1075 = 8'h33 == io_state_in_4 ? 8'hc3 : _GEN_1074; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1076 = 8'h34 == io_state_in_4 ? 8'h18 : _GEN_1075; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1077 = 8'h35 == io_state_in_4 ? 8'h96 : _GEN_1076; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1078 = 8'h36 == io_state_in_4 ? 8'h5 : _GEN_1077; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1079 = 8'h37 == io_state_in_4 ? 8'h9a : _GEN_1078; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1080 = 8'h38 == io_state_in_4 ? 8'h7 : _GEN_1079; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1081 = 8'h39 == io_state_in_4 ? 8'h12 : _GEN_1080; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1082 = 8'h3a == io_state_in_4 ? 8'h80 : _GEN_1081; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1083 = 8'h3b == io_state_in_4 ? 8'he2 : _GEN_1082; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1084 = 8'h3c == io_state_in_4 ? 8'heb : _GEN_1083; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1085 = 8'h3d == io_state_in_4 ? 8'h27 : _GEN_1084; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1086 = 8'h3e == io_state_in_4 ? 8'hb2 : _GEN_1085; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1087 = 8'h3f == io_state_in_4 ? 8'h75 : _GEN_1086; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1088 = 8'h40 == io_state_in_4 ? 8'h9 : _GEN_1087; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1089 = 8'h41 == io_state_in_4 ? 8'h83 : _GEN_1088; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1090 = 8'h42 == io_state_in_4 ? 8'h2c : _GEN_1089; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1091 = 8'h43 == io_state_in_4 ? 8'h1a : _GEN_1090; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1092 = 8'h44 == io_state_in_4 ? 8'h1b : _GEN_1091; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1093 = 8'h45 == io_state_in_4 ? 8'h6e : _GEN_1092; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1094 = 8'h46 == io_state_in_4 ? 8'h5a : _GEN_1093; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1095 = 8'h47 == io_state_in_4 ? 8'ha0 : _GEN_1094; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1096 = 8'h48 == io_state_in_4 ? 8'h52 : _GEN_1095; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1097 = 8'h49 == io_state_in_4 ? 8'h3b : _GEN_1096; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1098 = 8'h4a == io_state_in_4 ? 8'hd6 : _GEN_1097; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1099 = 8'h4b == io_state_in_4 ? 8'hb3 : _GEN_1098; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1100 = 8'h4c == io_state_in_4 ? 8'h29 : _GEN_1099; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1101 = 8'h4d == io_state_in_4 ? 8'he3 : _GEN_1100; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1102 = 8'h4e == io_state_in_4 ? 8'h2f : _GEN_1101; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1103 = 8'h4f == io_state_in_4 ? 8'h84 : _GEN_1102; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1104 = 8'h50 == io_state_in_4 ? 8'h53 : _GEN_1103; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1105 = 8'h51 == io_state_in_4 ? 8'hd1 : _GEN_1104; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1106 = 8'h52 == io_state_in_4 ? 8'h0 : _GEN_1105; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1107 = 8'h53 == io_state_in_4 ? 8'hed : _GEN_1106; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1108 = 8'h54 == io_state_in_4 ? 8'h20 : _GEN_1107; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1109 = 8'h55 == io_state_in_4 ? 8'hfc : _GEN_1108; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1110 = 8'h56 == io_state_in_4 ? 8'hb1 : _GEN_1109; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1111 = 8'h57 == io_state_in_4 ? 8'h5b : _GEN_1110; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1112 = 8'h58 == io_state_in_4 ? 8'h6a : _GEN_1111; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1113 = 8'h59 == io_state_in_4 ? 8'hcb : _GEN_1112; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1114 = 8'h5a == io_state_in_4 ? 8'hbe : _GEN_1113; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1115 = 8'h5b == io_state_in_4 ? 8'h39 : _GEN_1114; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1116 = 8'h5c == io_state_in_4 ? 8'h4a : _GEN_1115; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1117 = 8'h5d == io_state_in_4 ? 8'h4c : _GEN_1116; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1118 = 8'h5e == io_state_in_4 ? 8'h58 : _GEN_1117; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1119 = 8'h5f == io_state_in_4 ? 8'hcf : _GEN_1118; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1120 = 8'h60 == io_state_in_4 ? 8'hd0 : _GEN_1119; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1121 = 8'h61 == io_state_in_4 ? 8'hef : _GEN_1120; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1122 = 8'h62 == io_state_in_4 ? 8'haa : _GEN_1121; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1123 = 8'h63 == io_state_in_4 ? 8'hfb : _GEN_1122; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1124 = 8'h64 == io_state_in_4 ? 8'h43 : _GEN_1123; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1125 = 8'h65 == io_state_in_4 ? 8'h4d : _GEN_1124; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1126 = 8'h66 == io_state_in_4 ? 8'h33 : _GEN_1125; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1127 = 8'h67 == io_state_in_4 ? 8'h85 : _GEN_1126; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1128 = 8'h68 == io_state_in_4 ? 8'h45 : _GEN_1127; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1129 = 8'h69 == io_state_in_4 ? 8'hf9 : _GEN_1128; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1130 = 8'h6a == io_state_in_4 ? 8'h2 : _GEN_1129; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1131 = 8'h6b == io_state_in_4 ? 8'h7f : _GEN_1130; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1132 = 8'h6c == io_state_in_4 ? 8'h50 : _GEN_1131; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1133 = 8'h6d == io_state_in_4 ? 8'h3c : _GEN_1132; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1134 = 8'h6e == io_state_in_4 ? 8'h9f : _GEN_1133; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1135 = 8'h6f == io_state_in_4 ? 8'ha8 : _GEN_1134; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1136 = 8'h70 == io_state_in_4 ? 8'h51 : _GEN_1135; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1137 = 8'h71 == io_state_in_4 ? 8'ha3 : _GEN_1136; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1138 = 8'h72 == io_state_in_4 ? 8'h40 : _GEN_1137; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1139 = 8'h73 == io_state_in_4 ? 8'h8f : _GEN_1138; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1140 = 8'h74 == io_state_in_4 ? 8'h92 : _GEN_1139; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1141 = 8'h75 == io_state_in_4 ? 8'h9d : _GEN_1140; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1142 = 8'h76 == io_state_in_4 ? 8'h38 : _GEN_1141; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1143 = 8'h77 == io_state_in_4 ? 8'hf5 : _GEN_1142; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1144 = 8'h78 == io_state_in_4 ? 8'hbc : _GEN_1143; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1145 = 8'h79 == io_state_in_4 ? 8'hb6 : _GEN_1144; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1146 = 8'h7a == io_state_in_4 ? 8'hda : _GEN_1145; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1147 = 8'h7b == io_state_in_4 ? 8'h21 : _GEN_1146; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1148 = 8'h7c == io_state_in_4 ? 8'h10 : _GEN_1147; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1149 = 8'h7d == io_state_in_4 ? 8'hff : _GEN_1148; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1150 = 8'h7e == io_state_in_4 ? 8'hf3 : _GEN_1149; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1151 = 8'h7f == io_state_in_4 ? 8'hd2 : _GEN_1150; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1152 = 8'h80 == io_state_in_4 ? 8'hcd : _GEN_1151; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1153 = 8'h81 == io_state_in_4 ? 8'hc : _GEN_1152; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1154 = 8'h82 == io_state_in_4 ? 8'h13 : _GEN_1153; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1155 = 8'h83 == io_state_in_4 ? 8'hec : _GEN_1154; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1156 = 8'h84 == io_state_in_4 ? 8'h5f : _GEN_1155; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1157 = 8'h85 == io_state_in_4 ? 8'h97 : _GEN_1156; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1158 = 8'h86 == io_state_in_4 ? 8'h44 : _GEN_1157; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1159 = 8'h87 == io_state_in_4 ? 8'h17 : _GEN_1158; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1160 = 8'h88 == io_state_in_4 ? 8'hc4 : _GEN_1159; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1161 = 8'h89 == io_state_in_4 ? 8'ha7 : _GEN_1160; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1162 = 8'h8a == io_state_in_4 ? 8'h7e : _GEN_1161; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1163 = 8'h8b == io_state_in_4 ? 8'h3d : _GEN_1162; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1164 = 8'h8c == io_state_in_4 ? 8'h64 : _GEN_1163; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1165 = 8'h8d == io_state_in_4 ? 8'h5d : _GEN_1164; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1166 = 8'h8e == io_state_in_4 ? 8'h19 : _GEN_1165; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1167 = 8'h8f == io_state_in_4 ? 8'h73 : _GEN_1166; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1168 = 8'h90 == io_state_in_4 ? 8'h60 : _GEN_1167; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1169 = 8'h91 == io_state_in_4 ? 8'h81 : _GEN_1168; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1170 = 8'h92 == io_state_in_4 ? 8'h4f : _GEN_1169; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1171 = 8'h93 == io_state_in_4 ? 8'hdc : _GEN_1170; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1172 = 8'h94 == io_state_in_4 ? 8'h22 : _GEN_1171; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1173 = 8'h95 == io_state_in_4 ? 8'h2a : _GEN_1172; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1174 = 8'h96 == io_state_in_4 ? 8'h90 : _GEN_1173; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1175 = 8'h97 == io_state_in_4 ? 8'h88 : _GEN_1174; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1176 = 8'h98 == io_state_in_4 ? 8'h46 : _GEN_1175; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1177 = 8'h99 == io_state_in_4 ? 8'hee : _GEN_1176; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1178 = 8'h9a == io_state_in_4 ? 8'hb8 : _GEN_1177; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1179 = 8'h9b == io_state_in_4 ? 8'h14 : _GEN_1178; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1180 = 8'h9c == io_state_in_4 ? 8'hde : _GEN_1179; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1181 = 8'h9d == io_state_in_4 ? 8'h5e : _GEN_1180; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1182 = 8'h9e == io_state_in_4 ? 8'hb : _GEN_1181; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1183 = 8'h9f == io_state_in_4 ? 8'hdb : _GEN_1182; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1184 = 8'ha0 == io_state_in_4 ? 8'he0 : _GEN_1183; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1185 = 8'ha1 == io_state_in_4 ? 8'h32 : _GEN_1184; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1186 = 8'ha2 == io_state_in_4 ? 8'h3a : _GEN_1185; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1187 = 8'ha3 == io_state_in_4 ? 8'ha : _GEN_1186; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1188 = 8'ha4 == io_state_in_4 ? 8'h49 : _GEN_1187; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1189 = 8'ha5 == io_state_in_4 ? 8'h6 : _GEN_1188; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1190 = 8'ha6 == io_state_in_4 ? 8'h24 : _GEN_1189; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1191 = 8'ha7 == io_state_in_4 ? 8'h5c : _GEN_1190; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1192 = 8'ha8 == io_state_in_4 ? 8'hc2 : _GEN_1191; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1193 = 8'ha9 == io_state_in_4 ? 8'hd3 : _GEN_1192; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1194 = 8'haa == io_state_in_4 ? 8'hac : _GEN_1193; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1195 = 8'hab == io_state_in_4 ? 8'h62 : _GEN_1194; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1196 = 8'hac == io_state_in_4 ? 8'h91 : _GEN_1195; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1197 = 8'had == io_state_in_4 ? 8'h95 : _GEN_1196; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1198 = 8'hae == io_state_in_4 ? 8'he4 : _GEN_1197; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1199 = 8'haf == io_state_in_4 ? 8'h79 : _GEN_1198; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1200 = 8'hb0 == io_state_in_4 ? 8'he7 : _GEN_1199; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1201 = 8'hb1 == io_state_in_4 ? 8'hc8 : _GEN_1200; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1202 = 8'hb2 == io_state_in_4 ? 8'h37 : _GEN_1201; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1203 = 8'hb3 == io_state_in_4 ? 8'h6d : _GEN_1202; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1204 = 8'hb4 == io_state_in_4 ? 8'h8d : _GEN_1203; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1205 = 8'hb5 == io_state_in_4 ? 8'hd5 : _GEN_1204; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1206 = 8'hb6 == io_state_in_4 ? 8'h4e : _GEN_1205; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1207 = 8'hb7 == io_state_in_4 ? 8'ha9 : _GEN_1206; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1208 = 8'hb8 == io_state_in_4 ? 8'h6c : _GEN_1207; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1209 = 8'hb9 == io_state_in_4 ? 8'h56 : _GEN_1208; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1210 = 8'hba == io_state_in_4 ? 8'hf4 : _GEN_1209; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1211 = 8'hbb == io_state_in_4 ? 8'hea : _GEN_1210; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1212 = 8'hbc == io_state_in_4 ? 8'h65 : _GEN_1211; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1213 = 8'hbd == io_state_in_4 ? 8'h7a : _GEN_1212; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1214 = 8'hbe == io_state_in_4 ? 8'hae : _GEN_1213; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1215 = 8'hbf == io_state_in_4 ? 8'h8 : _GEN_1214; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1216 = 8'hc0 == io_state_in_4 ? 8'hba : _GEN_1215; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1217 = 8'hc1 == io_state_in_4 ? 8'h78 : _GEN_1216; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1218 = 8'hc2 == io_state_in_4 ? 8'h25 : _GEN_1217; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1219 = 8'hc3 == io_state_in_4 ? 8'h2e : _GEN_1218; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1220 = 8'hc4 == io_state_in_4 ? 8'h1c : _GEN_1219; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1221 = 8'hc5 == io_state_in_4 ? 8'ha6 : _GEN_1220; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1222 = 8'hc6 == io_state_in_4 ? 8'hb4 : _GEN_1221; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1223 = 8'hc7 == io_state_in_4 ? 8'hc6 : _GEN_1222; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1224 = 8'hc8 == io_state_in_4 ? 8'he8 : _GEN_1223; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1225 = 8'hc9 == io_state_in_4 ? 8'hdd : _GEN_1224; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1226 = 8'hca == io_state_in_4 ? 8'h74 : _GEN_1225; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1227 = 8'hcb == io_state_in_4 ? 8'h1f : _GEN_1226; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1228 = 8'hcc == io_state_in_4 ? 8'h4b : _GEN_1227; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1229 = 8'hcd == io_state_in_4 ? 8'hbd : _GEN_1228; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1230 = 8'hce == io_state_in_4 ? 8'h8b : _GEN_1229; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1231 = 8'hcf == io_state_in_4 ? 8'h8a : _GEN_1230; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1232 = 8'hd0 == io_state_in_4 ? 8'h70 : _GEN_1231; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1233 = 8'hd1 == io_state_in_4 ? 8'h3e : _GEN_1232; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1234 = 8'hd2 == io_state_in_4 ? 8'hb5 : _GEN_1233; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1235 = 8'hd3 == io_state_in_4 ? 8'h66 : _GEN_1234; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1236 = 8'hd4 == io_state_in_4 ? 8'h48 : _GEN_1235; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1237 = 8'hd5 == io_state_in_4 ? 8'h3 : _GEN_1236; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1238 = 8'hd6 == io_state_in_4 ? 8'hf6 : _GEN_1237; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1239 = 8'hd7 == io_state_in_4 ? 8'he : _GEN_1238; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1240 = 8'hd8 == io_state_in_4 ? 8'h61 : _GEN_1239; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1241 = 8'hd9 == io_state_in_4 ? 8'h35 : _GEN_1240; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1242 = 8'hda == io_state_in_4 ? 8'h57 : _GEN_1241; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1243 = 8'hdb == io_state_in_4 ? 8'hb9 : _GEN_1242; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1244 = 8'hdc == io_state_in_4 ? 8'h86 : _GEN_1243; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1245 = 8'hdd == io_state_in_4 ? 8'hc1 : _GEN_1244; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1246 = 8'hde == io_state_in_4 ? 8'h1d : _GEN_1245; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1247 = 8'hdf == io_state_in_4 ? 8'h9e : _GEN_1246; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1248 = 8'he0 == io_state_in_4 ? 8'he1 : _GEN_1247; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1249 = 8'he1 == io_state_in_4 ? 8'hf8 : _GEN_1248; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1250 = 8'he2 == io_state_in_4 ? 8'h98 : _GEN_1249; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1251 = 8'he3 == io_state_in_4 ? 8'h11 : _GEN_1250; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1252 = 8'he4 == io_state_in_4 ? 8'h69 : _GEN_1251; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1253 = 8'he5 == io_state_in_4 ? 8'hd9 : _GEN_1252; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1254 = 8'he6 == io_state_in_4 ? 8'h8e : _GEN_1253; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1255 = 8'he7 == io_state_in_4 ? 8'h94 : _GEN_1254; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1256 = 8'he8 == io_state_in_4 ? 8'h9b : _GEN_1255; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1257 = 8'he9 == io_state_in_4 ? 8'h1e : _GEN_1256; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1258 = 8'hea == io_state_in_4 ? 8'h87 : _GEN_1257; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1259 = 8'heb == io_state_in_4 ? 8'he9 : _GEN_1258; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1260 = 8'hec == io_state_in_4 ? 8'hce : _GEN_1259; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1261 = 8'hed == io_state_in_4 ? 8'h55 : _GEN_1260; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1262 = 8'hee == io_state_in_4 ? 8'h28 : _GEN_1261; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1263 = 8'hef == io_state_in_4 ? 8'hdf : _GEN_1262; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1264 = 8'hf0 == io_state_in_4 ? 8'h8c : _GEN_1263; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1265 = 8'hf1 == io_state_in_4 ? 8'ha1 : _GEN_1264; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1266 = 8'hf2 == io_state_in_4 ? 8'h89 : _GEN_1265; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1267 = 8'hf3 == io_state_in_4 ? 8'hd : _GEN_1266; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1268 = 8'hf4 == io_state_in_4 ? 8'hbf : _GEN_1267; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1269 = 8'hf5 == io_state_in_4 ? 8'he6 : _GEN_1268; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1270 = 8'hf6 == io_state_in_4 ? 8'h42 : _GEN_1269; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1271 = 8'hf7 == io_state_in_4 ? 8'h68 : _GEN_1270; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1272 = 8'hf8 == io_state_in_4 ? 8'h41 : _GEN_1271; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1273 = 8'hf9 == io_state_in_4 ? 8'h99 : _GEN_1272; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1274 = 8'hfa == io_state_in_4 ? 8'h2d : _GEN_1273; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1275 = 8'hfb == io_state_in_4 ? 8'hf : _GEN_1274; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1276 = 8'hfc == io_state_in_4 ? 8'hb0 : _GEN_1275; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1277 = 8'hfd == io_state_in_4 ? 8'h54 : _GEN_1276; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1278 = 8'hfe == io_state_in_4 ? 8'hbb : _GEN_1277; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1281 = 8'h1 == io_state_in_5 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1282 = 8'h2 == io_state_in_5 ? 8'h77 : _GEN_1281; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1283 = 8'h3 == io_state_in_5 ? 8'h7b : _GEN_1282; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1284 = 8'h4 == io_state_in_5 ? 8'hf2 : _GEN_1283; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1285 = 8'h5 == io_state_in_5 ? 8'h6b : _GEN_1284; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1286 = 8'h6 == io_state_in_5 ? 8'h6f : _GEN_1285; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1287 = 8'h7 == io_state_in_5 ? 8'hc5 : _GEN_1286; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1288 = 8'h8 == io_state_in_5 ? 8'h30 : _GEN_1287; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1289 = 8'h9 == io_state_in_5 ? 8'h1 : _GEN_1288; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1290 = 8'ha == io_state_in_5 ? 8'h67 : _GEN_1289; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1291 = 8'hb == io_state_in_5 ? 8'h2b : _GEN_1290; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1292 = 8'hc == io_state_in_5 ? 8'hfe : _GEN_1291; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1293 = 8'hd == io_state_in_5 ? 8'hd7 : _GEN_1292; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1294 = 8'he == io_state_in_5 ? 8'hab : _GEN_1293; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1295 = 8'hf == io_state_in_5 ? 8'h76 : _GEN_1294; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1296 = 8'h10 == io_state_in_5 ? 8'hca : _GEN_1295; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1297 = 8'h11 == io_state_in_5 ? 8'h82 : _GEN_1296; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1298 = 8'h12 == io_state_in_5 ? 8'hc9 : _GEN_1297; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1299 = 8'h13 == io_state_in_5 ? 8'h7d : _GEN_1298; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1300 = 8'h14 == io_state_in_5 ? 8'hfa : _GEN_1299; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1301 = 8'h15 == io_state_in_5 ? 8'h59 : _GEN_1300; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1302 = 8'h16 == io_state_in_5 ? 8'h47 : _GEN_1301; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1303 = 8'h17 == io_state_in_5 ? 8'hf0 : _GEN_1302; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1304 = 8'h18 == io_state_in_5 ? 8'had : _GEN_1303; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1305 = 8'h19 == io_state_in_5 ? 8'hd4 : _GEN_1304; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1306 = 8'h1a == io_state_in_5 ? 8'ha2 : _GEN_1305; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1307 = 8'h1b == io_state_in_5 ? 8'haf : _GEN_1306; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1308 = 8'h1c == io_state_in_5 ? 8'h9c : _GEN_1307; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1309 = 8'h1d == io_state_in_5 ? 8'ha4 : _GEN_1308; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1310 = 8'h1e == io_state_in_5 ? 8'h72 : _GEN_1309; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1311 = 8'h1f == io_state_in_5 ? 8'hc0 : _GEN_1310; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1312 = 8'h20 == io_state_in_5 ? 8'hb7 : _GEN_1311; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1313 = 8'h21 == io_state_in_5 ? 8'hfd : _GEN_1312; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1314 = 8'h22 == io_state_in_5 ? 8'h93 : _GEN_1313; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1315 = 8'h23 == io_state_in_5 ? 8'h26 : _GEN_1314; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1316 = 8'h24 == io_state_in_5 ? 8'h36 : _GEN_1315; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1317 = 8'h25 == io_state_in_5 ? 8'h3f : _GEN_1316; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1318 = 8'h26 == io_state_in_5 ? 8'hf7 : _GEN_1317; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1319 = 8'h27 == io_state_in_5 ? 8'hcc : _GEN_1318; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1320 = 8'h28 == io_state_in_5 ? 8'h34 : _GEN_1319; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1321 = 8'h29 == io_state_in_5 ? 8'ha5 : _GEN_1320; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1322 = 8'h2a == io_state_in_5 ? 8'he5 : _GEN_1321; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1323 = 8'h2b == io_state_in_5 ? 8'hf1 : _GEN_1322; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1324 = 8'h2c == io_state_in_5 ? 8'h71 : _GEN_1323; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1325 = 8'h2d == io_state_in_5 ? 8'hd8 : _GEN_1324; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1326 = 8'h2e == io_state_in_5 ? 8'h31 : _GEN_1325; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1327 = 8'h2f == io_state_in_5 ? 8'h15 : _GEN_1326; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1328 = 8'h30 == io_state_in_5 ? 8'h4 : _GEN_1327; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1329 = 8'h31 == io_state_in_5 ? 8'hc7 : _GEN_1328; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1330 = 8'h32 == io_state_in_5 ? 8'h23 : _GEN_1329; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1331 = 8'h33 == io_state_in_5 ? 8'hc3 : _GEN_1330; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1332 = 8'h34 == io_state_in_5 ? 8'h18 : _GEN_1331; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1333 = 8'h35 == io_state_in_5 ? 8'h96 : _GEN_1332; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1334 = 8'h36 == io_state_in_5 ? 8'h5 : _GEN_1333; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1335 = 8'h37 == io_state_in_5 ? 8'h9a : _GEN_1334; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1336 = 8'h38 == io_state_in_5 ? 8'h7 : _GEN_1335; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1337 = 8'h39 == io_state_in_5 ? 8'h12 : _GEN_1336; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1338 = 8'h3a == io_state_in_5 ? 8'h80 : _GEN_1337; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1339 = 8'h3b == io_state_in_5 ? 8'he2 : _GEN_1338; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1340 = 8'h3c == io_state_in_5 ? 8'heb : _GEN_1339; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1341 = 8'h3d == io_state_in_5 ? 8'h27 : _GEN_1340; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1342 = 8'h3e == io_state_in_5 ? 8'hb2 : _GEN_1341; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1343 = 8'h3f == io_state_in_5 ? 8'h75 : _GEN_1342; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1344 = 8'h40 == io_state_in_5 ? 8'h9 : _GEN_1343; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1345 = 8'h41 == io_state_in_5 ? 8'h83 : _GEN_1344; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1346 = 8'h42 == io_state_in_5 ? 8'h2c : _GEN_1345; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1347 = 8'h43 == io_state_in_5 ? 8'h1a : _GEN_1346; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1348 = 8'h44 == io_state_in_5 ? 8'h1b : _GEN_1347; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1349 = 8'h45 == io_state_in_5 ? 8'h6e : _GEN_1348; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1350 = 8'h46 == io_state_in_5 ? 8'h5a : _GEN_1349; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1351 = 8'h47 == io_state_in_5 ? 8'ha0 : _GEN_1350; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1352 = 8'h48 == io_state_in_5 ? 8'h52 : _GEN_1351; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1353 = 8'h49 == io_state_in_5 ? 8'h3b : _GEN_1352; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1354 = 8'h4a == io_state_in_5 ? 8'hd6 : _GEN_1353; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1355 = 8'h4b == io_state_in_5 ? 8'hb3 : _GEN_1354; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1356 = 8'h4c == io_state_in_5 ? 8'h29 : _GEN_1355; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1357 = 8'h4d == io_state_in_5 ? 8'he3 : _GEN_1356; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1358 = 8'h4e == io_state_in_5 ? 8'h2f : _GEN_1357; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1359 = 8'h4f == io_state_in_5 ? 8'h84 : _GEN_1358; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1360 = 8'h50 == io_state_in_5 ? 8'h53 : _GEN_1359; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1361 = 8'h51 == io_state_in_5 ? 8'hd1 : _GEN_1360; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1362 = 8'h52 == io_state_in_5 ? 8'h0 : _GEN_1361; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1363 = 8'h53 == io_state_in_5 ? 8'hed : _GEN_1362; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1364 = 8'h54 == io_state_in_5 ? 8'h20 : _GEN_1363; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1365 = 8'h55 == io_state_in_5 ? 8'hfc : _GEN_1364; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1366 = 8'h56 == io_state_in_5 ? 8'hb1 : _GEN_1365; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1367 = 8'h57 == io_state_in_5 ? 8'h5b : _GEN_1366; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1368 = 8'h58 == io_state_in_5 ? 8'h6a : _GEN_1367; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1369 = 8'h59 == io_state_in_5 ? 8'hcb : _GEN_1368; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1370 = 8'h5a == io_state_in_5 ? 8'hbe : _GEN_1369; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1371 = 8'h5b == io_state_in_5 ? 8'h39 : _GEN_1370; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1372 = 8'h5c == io_state_in_5 ? 8'h4a : _GEN_1371; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1373 = 8'h5d == io_state_in_5 ? 8'h4c : _GEN_1372; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1374 = 8'h5e == io_state_in_5 ? 8'h58 : _GEN_1373; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1375 = 8'h5f == io_state_in_5 ? 8'hcf : _GEN_1374; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1376 = 8'h60 == io_state_in_5 ? 8'hd0 : _GEN_1375; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1377 = 8'h61 == io_state_in_5 ? 8'hef : _GEN_1376; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1378 = 8'h62 == io_state_in_5 ? 8'haa : _GEN_1377; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1379 = 8'h63 == io_state_in_5 ? 8'hfb : _GEN_1378; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1380 = 8'h64 == io_state_in_5 ? 8'h43 : _GEN_1379; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1381 = 8'h65 == io_state_in_5 ? 8'h4d : _GEN_1380; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1382 = 8'h66 == io_state_in_5 ? 8'h33 : _GEN_1381; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1383 = 8'h67 == io_state_in_5 ? 8'h85 : _GEN_1382; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1384 = 8'h68 == io_state_in_5 ? 8'h45 : _GEN_1383; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1385 = 8'h69 == io_state_in_5 ? 8'hf9 : _GEN_1384; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1386 = 8'h6a == io_state_in_5 ? 8'h2 : _GEN_1385; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1387 = 8'h6b == io_state_in_5 ? 8'h7f : _GEN_1386; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1388 = 8'h6c == io_state_in_5 ? 8'h50 : _GEN_1387; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1389 = 8'h6d == io_state_in_5 ? 8'h3c : _GEN_1388; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1390 = 8'h6e == io_state_in_5 ? 8'h9f : _GEN_1389; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1391 = 8'h6f == io_state_in_5 ? 8'ha8 : _GEN_1390; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1392 = 8'h70 == io_state_in_5 ? 8'h51 : _GEN_1391; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1393 = 8'h71 == io_state_in_5 ? 8'ha3 : _GEN_1392; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1394 = 8'h72 == io_state_in_5 ? 8'h40 : _GEN_1393; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1395 = 8'h73 == io_state_in_5 ? 8'h8f : _GEN_1394; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1396 = 8'h74 == io_state_in_5 ? 8'h92 : _GEN_1395; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1397 = 8'h75 == io_state_in_5 ? 8'h9d : _GEN_1396; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1398 = 8'h76 == io_state_in_5 ? 8'h38 : _GEN_1397; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1399 = 8'h77 == io_state_in_5 ? 8'hf5 : _GEN_1398; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1400 = 8'h78 == io_state_in_5 ? 8'hbc : _GEN_1399; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1401 = 8'h79 == io_state_in_5 ? 8'hb6 : _GEN_1400; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1402 = 8'h7a == io_state_in_5 ? 8'hda : _GEN_1401; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1403 = 8'h7b == io_state_in_5 ? 8'h21 : _GEN_1402; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1404 = 8'h7c == io_state_in_5 ? 8'h10 : _GEN_1403; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1405 = 8'h7d == io_state_in_5 ? 8'hff : _GEN_1404; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1406 = 8'h7e == io_state_in_5 ? 8'hf3 : _GEN_1405; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1407 = 8'h7f == io_state_in_5 ? 8'hd2 : _GEN_1406; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1408 = 8'h80 == io_state_in_5 ? 8'hcd : _GEN_1407; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1409 = 8'h81 == io_state_in_5 ? 8'hc : _GEN_1408; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1410 = 8'h82 == io_state_in_5 ? 8'h13 : _GEN_1409; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1411 = 8'h83 == io_state_in_5 ? 8'hec : _GEN_1410; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1412 = 8'h84 == io_state_in_5 ? 8'h5f : _GEN_1411; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1413 = 8'h85 == io_state_in_5 ? 8'h97 : _GEN_1412; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1414 = 8'h86 == io_state_in_5 ? 8'h44 : _GEN_1413; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1415 = 8'h87 == io_state_in_5 ? 8'h17 : _GEN_1414; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1416 = 8'h88 == io_state_in_5 ? 8'hc4 : _GEN_1415; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1417 = 8'h89 == io_state_in_5 ? 8'ha7 : _GEN_1416; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1418 = 8'h8a == io_state_in_5 ? 8'h7e : _GEN_1417; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1419 = 8'h8b == io_state_in_5 ? 8'h3d : _GEN_1418; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1420 = 8'h8c == io_state_in_5 ? 8'h64 : _GEN_1419; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1421 = 8'h8d == io_state_in_5 ? 8'h5d : _GEN_1420; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1422 = 8'h8e == io_state_in_5 ? 8'h19 : _GEN_1421; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1423 = 8'h8f == io_state_in_5 ? 8'h73 : _GEN_1422; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1424 = 8'h90 == io_state_in_5 ? 8'h60 : _GEN_1423; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1425 = 8'h91 == io_state_in_5 ? 8'h81 : _GEN_1424; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1426 = 8'h92 == io_state_in_5 ? 8'h4f : _GEN_1425; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1427 = 8'h93 == io_state_in_5 ? 8'hdc : _GEN_1426; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1428 = 8'h94 == io_state_in_5 ? 8'h22 : _GEN_1427; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1429 = 8'h95 == io_state_in_5 ? 8'h2a : _GEN_1428; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1430 = 8'h96 == io_state_in_5 ? 8'h90 : _GEN_1429; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1431 = 8'h97 == io_state_in_5 ? 8'h88 : _GEN_1430; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1432 = 8'h98 == io_state_in_5 ? 8'h46 : _GEN_1431; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1433 = 8'h99 == io_state_in_5 ? 8'hee : _GEN_1432; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1434 = 8'h9a == io_state_in_5 ? 8'hb8 : _GEN_1433; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1435 = 8'h9b == io_state_in_5 ? 8'h14 : _GEN_1434; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1436 = 8'h9c == io_state_in_5 ? 8'hde : _GEN_1435; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1437 = 8'h9d == io_state_in_5 ? 8'h5e : _GEN_1436; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1438 = 8'h9e == io_state_in_5 ? 8'hb : _GEN_1437; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1439 = 8'h9f == io_state_in_5 ? 8'hdb : _GEN_1438; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1440 = 8'ha0 == io_state_in_5 ? 8'he0 : _GEN_1439; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1441 = 8'ha1 == io_state_in_5 ? 8'h32 : _GEN_1440; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1442 = 8'ha2 == io_state_in_5 ? 8'h3a : _GEN_1441; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1443 = 8'ha3 == io_state_in_5 ? 8'ha : _GEN_1442; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1444 = 8'ha4 == io_state_in_5 ? 8'h49 : _GEN_1443; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1445 = 8'ha5 == io_state_in_5 ? 8'h6 : _GEN_1444; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1446 = 8'ha6 == io_state_in_5 ? 8'h24 : _GEN_1445; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1447 = 8'ha7 == io_state_in_5 ? 8'h5c : _GEN_1446; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1448 = 8'ha8 == io_state_in_5 ? 8'hc2 : _GEN_1447; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1449 = 8'ha9 == io_state_in_5 ? 8'hd3 : _GEN_1448; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1450 = 8'haa == io_state_in_5 ? 8'hac : _GEN_1449; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1451 = 8'hab == io_state_in_5 ? 8'h62 : _GEN_1450; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1452 = 8'hac == io_state_in_5 ? 8'h91 : _GEN_1451; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1453 = 8'had == io_state_in_5 ? 8'h95 : _GEN_1452; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1454 = 8'hae == io_state_in_5 ? 8'he4 : _GEN_1453; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1455 = 8'haf == io_state_in_5 ? 8'h79 : _GEN_1454; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1456 = 8'hb0 == io_state_in_5 ? 8'he7 : _GEN_1455; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1457 = 8'hb1 == io_state_in_5 ? 8'hc8 : _GEN_1456; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1458 = 8'hb2 == io_state_in_5 ? 8'h37 : _GEN_1457; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1459 = 8'hb3 == io_state_in_5 ? 8'h6d : _GEN_1458; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1460 = 8'hb4 == io_state_in_5 ? 8'h8d : _GEN_1459; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1461 = 8'hb5 == io_state_in_5 ? 8'hd5 : _GEN_1460; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1462 = 8'hb6 == io_state_in_5 ? 8'h4e : _GEN_1461; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1463 = 8'hb7 == io_state_in_5 ? 8'ha9 : _GEN_1462; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1464 = 8'hb8 == io_state_in_5 ? 8'h6c : _GEN_1463; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1465 = 8'hb9 == io_state_in_5 ? 8'h56 : _GEN_1464; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1466 = 8'hba == io_state_in_5 ? 8'hf4 : _GEN_1465; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1467 = 8'hbb == io_state_in_5 ? 8'hea : _GEN_1466; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1468 = 8'hbc == io_state_in_5 ? 8'h65 : _GEN_1467; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1469 = 8'hbd == io_state_in_5 ? 8'h7a : _GEN_1468; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1470 = 8'hbe == io_state_in_5 ? 8'hae : _GEN_1469; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1471 = 8'hbf == io_state_in_5 ? 8'h8 : _GEN_1470; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1472 = 8'hc0 == io_state_in_5 ? 8'hba : _GEN_1471; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1473 = 8'hc1 == io_state_in_5 ? 8'h78 : _GEN_1472; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1474 = 8'hc2 == io_state_in_5 ? 8'h25 : _GEN_1473; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1475 = 8'hc3 == io_state_in_5 ? 8'h2e : _GEN_1474; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1476 = 8'hc4 == io_state_in_5 ? 8'h1c : _GEN_1475; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1477 = 8'hc5 == io_state_in_5 ? 8'ha6 : _GEN_1476; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1478 = 8'hc6 == io_state_in_5 ? 8'hb4 : _GEN_1477; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1479 = 8'hc7 == io_state_in_5 ? 8'hc6 : _GEN_1478; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1480 = 8'hc8 == io_state_in_5 ? 8'he8 : _GEN_1479; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1481 = 8'hc9 == io_state_in_5 ? 8'hdd : _GEN_1480; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1482 = 8'hca == io_state_in_5 ? 8'h74 : _GEN_1481; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1483 = 8'hcb == io_state_in_5 ? 8'h1f : _GEN_1482; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1484 = 8'hcc == io_state_in_5 ? 8'h4b : _GEN_1483; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1485 = 8'hcd == io_state_in_5 ? 8'hbd : _GEN_1484; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1486 = 8'hce == io_state_in_5 ? 8'h8b : _GEN_1485; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1487 = 8'hcf == io_state_in_5 ? 8'h8a : _GEN_1486; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1488 = 8'hd0 == io_state_in_5 ? 8'h70 : _GEN_1487; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1489 = 8'hd1 == io_state_in_5 ? 8'h3e : _GEN_1488; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1490 = 8'hd2 == io_state_in_5 ? 8'hb5 : _GEN_1489; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1491 = 8'hd3 == io_state_in_5 ? 8'h66 : _GEN_1490; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1492 = 8'hd4 == io_state_in_5 ? 8'h48 : _GEN_1491; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1493 = 8'hd5 == io_state_in_5 ? 8'h3 : _GEN_1492; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1494 = 8'hd6 == io_state_in_5 ? 8'hf6 : _GEN_1493; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1495 = 8'hd7 == io_state_in_5 ? 8'he : _GEN_1494; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1496 = 8'hd8 == io_state_in_5 ? 8'h61 : _GEN_1495; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1497 = 8'hd9 == io_state_in_5 ? 8'h35 : _GEN_1496; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1498 = 8'hda == io_state_in_5 ? 8'h57 : _GEN_1497; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1499 = 8'hdb == io_state_in_5 ? 8'hb9 : _GEN_1498; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1500 = 8'hdc == io_state_in_5 ? 8'h86 : _GEN_1499; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1501 = 8'hdd == io_state_in_5 ? 8'hc1 : _GEN_1500; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1502 = 8'hde == io_state_in_5 ? 8'h1d : _GEN_1501; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1503 = 8'hdf == io_state_in_5 ? 8'h9e : _GEN_1502; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1504 = 8'he0 == io_state_in_5 ? 8'he1 : _GEN_1503; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1505 = 8'he1 == io_state_in_5 ? 8'hf8 : _GEN_1504; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1506 = 8'he2 == io_state_in_5 ? 8'h98 : _GEN_1505; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1507 = 8'he3 == io_state_in_5 ? 8'h11 : _GEN_1506; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1508 = 8'he4 == io_state_in_5 ? 8'h69 : _GEN_1507; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1509 = 8'he5 == io_state_in_5 ? 8'hd9 : _GEN_1508; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1510 = 8'he6 == io_state_in_5 ? 8'h8e : _GEN_1509; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1511 = 8'he7 == io_state_in_5 ? 8'h94 : _GEN_1510; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1512 = 8'he8 == io_state_in_5 ? 8'h9b : _GEN_1511; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1513 = 8'he9 == io_state_in_5 ? 8'h1e : _GEN_1512; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1514 = 8'hea == io_state_in_5 ? 8'h87 : _GEN_1513; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1515 = 8'heb == io_state_in_5 ? 8'he9 : _GEN_1514; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1516 = 8'hec == io_state_in_5 ? 8'hce : _GEN_1515; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1517 = 8'hed == io_state_in_5 ? 8'h55 : _GEN_1516; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1518 = 8'hee == io_state_in_5 ? 8'h28 : _GEN_1517; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1519 = 8'hef == io_state_in_5 ? 8'hdf : _GEN_1518; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1520 = 8'hf0 == io_state_in_5 ? 8'h8c : _GEN_1519; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1521 = 8'hf1 == io_state_in_5 ? 8'ha1 : _GEN_1520; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1522 = 8'hf2 == io_state_in_5 ? 8'h89 : _GEN_1521; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1523 = 8'hf3 == io_state_in_5 ? 8'hd : _GEN_1522; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1524 = 8'hf4 == io_state_in_5 ? 8'hbf : _GEN_1523; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1525 = 8'hf5 == io_state_in_5 ? 8'he6 : _GEN_1524; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1526 = 8'hf6 == io_state_in_5 ? 8'h42 : _GEN_1525; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1527 = 8'hf7 == io_state_in_5 ? 8'h68 : _GEN_1526; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1528 = 8'hf8 == io_state_in_5 ? 8'h41 : _GEN_1527; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1529 = 8'hf9 == io_state_in_5 ? 8'h99 : _GEN_1528; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1530 = 8'hfa == io_state_in_5 ? 8'h2d : _GEN_1529; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1531 = 8'hfb == io_state_in_5 ? 8'hf : _GEN_1530; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1532 = 8'hfc == io_state_in_5 ? 8'hb0 : _GEN_1531; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1533 = 8'hfd == io_state_in_5 ? 8'h54 : _GEN_1532; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1534 = 8'hfe == io_state_in_5 ? 8'hbb : _GEN_1533; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1537 = 8'h1 == io_state_in_6 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1538 = 8'h2 == io_state_in_6 ? 8'h77 : _GEN_1537; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1539 = 8'h3 == io_state_in_6 ? 8'h7b : _GEN_1538; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1540 = 8'h4 == io_state_in_6 ? 8'hf2 : _GEN_1539; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1541 = 8'h5 == io_state_in_6 ? 8'h6b : _GEN_1540; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1542 = 8'h6 == io_state_in_6 ? 8'h6f : _GEN_1541; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1543 = 8'h7 == io_state_in_6 ? 8'hc5 : _GEN_1542; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1544 = 8'h8 == io_state_in_6 ? 8'h30 : _GEN_1543; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1545 = 8'h9 == io_state_in_6 ? 8'h1 : _GEN_1544; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1546 = 8'ha == io_state_in_6 ? 8'h67 : _GEN_1545; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1547 = 8'hb == io_state_in_6 ? 8'h2b : _GEN_1546; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1548 = 8'hc == io_state_in_6 ? 8'hfe : _GEN_1547; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1549 = 8'hd == io_state_in_6 ? 8'hd7 : _GEN_1548; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1550 = 8'he == io_state_in_6 ? 8'hab : _GEN_1549; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1551 = 8'hf == io_state_in_6 ? 8'h76 : _GEN_1550; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1552 = 8'h10 == io_state_in_6 ? 8'hca : _GEN_1551; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1553 = 8'h11 == io_state_in_6 ? 8'h82 : _GEN_1552; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1554 = 8'h12 == io_state_in_6 ? 8'hc9 : _GEN_1553; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1555 = 8'h13 == io_state_in_6 ? 8'h7d : _GEN_1554; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1556 = 8'h14 == io_state_in_6 ? 8'hfa : _GEN_1555; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1557 = 8'h15 == io_state_in_6 ? 8'h59 : _GEN_1556; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1558 = 8'h16 == io_state_in_6 ? 8'h47 : _GEN_1557; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1559 = 8'h17 == io_state_in_6 ? 8'hf0 : _GEN_1558; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1560 = 8'h18 == io_state_in_6 ? 8'had : _GEN_1559; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1561 = 8'h19 == io_state_in_6 ? 8'hd4 : _GEN_1560; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1562 = 8'h1a == io_state_in_6 ? 8'ha2 : _GEN_1561; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1563 = 8'h1b == io_state_in_6 ? 8'haf : _GEN_1562; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1564 = 8'h1c == io_state_in_6 ? 8'h9c : _GEN_1563; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1565 = 8'h1d == io_state_in_6 ? 8'ha4 : _GEN_1564; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1566 = 8'h1e == io_state_in_6 ? 8'h72 : _GEN_1565; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1567 = 8'h1f == io_state_in_6 ? 8'hc0 : _GEN_1566; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1568 = 8'h20 == io_state_in_6 ? 8'hb7 : _GEN_1567; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1569 = 8'h21 == io_state_in_6 ? 8'hfd : _GEN_1568; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1570 = 8'h22 == io_state_in_6 ? 8'h93 : _GEN_1569; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1571 = 8'h23 == io_state_in_6 ? 8'h26 : _GEN_1570; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1572 = 8'h24 == io_state_in_6 ? 8'h36 : _GEN_1571; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1573 = 8'h25 == io_state_in_6 ? 8'h3f : _GEN_1572; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1574 = 8'h26 == io_state_in_6 ? 8'hf7 : _GEN_1573; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1575 = 8'h27 == io_state_in_6 ? 8'hcc : _GEN_1574; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1576 = 8'h28 == io_state_in_6 ? 8'h34 : _GEN_1575; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1577 = 8'h29 == io_state_in_6 ? 8'ha5 : _GEN_1576; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1578 = 8'h2a == io_state_in_6 ? 8'he5 : _GEN_1577; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1579 = 8'h2b == io_state_in_6 ? 8'hf1 : _GEN_1578; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1580 = 8'h2c == io_state_in_6 ? 8'h71 : _GEN_1579; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1581 = 8'h2d == io_state_in_6 ? 8'hd8 : _GEN_1580; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1582 = 8'h2e == io_state_in_6 ? 8'h31 : _GEN_1581; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1583 = 8'h2f == io_state_in_6 ? 8'h15 : _GEN_1582; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1584 = 8'h30 == io_state_in_6 ? 8'h4 : _GEN_1583; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1585 = 8'h31 == io_state_in_6 ? 8'hc7 : _GEN_1584; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1586 = 8'h32 == io_state_in_6 ? 8'h23 : _GEN_1585; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1587 = 8'h33 == io_state_in_6 ? 8'hc3 : _GEN_1586; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1588 = 8'h34 == io_state_in_6 ? 8'h18 : _GEN_1587; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1589 = 8'h35 == io_state_in_6 ? 8'h96 : _GEN_1588; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1590 = 8'h36 == io_state_in_6 ? 8'h5 : _GEN_1589; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1591 = 8'h37 == io_state_in_6 ? 8'h9a : _GEN_1590; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1592 = 8'h38 == io_state_in_6 ? 8'h7 : _GEN_1591; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1593 = 8'h39 == io_state_in_6 ? 8'h12 : _GEN_1592; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1594 = 8'h3a == io_state_in_6 ? 8'h80 : _GEN_1593; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1595 = 8'h3b == io_state_in_6 ? 8'he2 : _GEN_1594; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1596 = 8'h3c == io_state_in_6 ? 8'heb : _GEN_1595; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1597 = 8'h3d == io_state_in_6 ? 8'h27 : _GEN_1596; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1598 = 8'h3e == io_state_in_6 ? 8'hb2 : _GEN_1597; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1599 = 8'h3f == io_state_in_6 ? 8'h75 : _GEN_1598; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1600 = 8'h40 == io_state_in_6 ? 8'h9 : _GEN_1599; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1601 = 8'h41 == io_state_in_6 ? 8'h83 : _GEN_1600; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1602 = 8'h42 == io_state_in_6 ? 8'h2c : _GEN_1601; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1603 = 8'h43 == io_state_in_6 ? 8'h1a : _GEN_1602; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1604 = 8'h44 == io_state_in_6 ? 8'h1b : _GEN_1603; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1605 = 8'h45 == io_state_in_6 ? 8'h6e : _GEN_1604; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1606 = 8'h46 == io_state_in_6 ? 8'h5a : _GEN_1605; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1607 = 8'h47 == io_state_in_6 ? 8'ha0 : _GEN_1606; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1608 = 8'h48 == io_state_in_6 ? 8'h52 : _GEN_1607; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1609 = 8'h49 == io_state_in_6 ? 8'h3b : _GEN_1608; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1610 = 8'h4a == io_state_in_6 ? 8'hd6 : _GEN_1609; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1611 = 8'h4b == io_state_in_6 ? 8'hb3 : _GEN_1610; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1612 = 8'h4c == io_state_in_6 ? 8'h29 : _GEN_1611; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1613 = 8'h4d == io_state_in_6 ? 8'he3 : _GEN_1612; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1614 = 8'h4e == io_state_in_6 ? 8'h2f : _GEN_1613; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1615 = 8'h4f == io_state_in_6 ? 8'h84 : _GEN_1614; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1616 = 8'h50 == io_state_in_6 ? 8'h53 : _GEN_1615; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1617 = 8'h51 == io_state_in_6 ? 8'hd1 : _GEN_1616; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1618 = 8'h52 == io_state_in_6 ? 8'h0 : _GEN_1617; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1619 = 8'h53 == io_state_in_6 ? 8'hed : _GEN_1618; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1620 = 8'h54 == io_state_in_6 ? 8'h20 : _GEN_1619; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1621 = 8'h55 == io_state_in_6 ? 8'hfc : _GEN_1620; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1622 = 8'h56 == io_state_in_6 ? 8'hb1 : _GEN_1621; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1623 = 8'h57 == io_state_in_6 ? 8'h5b : _GEN_1622; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1624 = 8'h58 == io_state_in_6 ? 8'h6a : _GEN_1623; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1625 = 8'h59 == io_state_in_6 ? 8'hcb : _GEN_1624; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1626 = 8'h5a == io_state_in_6 ? 8'hbe : _GEN_1625; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1627 = 8'h5b == io_state_in_6 ? 8'h39 : _GEN_1626; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1628 = 8'h5c == io_state_in_6 ? 8'h4a : _GEN_1627; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1629 = 8'h5d == io_state_in_6 ? 8'h4c : _GEN_1628; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1630 = 8'h5e == io_state_in_6 ? 8'h58 : _GEN_1629; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1631 = 8'h5f == io_state_in_6 ? 8'hcf : _GEN_1630; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1632 = 8'h60 == io_state_in_6 ? 8'hd0 : _GEN_1631; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1633 = 8'h61 == io_state_in_6 ? 8'hef : _GEN_1632; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1634 = 8'h62 == io_state_in_6 ? 8'haa : _GEN_1633; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1635 = 8'h63 == io_state_in_6 ? 8'hfb : _GEN_1634; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1636 = 8'h64 == io_state_in_6 ? 8'h43 : _GEN_1635; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1637 = 8'h65 == io_state_in_6 ? 8'h4d : _GEN_1636; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1638 = 8'h66 == io_state_in_6 ? 8'h33 : _GEN_1637; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1639 = 8'h67 == io_state_in_6 ? 8'h85 : _GEN_1638; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1640 = 8'h68 == io_state_in_6 ? 8'h45 : _GEN_1639; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1641 = 8'h69 == io_state_in_6 ? 8'hf9 : _GEN_1640; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1642 = 8'h6a == io_state_in_6 ? 8'h2 : _GEN_1641; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1643 = 8'h6b == io_state_in_6 ? 8'h7f : _GEN_1642; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1644 = 8'h6c == io_state_in_6 ? 8'h50 : _GEN_1643; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1645 = 8'h6d == io_state_in_6 ? 8'h3c : _GEN_1644; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1646 = 8'h6e == io_state_in_6 ? 8'h9f : _GEN_1645; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1647 = 8'h6f == io_state_in_6 ? 8'ha8 : _GEN_1646; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1648 = 8'h70 == io_state_in_6 ? 8'h51 : _GEN_1647; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1649 = 8'h71 == io_state_in_6 ? 8'ha3 : _GEN_1648; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1650 = 8'h72 == io_state_in_6 ? 8'h40 : _GEN_1649; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1651 = 8'h73 == io_state_in_6 ? 8'h8f : _GEN_1650; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1652 = 8'h74 == io_state_in_6 ? 8'h92 : _GEN_1651; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1653 = 8'h75 == io_state_in_6 ? 8'h9d : _GEN_1652; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1654 = 8'h76 == io_state_in_6 ? 8'h38 : _GEN_1653; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1655 = 8'h77 == io_state_in_6 ? 8'hf5 : _GEN_1654; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1656 = 8'h78 == io_state_in_6 ? 8'hbc : _GEN_1655; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1657 = 8'h79 == io_state_in_6 ? 8'hb6 : _GEN_1656; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1658 = 8'h7a == io_state_in_6 ? 8'hda : _GEN_1657; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1659 = 8'h7b == io_state_in_6 ? 8'h21 : _GEN_1658; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1660 = 8'h7c == io_state_in_6 ? 8'h10 : _GEN_1659; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1661 = 8'h7d == io_state_in_6 ? 8'hff : _GEN_1660; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1662 = 8'h7e == io_state_in_6 ? 8'hf3 : _GEN_1661; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1663 = 8'h7f == io_state_in_6 ? 8'hd2 : _GEN_1662; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1664 = 8'h80 == io_state_in_6 ? 8'hcd : _GEN_1663; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1665 = 8'h81 == io_state_in_6 ? 8'hc : _GEN_1664; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1666 = 8'h82 == io_state_in_6 ? 8'h13 : _GEN_1665; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1667 = 8'h83 == io_state_in_6 ? 8'hec : _GEN_1666; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1668 = 8'h84 == io_state_in_6 ? 8'h5f : _GEN_1667; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1669 = 8'h85 == io_state_in_6 ? 8'h97 : _GEN_1668; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1670 = 8'h86 == io_state_in_6 ? 8'h44 : _GEN_1669; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1671 = 8'h87 == io_state_in_6 ? 8'h17 : _GEN_1670; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1672 = 8'h88 == io_state_in_6 ? 8'hc4 : _GEN_1671; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1673 = 8'h89 == io_state_in_6 ? 8'ha7 : _GEN_1672; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1674 = 8'h8a == io_state_in_6 ? 8'h7e : _GEN_1673; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1675 = 8'h8b == io_state_in_6 ? 8'h3d : _GEN_1674; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1676 = 8'h8c == io_state_in_6 ? 8'h64 : _GEN_1675; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1677 = 8'h8d == io_state_in_6 ? 8'h5d : _GEN_1676; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1678 = 8'h8e == io_state_in_6 ? 8'h19 : _GEN_1677; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1679 = 8'h8f == io_state_in_6 ? 8'h73 : _GEN_1678; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1680 = 8'h90 == io_state_in_6 ? 8'h60 : _GEN_1679; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1681 = 8'h91 == io_state_in_6 ? 8'h81 : _GEN_1680; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1682 = 8'h92 == io_state_in_6 ? 8'h4f : _GEN_1681; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1683 = 8'h93 == io_state_in_6 ? 8'hdc : _GEN_1682; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1684 = 8'h94 == io_state_in_6 ? 8'h22 : _GEN_1683; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1685 = 8'h95 == io_state_in_6 ? 8'h2a : _GEN_1684; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1686 = 8'h96 == io_state_in_6 ? 8'h90 : _GEN_1685; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1687 = 8'h97 == io_state_in_6 ? 8'h88 : _GEN_1686; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1688 = 8'h98 == io_state_in_6 ? 8'h46 : _GEN_1687; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1689 = 8'h99 == io_state_in_6 ? 8'hee : _GEN_1688; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1690 = 8'h9a == io_state_in_6 ? 8'hb8 : _GEN_1689; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1691 = 8'h9b == io_state_in_6 ? 8'h14 : _GEN_1690; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1692 = 8'h9c == io_state_in_6 ? 8'hde : _GEN_1691; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1693 = 8'h9d == io_state_in_6 ? 8'h5e : _GEN_1692; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1694 = 8'h9e == io_state_in_6 ? 8'hb : _GEN_1693; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1695 = 8'h9f == io_state_in_6 ? 8'hdb : _GEN_1694; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1696 = 8'ha0 == io_state_in_6 ? 8'he0 : _GEN_1695; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1697 = 8'ha1 == io_state_in_6 ? 8'h32 : _GEN_1696; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1698 = 8'ha2 == io_state_in_6 ? 8'h3a : _GEN_1697; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1699 = 8'ha3 == io_state_in_6 ? 8'ha : _GEN_1698; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1700 = 8'ha4 == io_state_in_6 ? 8'h49 : _GEN_1699; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1701 = 8'ha5 == io_state_in_6 ? 8'h6 : _GEN_1700; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1702 = 8'ha6 == io_state_in_6 ? 8'h24 : _GEN_1701; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1703 = 8'ha7 == io_state_in_6 ? 8'h5c : _GEN_1702; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1704 = 8'ha8 == io_state_in_6 ? 8'hc2 : _GEN_1703; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1705 = 8'ha9 == io_state_in_6 ? 8'hd3 : _GEN_1704; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1706 = 8'haa == io_state_in_6 ? 8'hac : _GEN_1705; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1707 = 8'hab == io_state_in_6 ? 8'h62 : _GEN_1706; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1708 = 8'hac == io_state_in_6 ? 8'h91 : _GEN_1707; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1709 = 8'had == io_state_in_6 ? 8'h95 : _GEN_1708; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1710 = 8'hae == io_state_in_6 ? 8'he4 : _GEN_1709; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1711 = 8'haf == io_state_in_6 ? 8'h79 : _GEN_1710; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1712 = 8'hb0 == io_state_in_6 ? 8'he7 : _GEN_1711; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1713 = 8'hb1 == io_state_in_6 ? 8'hc8 : _GEN_1712; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1714 = 8'hb2 == io_state_in_6 ? 8'h37 : _GEN_1713; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1715 = 8'hb3 == io_state_in_6 ? 8'h6d : _GEN_1714; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1716 = 8'hb4 == io_state_in_6 ? 8'h8d : _GEN_1715; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1717 = 8'hb5 == io_state_in_6 ? 8'hd5 : _GEN_1716; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1718 = 8'hb6 == io_state_in_6 ? 8'h4e : _GEN_1717; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1719 = 8'hb7 == io_state_in_6 ? 8'ha9 : _GEN_1718; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1720 = 8'hb8 == io_state_in_6 ? 8'h6c : _GEN_1719; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1721 = 8'hb9 == io_state_in_6 ? 8'h56 : _GEN_1720; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1722 = 8'hba == io_state_in_6 ? 8'hf4 : _GEN_1721; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1723 = 8'hbb == io_state_in_6 ? 8'hea : _GEN_1722; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1724 = 8'hbc == io_state_in_6 ? 8'h65 : _GEN_1723; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1725 = 8'hbd == io_state_in_6 ? 8'h7a : _GEN_1724; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1726 = 8'hbe == io_state_in_6 ? 8'hae : _GEN_1725; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1727 = 8'hbf == io_state_in_6 ? 8'h8 : _GEN_1726; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1728 = 8'hc0 == io_state_in_6 ? 8'hba : _GEN_1727; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1729 = 8'hc1 == io_state_in_6 ? 8'h78 : _GEN_1728; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1730 = 8'hc2 == io_state_in_6 ? 8'h25 : _GEN_1729; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1731 = 8'hc3 == io_state_in_6 ? 8'h2e : _GEN_1730; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1732 = 8'hc4 == io_state_in_6 ? 8'h1c : _GEN_1731; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1733 = 8'hc5 == io_state_in_6 ? 8'ha6 : _GEN_1732; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1734 = 8'hc6 == io_state_in_6 ? 8'hb4 : _GEN_1733; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1735 = 8'hc7 == io_state_in_6 ? 8'hc6 : _GEN_1734; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1736 = 8'hc8 == io_state_in_6 ? 8'he8 : _GEN_1735; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1737 = 8'hc9 == io_state_in_6 ? 8'hdd : _GEN_1736; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1738 = 8'hca == io_state_in_6 ? 8'h74 : _GEN_1737; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1739 = 8'hcb == io_state_in_6 ? 8'h1f : _GEN_1738; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1740 = 8'hcc == io_state_in_6 ? 8'h4b : _GEN_1739; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1741 = 8'hcd == io_state_in_6 ? 8'hbd : _GEN_1740; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1742 = 8'hce == io_state_in_6 ? 8'h8b : _GEN_1741; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1743 = 8'hcf == io_state_in_6 ? 8'h8a : _GEN_1742; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1744 = 8'hd0 == io_state_in_6 ? 8'h70 : _GEN_1743; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1745 = 8'hd1 == io_state_in_6 ? 8'h3e : _GEN_1744; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1746 = 8'hd2 == io_state_in_6 ? 8'hb5 : _GEN_1745; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1747 = 8'hd3 == io_state_in_6 ? 8'h66 : _GEN_1746; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1748 = 8'hd4 == io_state_in_6 ? 8'h48 : _GEN_1747; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1749 = 8'hd5 == io_state_in_6 ? 8'h3 : _GEN_1748; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1750 = 8'hd6 == io_state_in_6 ? 8'hf6 : _GEN_1749; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1751 = 8'hd7 == io_state_in_6 ? 8'he : _GEN_1750; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1752 = 8'hd8 == io_state_in_6 ? 8'h61 : _GEN_1751; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1753 = 8'hd9 == io_state_in_6 ? 8'h35 : _GEN_1752; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1754 = 8'hda == io_state_in_6 ? 8'h57 : _GEN_1753; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1755 = 8'hdb == io_state_in_6 ? 8'hb9 : _GEN_1754; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1756 = 8'hdc == io_state_in_6 ? 8'h86 : _GEN_1755; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1757 = 8'hdd == io_state_in_6 ? 8'hc1 : _GEN_1756; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1758 = 8'hde == io_state_in_6 ? 8'h1d : _GEN_1757; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1759 = 8'hdf == io_state_in_6 ? 8'h9e : _GEN_1758; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1760 = 8'he0 == io_state_in_6 ? 8'he1 : _GEN_1759; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1761 = 8'he1 == io_state_in_6 ? 8'hf8 : _GEN_1760; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1762 = 8'he2 == io_state_in_6 ? 8'h98 : _GEN_1761; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1763 = 8'he3 == io_state_in_6 ? 8'h11 : _GEN_1762; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1764 = 8'he4 == io_state_in_6 ? 8'h69 : _GEN_1763; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1765 = 8'he5 == io_state_in_6 ? 8'hd9 : _GEN_1764; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1766 = 8'he6 == io_state_in_6 ? 8'h8e : _GEN_1765; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1767 = 8'he7 == io_state_in_6 ? 8'h94 : _GEN_1766; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1768 = 8'he8 == io_state_in_6 ? 8'h9b : _GEN_1767; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1769 = 8'he9 == io_state_in_6 ? 8'h1e : _GEN_1768; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1770 = 8'hea == io_state_in_6 ? 8'h87 : _GEN_1769; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1771 = 8'heb == io_state_in_6 ? 8'he9 : _GEN_1770; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1772 = 8'hec == io_state_in_6 ? 8'hce : _GEN_1771; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1773 = 8'hed == io_state_in_6 ? 8'h55 : _GEN_1772; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1774 = 8'hee == io_state_in_6 ? 8'h28 : _GEN_1773; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1775 = 8'hef == io_state_in_6 ? 8'hdf : _GEN_1774; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1776 = 8'hf0 == io_state_in_6 ? 8'h8c : _GEN_1775; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1777 = 8'hf1 == io_state_in_6 ? 8'ha1 : _GEN_1776; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1778 = 8'hf2 == io_state_in_6 ? 8'h89 : _GEN_1777; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1779 = 8'hf3 == io_state_in_6 ? 8'hd : _GEN_1778; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1780 = 8'hf4 == io_state_in_6 ? 8'hbf : _GEN_1779; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1781 = 8'hf5 == io_state_in_6 ? 8'he6 : _GEN_1780; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1782 = 8'hf6 == io_state_in_6 ? 8'h42 : _GEN_1781; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1783 = 8'hf7 == io_state_in_6 ? 8'h68 : _GEN_1782; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1784 = 8'hf8 == io_state_in_6 ? 8'h41 : _GEN_1783; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1785 = 8'hf9 == io_state_in_6 ? 8'h99 : _GEN_1784; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1786 = 8'hfa == io_state_in_6 ? 8'h2d : _GEN_1785; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1787 = 8'hfb == io_state_in_6 ? 8'hf : _GEN_1786; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1788 = 8'hfc == io_state_in_6 ? 8'hb0 : _GEN_1787; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1789 = 8'hfd == io_state_in_6 ? 8'h54 : _GEN_1788; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1790 = 8'hfe == io_state_in_6 ? 8'hbb : _GEN_1789; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1793 = 8'h1 == io_state_in_7 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1794 = 8'h2 == io_state_in_7 ? 8'h77 : _GEN_1793; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1795 = 8'h3 == io_state_in_7 ? 8'h7b : _GEN_1794; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1796 = 8'h4 == io_state_in_7 ? 8'hf2 : _GEN_1795; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1797 = 8'h5 == io_state_in_7 ? 8'h6b : _GEN_1796; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1798 = 8'h6 == io_state_in_7 ? 8'h6f : _GEN_1797; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1799 = 8'h7 == io_state_in_7 ? 8'hc5 : _GEN_1798; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1800 = 8'h8 == io_state_in_7 ? 8'h30 : _GEN_1799; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1801 = 8'h9 == io_state_in_7 ? 8'h1 : _GEN_1800; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1802 = 8'ha == io_state_in_7 ? 8'h67 : _GEN_1801; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1803 = 8'hb == io_state_in_7 ? 8'h2b : _GEN_1802; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1804 = 8'hc == io_state_in_7 ? 8'hfe : _GEN_1803; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1805 = 8'hd == io_state_in_7 ? 8'hd7 : _GEN_1804; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1806 = 8'he == io_state_in_7 ? 8'hab : _GEN_1805; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1807 = 8'hf == io_state_in_7 ? 8'h76 : _GEN_1806; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1808 = 8'h10 == io_state_in_7 ? 8'hca : _GEN_1807; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1809 = 8'h11 == io_state_in_7 ? 8'h82 : _GEN_1808; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1810 = 8'h12 == io_state_in_7 ? 8'hc9 : _GEN_1809; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1811 = 8'h13 == io_state_in_7 ? 8'h7d : _GEN_1810; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1812 = 8'h14 == io_state_in_7 ? 8'hfa : _GEN_1811; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1813 = 8'h15 == io_state_in_7 ? 8'h59 : _GEN_1812; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1814 = 8'h16 == io_state_in_7 ? 8'h47 : _GEN_1813; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1815 = 8'h17 == io_state_in_7 ? 8'hf0 : _GEN_1814; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1816 = 8'h18 == io_state_in_7 ? 8'had : _GEN_1815; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1817 = 8'h19 == io_state_in_7 ? 8'hd4 : _GEN_1816; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1818 = 8'h1a == io_state_in_7 ? 8'ha2 : _GEN_1817; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1819 = 8'h1b == io_state_in_7 ? 8'haf : _GEN_1818; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1820 = 8'h1c == io_state_in_7 ? 8'h9c : _GEN_1819; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1821 = 8'h1d == io_state_in_7 ? 8'ha4 : _GEN_1820; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1822 = 8'h1e == io_state_in_7 ? 8'h72 : _GEN_1821; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1823 = 8'h1f == io_state_in_7 ? 8'hc0 : _GEN_1822; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1824 = 8'h20 == io_state_in_7 ? 8'hb7 : _GEN_1823; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1825 = 8'h21 == io_state_in_7 ? 8'hfd : _GEN_1824; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1826 = 8'h22 == io_state_in_7 ? 8'h93 : _GEN_1825; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1827 = 8'h23 == io_state_in_7 ? 8'h26 : _GEN_1826; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1828 = 8'h24 == io_state_in_7 ? 8'h36 : _GEN_1827; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1829 = 8'h25 == io_state_in_7 ? 8'h3f : _GEN_1828; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1830 = 8'h26 == io_state_in_7 ? 8'hf7 : _GEN_1829; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1831 = 8'h27 == io_state_in_7 ? 8'hcc : _GEN_1830; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1832 = 8'h28 == io_state_in_7 ? 8'h34 : _GEN_1831; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1833 = 8'h29 == io_state_in_7 ? 8'ha5 : _GEN_1832; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1834 = 8'h2a == io_state_in_7 ? 8'he5 : _GEN_1833; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1835 = 8'h2b == io_state_in_7 ? 8'hf1 : _GEN_1834; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1836 = 8'h2c == io_state_in_7 ? 8'h71 : _GEN_1835; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1837 = 8'h2d == io_state_in_7 ? 8'hd8 : _GEN_1836; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1838 = 8'h2e == io_state_in_7 ? 8'h31 : _GEN_1837; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1839 = 8'h2f == io_state_in_7 ? 8'h15 : _GEN_1838; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1840 = 8'h30 == io_state_in_7 ? 8'h4 : _GEN_1839; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1841 = 8'h31 == io_state_in_7 ? 8'hc7 : _GEN_1840; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1842 = 8'h32 == io_state_in_7 ? 8'h23 : _GEN_1841; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1843 = 8'h33 == io_state_in_7 ? 8'hc3 : _GEN_1842; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1844 = 8'h34 == io_state_in_7 ? 8'h18 : _GEN_1843; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1845 = 8'h35 == io_state_in_7 ? 8'h96 : _GEN_1844; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1846 = 8'h36 == io_state_in_7 ? 8'h5 : _GEN_1845; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1847 = 8'h37 == io_state_in_7 ? 8'h9a : _GEN_1846; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1848 = 8'h38 == io_state_in_7 ? 8'h7 : _GEN_1847; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1849 = 8'h39 == io_state_in_7 ? 8'h12 : _GEN_1848; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1850 = 8'h3a == io_state_in_7 ? 8'h80 : _GEN_1849; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1851 = 8'h3b == io_state_in_7 ? 8'he2 : _GEN_1850; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1852 = 8'h3c == io_state_in_7 ? 8'heb : _GEN_1851; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1853 = 8'h3d == io_state_in_7 ? 8'h27 : _GEN_1852; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1854 = 8'h3e == io_state_in_7 ? 8'hb2 : _GEN_1853; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1855 = 8'h3f == io_state_in_7 ? 8'h75 : _GEN_1854; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1856 = 8'h40 == io_state_in_7 ? 8'h9 : _GEN_1855; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1857 = 8'h41 == io_state_in_7 ? 8'h83 : _GEN_1856; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1858 = 8'h42 == io_state_in_7 ? 8'h2c : _GEN_1857; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1859 = 8'h43 == io_state_in_7 ? 8'h1a : _GEN_1858; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1860 = 8'h44 == io_state_in_7 ? 8'h1b : _GEN_1859; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1861 = 8'h45 == io_state_in_7 ? 8'h6e : _GEN_1860; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1862 = 8'h46 == io_state_in_7 ? 8'h5a : _GEN_1861; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1863 = 8'h47 == io_state_in_7 ? 8'ha0 : _GEN_1862; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1864 = 8'h48 == io_state_in_7 ? 8'h52 : _GEN_1863; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1865 = 8'h49 == io_state_in_7 ? 8'h3b : _GEN_1864; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1866 = 8'h4a == io_state_in_7 ? 8'hd6 : _GEN_1865; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1867 = 8'h4b == io_state_in_7 ? 8'hb3 : _GEN_1866; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1868 = 8'h4c == io_state_in_7 ? 8'h29 : _GEN_1867; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1869 = 8'h4d == io_state_in_7 ? 8'he3 : _GEN_1868; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1870 = 8'h4e == io_state_in_7 ? 8'h2f : _GEN_1869; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1871 = 8'h4f == io_state_in_7 ? 8'h84 : _GEN_1870; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1872 = 8'h50 == io_state_in_7 ? 8'h53 : _GEN_1871; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1873 = 8'h51 == io_state_in_7 ? 8'hd1 : _GEN_1872; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1874 = 8'h52 == io_state_in_7 ? 8'h0 : _GEN_1873; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1875 = 8'h53 == io_state_in_7 ? 8'hed : _GEN_1874; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1876 = 8'h54 == io_state_in_7 ? 8'h20 : _GEN_1875; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1877 = 8'h55 == io_state_in_7 ? 8'hfc : _GEN_1876; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1878 = 8'h56 == io_state_in_7 ? 8'hb1 : _GEN_1877; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1879 = 8'h57 == io_state_in_7 ? 8'h5b : _GEN_1878; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1880 = 8'h58 == io_state_in_7 ? 8'h6a : _GEN_1879; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1881 = 8'h59 == io_state_in_7 ? 8'hcb : _GEN_1880; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1882 = 8'h5a == io_state_in_7 ? 8'hbe : _GEN_1881; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1883 = 8'h5b == io_state_in_7 ? 8'h39 : _GEN_1882; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1884 = 8'h5c == io_state_in_7 ? 8'h4a : _GEN_1883; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1885 = 8'h5d == io_state_in_7 ? 8'h4c : _GEN_1884; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1886 = 8'h5e == io_state_in_7 ? 8'h58 : _GEN_1885; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1887 = 8'h5f == io_state_in_7 ? 8'hcf : _GEN_1886; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1888 = 8'h60 == io_state_in_7 ? 8'hd0 : _GEN_1887; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1889 = 8'h61 == io_state_in_7 ? 8'hef : _GEN_1888; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1890 = 8'h62 == io_state_in_7 ? 8'haa : _GEN_1889; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1891 = 8'h63 == io_state_in_7 ? 8'hfb : _GEN_1890; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1892 = 8'h64 == io_state_in_7 ? 8'h43 : _GEN_1891; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1893 = 8'h65 == io_state_in_7 ? 8'h4d : _GEN_1892; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1894 = 8'h66 == io_state_in_7 ? 8'h33 : _GEN_1893; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1895 = 8'h67 == io_state_in_7 ? 8'h85 : _GEN_1894; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1896 = 8'h68 == io_state_in_7 ? 8'h45 : _GEN_1895; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1897 = 8'h69 == io_state_in_7 ? 8'hf9 : _GEN_1896; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1898 = 8'h6a == io_state_in_7 ? 8'h2 : _GEN_1897; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1899 = 8'h6b == io_state_in_7 ? 8'h7f : _GEN_1898; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1900 = 8'h6c == io_state_in_7 ? 8'h50 : _GEN_1899; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1901 = 8'h6d == io_state_in_7 ? 8'h3c : _GEN_1900; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1902 = 8'h6e == io_state_in_7 ? 8'h9f : _GEN_1901; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1903 = 8'h6f == io_state_in_7 ? 8'ha8 : _GEN_1902; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1904 = 8'h70 == io_state_in_7 ? 8'h51 : _GEN_1903; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1905 = 8'h71 == io_state_in_7 ? 8'ha3 : _GEN_1904; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1906 = 8'h72 == io_state_in_7 ? 8'h40 : _GEN_1905; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1907 = 8'h73 == io_state_in_7 ? 8'h8f : _GEN_1906; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1908 = 8'h74 == io_state_in_7 ? 8'h92 : _GEN_1907; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1909 = 8'h75 == io_state_in_7 ? 8'h9d : _GEN_1908; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1910 = 8'h76 == io_state_in_7 ? 8'h38 : _GEN_1909; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1911 = 8'h77 == io_state_in_7 ? 8'hf5 : _GEN_1910; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1912 = 8'h78 == io_state_in_7 ? 8'hbc : _GEN_1911; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1913 = 8'h79 == io_state_in_7 ? 8'hb6 : _GEN_1912; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1914 = 8'h7a == io_state_in_7 ? 8'hda : _GEN_1913; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1915 = 8'h7b == io_state_in_7 ? 8'h21 : _GEN_1914; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1916 = 8'h7c == io_state_in_7 ? 8'h10 : _GEN_1915; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1917 = 8'h7d == io_state_in_7 ? 8'hff : _GEN_1916; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1918 = 8'h7e == io_state_in_7 ? 8'hf3 : _GEN_1917; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1919 = 8'h7f == io_state_in_7 ? 8'hd2 : _GEN_1918; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1920 = 8'h80 == io_state_in_7 ? 8'hcd : _GEN_1919; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1921 = 8'h81 == io_state_in_7 ? 8'hc : _GEN_1920; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1922 = 8'h82 == io_state_in_7 ? 8'h13 : _GEN_1921; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1923 = 8'h83 == io_state_in_7 ? 8'hec : _GEN_1922; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1924 = 8'h84 == io_state_in_7 ? 8'h5f : _GEN_1923; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1925 = 8'h85 == io_state_in_7 ? 8'h97 : _GEN_1924; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1926 = 8'h86 == io_state_in_7 ? 8'h44 : _GEN_1925; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1927 = 8'h87 == io_state_in_7 ? 8'h17 : _GEN_1926; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1928 = 8'h88 == io_state_in_7 ? 8'hc4 : _GEN_1927; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1929 = 8'h89 == io_state_in_7 ? 8'ha7 : _GEN_1928; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1930 = 8'h8a == io_state_in_7 ? 8'h7e : _GEN_1929; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1931 = 8'h8b == io_state_in_7 ? 8'h3d : _GEN_1930; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1932 = 8'h8c == io_state_in_7 ? 8'h64 : _GEN_1931; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1933 = 8'h8d == io_state_in_7 ? 8'h5d : _GEN_1932; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1934 = 8'h8e == io_state_in_7 ? 8'h19 : _GEN_1933; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1935 = 8'h8f == io_state_in_7 ? 8'h73 : _GEN_1934; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1936 = 8'h90 == io_state_in_7 ? 8'h60 : _GEN_1935; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1937 = 8'h91 == io_state_in_7 ? 8'h81 : _GEN_1936; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1938 = 8'h92 == io_state_in_7 ? 8'h4f : _GEN_1937; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1939 = 8'h93 == io_state_in_7 ? 8'hdc : _GEN_1938; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1940 = 8'h94 == io_state_in_7 ? 8'h22 : _GEN_1939; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1941 = 8'h95 == io_state_in_7 ? 8'h2a : _GEN_1940; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1942 = 8'h96 == io_state_in_7 ? 8'h90 : _GEN_1941; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1943 = 8'h97 == io_state_in_7 ? 8'h88 : _GEN_1942; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1944 = 8'h98 == io_state_in_7 ? 8'h46 : _GEN_1943; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1945 = 8'h99 == io_state_in_7 ? 8'hee : _GEN_1944; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1946 = 8'h9a == io_state_in_7 ? 8'hb8 : _GEN_1945; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1947 = 8'h9b == io_state_in_7 ? 8'h14 : _GEN_1946; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1948 = 8'h9c == io_state_in_7 ? 8'hde : _GEN_1947; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1949 = 8'h9d == io_state_in_7 ? 8'h5e : _GEN_1948; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1950 = 8'h9e == io_state_in_7 ? 8'hb : _GEN_1949; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1951 = 8'h9f == io_state_in_7 ? 8'hdb : _GEN_1950; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1952 = 8'ha0 == io_state_in_7 ? 8'he0 : _GEN_1951; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1953 = 8'ha1 == io_state_in_7 ? 8'h32 : _GEN_1952; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1954 = 8'ha2 == io_state_in_7 ? 8'h3a : _GEN_1953; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1955 = 8'ha3 == io_state_in_7 ? 8'ha : _GEN_1954; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1956 = 8'ha4 == io_state_in_7 ? 8'h49 : _GEN_1955; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1957 = 8'ha5 == io_state_in_7 ? 8'h6 : _GEN_1956; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1958 = 8'ha6 == io_state_in_7 ? 8'h24 : _GEN_1957; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1959 = 8'ha7 == io_state_in_7 ? 8'h5c : _GEN_1958; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1960 = 8'ha8 == io_state_in_7 ? 8'hc2 : _GEN_1959; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1961 = 8'ha9 == io_state_in_7 ? 8'hd3 : _GEN_1960; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1962 = 8'haa == io_state_in_7 ? 8'hac : _GEN_1961; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1963 = 8'hab == io_state_in_7 ? 8'h62 : _GEN_1962; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1964 = 8'hac == io_state_in_7 ? 8'h91 : _GEN_1963; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1965 = 8'had == io_state_in_7 ? 8'h95 : _GEN_1964; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1966 = 8'hae == io_state_in_7 ? 8'he4 : _GEN_1965; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1967 = 8'haf == io_state_in_7 ? 8'h79 : _GEN_1966; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1968 = 8'hb0 == io_state_in_7 ? 8'he7 : _GEN_1967; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1969 = 8'hb1 == io_state_in_7 ? 8'hc8 : _GEN_1968; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1970 = 8'hb2 == io_state_in_7 ? 8'h37 : _GEN_1969; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1971 = 8'hb3 == io_state_in_7 ? 8'h6d : _GEN_1970; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1972 = 8'hb4 == io_state_in_7 ? 8'h8d : _GEN_1971; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1973 = 8'hb5 == io_state_in_7 ? 8'hd5 : _GEN_1972; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1974 = 8'hb6 == io_state_in_7 ? 8'h4e : _GEN_1973; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1975 = 8'hb7 == io_state_in_7 ? 8'ha9 : _GEN_1974; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1976 = 8'hb8 == io_state_in_7 ? 8'h6c : _GEN_1975; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1977 = 8'hb9 == io_state_in_7 ? 8'h56 : _GEN_1976; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1978 = 8'hba == io_state_in_7 ? 8'hf4 : _GEN_1977; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1979 = 8'hbb == io_state_in_7 ? 8'hea : _GEN_1978; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1980 = 8'hbc == io_state_in_7 ? 8'h65 : _GEN_1979; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1981 = 8'hbd == io_state_in_7 ? 8'h7a : _GEN_1980; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1982 = 8'hbe == io_state_in_7 ? 8'hae : _GEN_1981; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1983 = 8'hbf == io_state_in_7 ? 8'h8 : _GEN_1982; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1984 = 8'hc0 == io_state_in_7 ? 8'hba : _GEN_1983; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1985 = 8'hc1 == io_state_in_7 ? 8'h78 : _GEN_1984; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1986 = 8'hc2 == io_state_in_7 ? 8'h25 : _GEN_1985; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1987 = 8'hc3 == io_state_in_7 ? 8'h2e : _GEN_1986; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1988 = 8'hc4 == io_state_in_7 ? 8'h1c : _GEN_1987; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1989 = 8'hc5 == io_state_in_7 ? 8'ha6 : _GEN_1988; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1990 = 8'hc6 == io_state_in_7 ? 8'hb4 : _GEN_1989; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1991 = 8'hc7 == io_state_in_7 ? 8'hc6 : _GEN_1990; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1992 = 8'hc8 == io_state_in_7 ? 8'he8 : _GEN_1991; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1993 = 8'hc9 == io_state_in_7 ? 8'hdd : _GEN_1992; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1994 = 8'hca == io_state_in_7 ? 8'h74 : _GEN_1993; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1995 = 8'hcb == io_state_in_7 ? 8'h1f : _GEN_1994; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1996 = 8'hcc == io_state_in_7 ? 8'h4b : _GEN_1995; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1997 = 8'hcd == io_state_in_7 ? 8'hbd : _GEN_1996; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1998 = 8'hce == io_state_in_7 ? 8'h8b : _GEN_1997; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_1999 = 8'hcf == io_state_in_7 ? 8'h8a : _GEN_1998; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2000 = 8'hd0 == io_state_in_7 ? 8'h70 : _GEN_1999; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2001 = 8'hd1 == io_state_in_7 ? 8'h3e : _GEN_2000; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2002 = 8'hd2 == io_state_in_7 ? 8'hb5 : _GEN_2001; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2003 = 8'hd3 == io_state_in_7 ? 8'h66 : _GEN_2002; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2004 = 8'hd4 == io_state_in_7 ? 8'h48 : _GEN_2003; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2005 = 8'hd5 == io_state_in_7 ? 8'h3 : _GEN_2004; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2006 = 8'hd6 == io_state_in_7 ? 8'hf6 : _GEN_2005; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2007 = 8'hd7 == io_state_in_7 ? 8'he : _GEN_2006; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2008 = 8'hd8 == io_state_in_7 ? 8'h61 : _GEN_2007; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2009 = 8'hd9 == io_state_in_7 ? 8'h35 : _GEN_2008; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2010 = 8'hda == io_state_in_7 ? 8'h57 : _GEN_2009; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2011 = 8'hdb == io_state_in_7 ? 8'hb9 : _GEN_2010; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2012 = 8'hdc == io_state_in_7 ? 8'h86 : _GEN_2011; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2013 = 8'hdd == io_state_in_7 ? 8'hc1 : _GEN_2012; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2014 = 8'hde == io_state_in_7 ? 8'h1d : _GEN_2013; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2015 = 8'hdf == io_state_in_7 ? 8'h9e : _GEN_2014; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2016 = 8'he0 == io_state_in_7 ? 8'he1 : _GEN_2015; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2017 = 8'he1 == io_state_in_7 ? 8'hf8 : _GEN_2016; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2018 = 8'he2 == io_state_in_7 ? 8'h98 : _GEN_2017; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2019 = 8'he3 == io_state_in_7 ? 8'h11 : _GEN_2018; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2020 = 8'he4 == io_state_in_7 ? 8'h69 : _GEN_2019; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2021 = 8'he5 == io_state_in_7 ? 8'hd9 : _GEN_2020; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2022 = 8'he6 == io_state_in_7 ? 8'h8e : _GEN_2021; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2023 = 8'he7 == io_state_in_7 ? 8'h94 : _GEN_2022; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2024 = 8'he8 == io_state_in_7 ? 8'h9b : _GEN_2023; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2025 = 8'he9 == io_state_in_7 ? 8'h1e : _GEN_2024; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2026 = 8'hea == io_state_in_7 ? 8'h87 : _GEN_2025; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2027 = 8'heb == io_state_in_7 ? 8'he9 : _GEN_2026; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2028 = 8'hec == io_state_in_7 ? 8'hce : _GEN_2027; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2029 = 8'hed == io_state_in_7 ? 8'h55 : _GEN_2028; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2030 = 8'hee == io_state_in_7 ? 8'h28 : _GEN_2029; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2031 = 8'hef == io_state_in_7 ? 8'hdf : _GEN_2030; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2032 = 8'hf0 == io_state_in_7 ? 8'h8c : _GEN_2031; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2033 = 8'hf1 == io_state_in_7 ? 8'ha1 : _GEN_2032; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2034 = 8'hf2 == io_state_in_7 ? 8'h89 : _GEN_2033; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2035 = 8'hf3 == io_state_in_7 ? 8'hd : _GEN_2034; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2036 = 8'hf4 == io_state_in_7 ? 8'hbf : _GEN_2035; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2037 = 8'hf5 == io_state_in_7 ? 8'he6 : _GEN_2036; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2038 = 8'hf6 == io_state_in_7 ? 8'h42 : _GEN_2037; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2039 = 8'hf7 == io_state_in_7 ? 8'h68 : _GEN_2038; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2040 = 8'hf8 == io_state_in_7 ? 8'h41 : _GEN_2039; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2041 = 8'hf9 == io_state_in_7 ? 8'h99 : _GEN_2040; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2042 = 8'hfa == io_state_in_7 ? 8'h2d : _GEN_2041; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2043 = 8'hfb == io_state_in_7 ? 8'hf : _GEN_2042; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2044 = 8'hfc == io_state_in_7 ? 8'hb0 : _GEN_2043; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2045 = 8'hfd == io_state_in_7 ? 8'h54 : _GEN_2044; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2046 = 8'hfe == io_state_in_7 ? 8'hbb : _GEN_2045; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2049 = 8'h1 == io_state_in_8 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2050 = 8'h2 == io_state_in_8 ? 8'h77 : _GEN_2049; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2051 = 8'h3 == io_state_in_8 ? 8'h7b : _GEN_2050; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2052 = 8'h4 == io_state_in_8 ? 8'hf2 : _GEN_2051; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2053 = 8'h5 == io_state_in_8 ? 8'h6b : _GEN_2052; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2054 = 8'h6 == io_state_in_8 ? 8'h6f : _GEN_2053; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2055 = 8'h7 == io_state_in_8 ? 8'hc5 : _GEN_2054; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2056 = 8'h8 == io_state_in_8 ? 8'h30 : _GEN_2055; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2057 = 8'h9 == io_state_in_8 ? 8'h1 : _GEN_2056; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2058 = 8'ha == io_state_in_8 ? 8'h67 : _GEN_2057; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2059 = 8'hb == io_state_in_8 ? 8'h2b : _GEN_2058; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2060 = 8'hc == io_state_in_8 ? 8'hfe : _GEN_2059; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2061 = 8'hd == io_state_in_8 ? 8'hd7 : _GEN_2060; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2062 = 8'he == io_state_in_8 ? 8'hab : _GEN_2061; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2063 = 8'hf == io_state_in_8 ? 8'h76 : _GEN_2062; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2064 = 8'h10 == io_state_in_8 ? 8'hca : _GEN_2063; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2065 = 8'h11 == io_state_in_8 ? 8'h82 : _GEN_2064; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2066 = 8'h12 == io_state_in_8 ? 8'hc9 : _GEN_2065; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2067 = 8'h13 == io_state_in_8 ? 8'h7d : _GEN_2066; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2068 = 8'h14 == io_state_in_8 ? 8'hfa : _GEN_2067; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2069 = 8'h15 == io_state_in_8 ? 8'h59 : _GEN_2068; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2070 = 8'h16 == io_state_in_8 ? 8'h47 : _GEN_2069; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2071 = 8'h17 == io_state_in_8 ? 8'hf0 : _GEN_2070; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2072 = 8'h18 == io_state_in_8 ? 8'had : _GEN_2071; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2073 = 8'h19 == io_state_in_8 ? 8'hd4 : _GEN_2072; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2074 = 8'h1a == io_state_in_8 ? 8'ha2 : _GEN_2073; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2075 = 8'h1b == io_state_in_8 ? 8'haf : _GEN_2074; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2076 = 8'h1c == io_state_in_8 ? 8'h9c : _GEN_2075; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2077 = 8'h1d == io_state_in_8 ? 8'ha4 : _GEN_2076; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2078 = 8'h1e == io_state_in_8 ? 8'h72 : _GEN_2077; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2079 = 8'h1f == io_state_in_8 ? 8'hc0 : _GEN_2078; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2080 = 8'h20 == io_state_in_8 ? 8'hb7 : _GEN_2079; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2081 = 8'h21 == io_state_in_8 ? 8'hfd : _GEN_2080; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2082 = 8'h22 == io_state_in_8 ? 8'h93 : _GEN_2081; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2083 = 8'h23 == io_state_in_8 ? 8'h26 : _GEN_2082; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2084 = 8'h24 == io_state_in_8 ? 8'h36 : _GEN_2083; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2085 = 8'h25 == io_state_in_8 ? 8'h3f : _GEN_2084; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2086 = 8'h26 == io_state_in_8 ? 8'hf7 : _GEN_2085; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2087 = 8'h27 == io_state_in_8 ? 8'hcc : _GEN_2086; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2088 = 8'h28 == io_state_in_8 ? 8'h34 : _GEN_2087; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2089 = 8'h29 == io_state_in_8 ? 8'ha5 : _GEN_2088; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2090 = 8'h2a == io_state_in_8 ? 8'he5 : _GEN_2089; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2091 = 8'h2b == io_state_in_8 ? 8'hf1 : _GEN_2090; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2092 = 8'h2c == io_state_in_8 ? 8'h71 : _GEN_2091; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2093 = 8'h2d == io_state_in_8 ? 8'hd8 : _GEN_2092; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2094 = 8'h2e == io_state_in_8 ? 8'h31 : _GEN_2093; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2095 = 8'h2f == io_state_in_8 ? 8'h15 : _GEN_2094; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2096 = 8'h30 == io_state_in_8 ? 8'h4 : _GEN_2095; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2097 = 8'h31 == io_state_in_8 ? 8'hc7 : _GEN_2096; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2098 = 8'h32 == io_state_in_8 ? 8'h23 : _GEN_2097; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2099 = 8'h33 == io_state_in_8 ? 8'hc3 : _GEN_2098; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2100 = 8'h34 == io_state_in_8 ? 8'h18 : _GEN_2099; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2101 = 8'h35 == io_state_in_8 ? 8'h96 : _GEN_2100; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2102 = 8'h36 == io_state_in_8 ? 8'h5 : _GEN_2101; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2103 = 8'h37 == io_state_in_8 ? 8'h9a : _GEN_2102; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2104 = 8'h38 == io_state_in_8 ? 8'h7 : _GEN_2103; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2105 = 8'h39 == io_state_in_8 ? 8'h12 : _GEN_2104; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2106 = 8'h3a == io_state_in_8 ? 8'h80 : _GEN_2105; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2107 = 8'h3b == io_state_in_8 ? 8'he2 : _GEN_2106; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2108 = 8'h3c == io_state_in_8 ? 8'heb : _GEN_2107; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2109 = 8'h3d == io_state_in_8 ? 8'h27 : _GEN_2108; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2110 = 8'h3e == io_state_in_8 ? 8'hb2 : _GEN_2109; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2111 = 8'h3f == io_state_in_8 ? 8'h75 : _GEN_2110; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2112 = 8'h40 == io_state_in_8 ? 8'h9 : _GEN_2111; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2113 = 8'h41 == io_state_in_8 ? 8'h83 : _GEN_2112; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2114 = 8'h42 == io_state_in_8 ? 8'h2c : _GEN_2113; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2115 = 8'h43 == io_state_in_8 ? 8'h1a : _GEN_2114; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2116 = 8'h44 == io_state_in_8 ? 8'h1b : _GEN_2115; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2117 = 8'h45 == io_state_in_8 ? 8'h6e : _GEN_2116; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2118 = 8'h46 == io_state_in_8 ? 8'h5a : _GEN_2117; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2119 = 8'h47 == io_state_in_8 ? 8'ha0 : _GEN_2118; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2120 = 8'h48 == io_state_in_8 ? 8'h52 : _GEN_2119; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2121 = 8'h49 == io_state_in_8 ? 8'h3b : _GEN_2120; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2122 = 8'h4a == io_state_in_8 ? 8'hd6 : _GEN_2121; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2123 = 8'h4b == io_state_in_8 ? 8'hb3 : _GEN_2122; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2124 = 8'h4c == io_state_in_8 ? 8'h29 : _GEN_2123; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2125 = 8'h4d == io_state_in_8 ? 8'he3 : _GEN_2124; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2126 = 8'h4e == io_state_in_8 ? 8'h2f : _GEN_2125; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2127 = 8'h4f == io_state_in_8 ? 8'h84 : _GEN_2126; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2128 = 8'h50 == io_state_in_8 ? 8'h53 : _GEN_2127; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2129 = 8'h51 == io_state_in_8 ? 8'hd1 : _GEN_2128; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2130 = 8'h52 == io_state_in_8 ? 8'h0 : _GEN_2129; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2131 = 8'h53 == io_state_in_8 ? 8'hed : _GEN_2130; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2132 = 8'h54 == io_state_in_8 ? 8'h20 : _GEN_2131; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2133 = 8'h55 == io_state_in_8 ? 8'hfc : _GEN_2132; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2134 = 8'h56 == io_state_in_8 ? 8'hb1 : _GEN_2133; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2135 = 8'h57 == io_state_in_8 ? 8'h5b : _GEN_2134; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2136 = 8'h58 == io_state_in_8 ? 8'h6a : _GEN_2135; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2137 = 8'h59 == io_state_in_8 ? 8'hcb : _GEN_2136; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2138 = 8'h5a == io_state_in_8 ? 8'hbe : _GEN_2137; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2139 = 8'h5b == io_state_in_8 ? 8'h39 : _GEN_2138; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2140 = 8'h5c == io_state_in_8 ? 8'h4a : _GEN_2139; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2141 = 8'h5d == io_state_in_8 ? 8'h4c : _GEN_2140; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2142 = 8'h5e == io_state_in_8 ? 8'h58 : _GEN_2141; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2143 = 8'h5f == io_state_in_8 ? 8'hcf : _GEN_2142; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2144 = 8'h60 == io_state_in_8 ? 8'hd0 : _GEN_2143; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2145 = 8'h61 == io_state_in_8 ? 8'hef : _GEN_2144; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2146 = 8'h62 == io_state_in_8 ? 8'haa : _GEN_2145; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2147 = 8'h63 == io_state_in_8 ? 8'hfb : _GEN_2146; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2148 = 8'h64 == io_state_in_8 ? 8'h43 : _GEN_2147; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2149 = 8'h65 == io_state_in_8 ? 8'h4d : _GEN_2148; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2150 = 8'h66 == io_state_in_8 ? 8'h33 : _GEN_2149; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2151 = 8'h67 == io_state_in_8 ? 8'h85 : _GEN_2150; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2152 = 8'h68 == io_state_in_8 ? 8'h45 : _GEN_2151; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2153 = 8'h69 == io_state_in_8 ? 8'hf9 : _GEN_2152; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2154 = 8'h6a == io_state_in_8 ? 8'h2 : _GEN_2153; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2155 = 8'h6b == io_state_in_8 ? 8'h7f : _GEN_2154; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2156 = 8'h6c == io_state_in_8 ? 8'h50 : _GEN_2155; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2157 = 8'h6d == io_state_in_8 ? 8'h3c : _GEN_2156; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2158 = 8'h6e == io_state_in_8 ? 8'h9f : _GEN_2157; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2159 = 8'h6f == io_state_in_8 ? 8'ha8 : _GEN_2158; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2160 = 8'h70 == io_state_in_8 ? 8'h51 : _GEN_2159; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2161 = 8'h71 == io_state_in_8 ? 8'ha3 : _GEN_2160; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2162 = 8'h72 == io_state_in_8 ? 8'h40 : _GEN_2161; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2163 = 8'h73 == io_state_in_8 ? 8'h8f : _GEN_2162; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2164 = 8'h74 == io_state_in_8 ? 8'h92 : _GEN_2163; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2165 = 8'h75 == io_state_in_8 ? 8'h9d : _GEN_2164; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2166 = 8'h76 == io_state_in_8 ? 8'h38 : _GEN_2165; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2167 = 8'h77 == io_state_in_8 ? 8'hf5 : _GEN_2166; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2168 = 8'h78 == io_state_in_8 ? 8'hbc : _GEN_2167; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2169 = 8'h79 == io_state_in_8 ? 8'hb6 : _GEN_2168; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2170 = 8'h7a == io_state_in_8 ? 8'hda : _GEN_2169; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2171 = 8'h7b == io_state_in_8 ? 8'h21 : _GEN_2170; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2172 = 8'h7c == io_state_in_8 ? 8'h10 : _GEN_2171; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2173 = 8'h7d == io_state_in_8 ? 8'hff : _GEN_2172; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2174 = 8'h7e == io_state_in_8 ? 8'hf3 : _GEN_2173; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2175 = 8'h7f == io_state_in_8 ? 8'hd2 : _GEN_2174; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2176 = 8'h80 == io_state_in_8 ? 8'hcd : _GEN_2175; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2177 = 8'h81 == io_state_in_8 ? 8'hc : _GEN_2176; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2178 = 8'h82 == io_state_in_8 ? 8'h13 : _GEN_2177; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2179 = 8'h83 == io_state_in_8 ? 8'hec : _GEN_2178; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2180 = 8'h84 == io_state_in_8 ? 8'h5f : _GEN_2179; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2181 = 8'h85 == io_state_in_8 ? 8'h97 : _GEN_2180; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2182 = 8'h86 == io_state_in_8 ? 8'h44 : _GEN_2181; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2183 = 8'h87 == io_state_in_8 ? 8'h17 : _GEN_2182; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2184 = 8'h88 == io_state_in_8 ? 8'hc4 : _GEN_2183; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2185 = 8'h89 == io_state_in_8 ? 8'ha7 : _GEN_2184; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2186 = 8'h8a == io_state_in_8 ? 8'h7e : _GEN_2185; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2187 = 8'h8b == io_state_in_8 ? 8'h3d : _GEN_2186; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2188 = 8'h8c == io_state_in_8 ? 8'h64 : _GEN_2187; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2189 = 8'h8d == io_state_in_8 ? 8'h5d : _GEN_2188; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2190 = 8'h8e == io_state_in_8 ? 8'h19 : _GEN_2189; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2191 = 8'h8f == io_state_in_8 ? 8'h73 : _GEN_2190; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2192 = 8'h90 == io_state_in_8 ? 8'h60 : _GEN_2191; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2193 = 8'h91 == io_state_in_8 ? 8'h81 : _GEN_2192; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2194 = 8'h92 == io_state_in_8 ? 8'h4f : _GEN_2193; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2195 = 8'h93 == io_state_in_8 ? 8'hdc : _GEN_2194; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2196 = 8'h94 == io_state_in_8 ? 8'h22 : _GEN_2195; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2197 = 8'h95 == io_state_in_8 ? 8'h2a : _GEN_2196; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2198 = 8'h96 == io_state_in_8 ? 8'h90 : _GEN_2197; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2199 = 8'h97 == io_state_in_8 ? 8'h88 : _GEN_2198; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2200 = 8'h98 == io_state_in_8 ? 8'h46 : _GEN_2199; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2201 = 8'h99 == io_state_in_8 ? 8'hee : _GEN_2200; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2202 = 8'h9a == io_state_in_8 ? 8'hb8 : _GEN_2201; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2203 = 8'h9b == io_state_in_8 ? 8'h14 : _GEN_2202; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2204 = 8'h9c == io_state_in_8 ? 8'hde : _GEN_2203; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2205 = 8'h9d == io_state_in_8 ? 8'h5e : _GEN_2204; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2206 = 8'h9e == io_state_in_8 ? 8'hb : _GEN_2205; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2207 = 8'h9f == io_state_in_8 ? 8'hdb : _GEN_2206; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2208 = 8'ha0 == io_state_in_8 ? 8'he0 : _GEN_2207; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2209 = 8'ha1 == io_state_in_8 ? 8'h32 : _GEN_2208; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2210 = 8'ha2 == io_state_in_8 ? 8'h3a : _GEN_2209; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2211 = 8'ha3 == io_state_in_8 ? 8'ha : _GEN_2210; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2212 = 8'ha4 == io_state_in_8 ? 8'h49 : _GEN_2211; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2213 = 8'ha5 == io_state_in_8 ? 8'h6 : _GEN_2212; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2214 = 8'ha6 == io_state_in_8 ? 8'h24 : _GEN_2213; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2215 = 8'ha7 == io_state_in_8 ? 8'h5c : _GEN_2214; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2216 = 8'ha8 == io_state_in_8 ? 8'hc2 : _GEN_2215; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2217 = 8'ha9 == io_state_in_8 ? 8'hd3 : _GEN_2216; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2218 = 8'haa == io_state_in_8 ? 8'hac : _GEN_2217; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2219 = 8'hab == io_state_in_8 ? 8'h62 : _GEN_2218; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2220 = 8'hac == io_state_in_8 ? 8'h91 : _GEN_2219; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2221 = 8'had == io_state_in_8 ? 8'h95 : _GEN_2220; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2222 = 8'hae == io_state_in_8 ? 8'he4 : _GEN_2221; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2223 = 8'haf == io_state_in_8 ? 8'h79 : _GEN_2222; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2224 = 8'hb0 == io_state_in_8 ? 8'he7 : _GEN_2223; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2225 = 8'hb1 == io_state_in_8 ? 8'hc8 : _GEN_2224; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2226 = 8'hb2 == io_state_in_8 ? 8'h37 : _GEN_2225; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2227 = 8'hb3 == io_state_in_8 ? 8'h6d : _GEN_2226; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2228 = 8'hb4 == io_state_in_8 ? 8'h8d : _GEN_2227; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2229 = 8'hb5 == io_state_in_8 ? 8'hd5 : _GEN_2228; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2230 = 8'hb6 == io_state_in_8 ? 8'h4e : _GEN_2229; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2231 = 8'hb7 == io_state_in_8 ? 8'ha9 : _GEN_2230; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2232 = 8'hb8 == io_state_in_8 ? 8'h6c : _GEN_2231; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2233 = 8'hb9 == io_state_in_8 ? 8'h56 : _GEN_2232; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2234 = 8'hba == io_state_in_8 ? 8'hf4 : _GEN_2233; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2235 = 8'hbb == io_state_in_8 ? 8'hea : _GEN_2234; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2236 = 8'hbc == io_state_in_8 ? 8'h65 : _GEN_2235; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2237 = 8'hbd == io_state_in_8 ? 8'h7a : _GEN_2236; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2238 = 8'hbe == io_state_in_8 ? 8'hae : _GEN_2237; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2239 = 8'hbf == io_state_in_8 ? 8'h8 : _GEN_2238; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2240 = 8'hc0 == io_state_in_8 ? 8'hba : _GEN_2239; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2241 = 8'hc1 == io_state_in_8 ? 8'h78 : _GEN_2240; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2242 = 8'hc2 == io_state_in_8 ? 8'h25 : _GEN_2241; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2243 = 8'hc3 == io_state_in_8 ? 8'h2e : _GEN_2242; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2244 = 8'hc4 == io_state_in_8 ? 8'h1c : _GEN_2243; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2245 = 8'hc5 == io_state_in_8 ? 8'ha6 : _GEN_2244; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2246 = 8'hc6 == io_state_in_8 ? 8'hb4 : _GEN_2245; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2247 = 8'hc7 == io_state_in_8 ? 8'hc6 : _GEN_2246; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2248 = 8'hc8 == io_state_in_8 ? 8'he8 : _GEN_2247; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2249 = 8'hc9 == io_state_in_8 ? 8'hdd : _GEN_2248; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2250 = 8'hca == io_state_in_8 ? 8'h74 : _GEN_2249; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2251 = 8'hcb == io_state_in_8 ? 8'h1f : _GEN_2250; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2252 = 8'hcc == io_state_in_8 ? 8'h4b : _GEN_2251; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2253 = 8'hcd == io_state_in_8 ? 8'hbd : _GEN_2252; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2254 = 8'hce == io_state_in_8 ? 8'h8b : _GEN_2253; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2255 = 8'hcf == io_state_in_8 ? 8'h8a : _GEN_2254; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2256 = 8'hd0 == io_state_in_8 ? 8'h70 : _GEN_2255; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2257 = 8'hd1 == io_state_in_8 ? 8'h3e : _GEN_2256; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2258 = 8'hd2 == io_state_in_8 ? 8'hb5 : _GEN_2257; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2259 = 8'hd3 == io_state_in_8 ? 8'h66 : _GEN_2258; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2260 = 8'hd4 == io_state_in_8 ? 8'h48 : _GEN_2259; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2261 = 8'hd5 == io_state_in_8 ? 8'h3 : _GEN_2260; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2262 = 8'hd6 == io_state_in_8 ? 8'hf6 : _GEN_2261; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2263 = 8'hd7 == io_state_in_8 ? 8'he : _GEN_2262; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2264 = 8'hd8 == io_state_in_8 ? 8'h61 : _GEN_2263; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2265 = 8'hd9 == io_state_in_8 ? 8'h35 : _GEN_2264; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2266 = 8'hda == io_state_in_8 ? 8'h57 : _GEN_2265; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2267 = 8'hdb == io_state_in_8 ? 8'hb9 : _GEN_2266; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2268 = 8'hdc == io_state_in_8 ? 8'h86 : _GEN_2267; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2269 = 8'hdd == io_state_in_8 ? 8'hc1 : _GEN_2268; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2270 = 8'hde == io_state_in_8 ? 8'h1d : _GEN_2269; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2271 = 8'hdf == io_state_in_8 ? 8'h9e : _GEN_2270; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2272 = 8'he0 == io_state_in_8 ? 8'he1 : _GEN_2271; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2273 = 8'he1 == io_state_in_8 ? 8'hf8 : _GEN_2272; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2274 = 8'he2 == io_state_in_8 ? 8'h98 : _GEN_2273; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2275 = 8'he3 == io_state_in_8 ? 8'h11 : _GEN_2274; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2276 = 8'he4 == io_state_in_8 ? 8'h69 : _GEN_2275; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2277 = 8'he5 == io_state_in_8 ? 8'hd9 : _GEN_2276; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2278 = 8'he6 == io_state_in_8 ? 8'h8e : _GEN_2277; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2279 = 8'he7 == io_state_in_8 ? 8'h94 : _GEN_2278; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2280 = 8'he8 == io_state_in_8 ? 8'h9b : _GEN_2279; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2281 = 8'he9 == io_state_in_8 ? 8'h1e : _GEN_2280; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2282 = 8'hea == io_state_in_8 ? 8'h87 : _GEN_2281; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2283 = 8'heb == io_state_in_8 ? 8'he9 : _GEN_2282; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2284 = 8'hec == io_state_in_8 ? 8'hce : _GEN_2283; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2285 = 8'hed == io_state_in_8 ? 8'h55 : _GEN_2284; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2286 = 8'hee == io_state_in_8 ? 8'h28 : _GEN_2285; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2287 = 8'hef == io_state_in_8 ? 8'hdf : _GEN_2286; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2288 = 8'hf0 == io_state_in_8 ? 8'h8c : _GEN_2287; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2289 = 8'hf1 == io_state_in_8 ? 8'ha1 : _GEN_2288; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2290 = 8'hf2 == io_state_in_8 ? 8'h89 : _GEN_2289; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2291 = 8'hf3 == io_state_in_8 ? 8'hd : _GEN_2290; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2292 = 8'hf4 == io_state_in_8 ? 8'hbf : _GEN_2291; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2293 = 8'hf5 == io_state_in_8 ? 8'he6 : _GEN_2292; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2294 = 8'hf6 == io_state_in_8 ? 8'h42 : _GEN_2293; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2295 = 8'hf7 == io_state_in_8 ? 8'h68 : _GEN_2294; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2296 = 8'hf8 == io_state_in_8 ? 8'h41 : _GEN_2295; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2297 = 8'hf9 == io_state_in_8 ? 8'h99 : _GEN_2296; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2298 = 8'hfa == io_state_in_8 ? 8'h2d : _GEN_2297; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2299 = 8'hfb == io_state_in_8 ? 8'hf : _GEN_2298; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2300 = 8'hfc == io_state_in_8 ? 8'hb0 : _GEN_2299; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2301 = 8'hfd == io_state_in_8 ? 8'h54 : _GEN_2300; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2302 = 8'hfe == io_state_in_8 ? 8'hbb : _GEN_2301; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2305 = 8'h1 == io_state_in_9 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2306 = 8'h2 == io_state_in_9 ? 8'h77 : _GEN_2305; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2307 = 8'h3 == io_state_in_9 ? 8'h7b : _GEN_2306; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2308 = 8'h4 == io_state_in_9 ? 8'hf2 : _GEN_2307; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2309 = 8'h5 == io_state_in_9 ? 8'h6b : _GEN_2308; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2310 = 8'h6 == io_state_in_9 ? 8'h6f : _GEN_2309; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2311 = 8'h7 == io_state_in_9 ? 8'hc5 : _GEN_2310; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2312 = 8'h8 == io_state_in_9 ? 8'h30 : _GEN_2311; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2313 = 8'h9 == io_state_in_9 ? 8'h1 : _GEN_2312; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2314 = 8'ha == io_state_in_9 ? 8'h67 : _GEN_2313; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2315 = 8'hb == io_state_in_9 ? 8'h2b : _GEN_2314; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2316 = 8'hc == io_state_in_9 ? 8'hfe : _GEN_2315; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2317 = 8'hd == io_state_in_9 ? 8'hd7 : _GEN_2316; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2318 = 8'he == io_state_in_9 ? 8'hab : _GEN_2317; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2319 = 8'hf == io_state_in_9 ? 8'h76 : _GEN_2318; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2320 = 8'h10 == io_state_in_9 ? 8'hca : _GEN_2319; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2321 = 8'h11 == io_state_in_9 ? 8'h82 : _GEN_2320; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2322 = 8'h12 == io_state_in_9 ? 8'hc9 : _GEN_2321; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2323 = 8'h13 == io_state_in_9 ? 8'h7d : _GEN_2322; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2324 = 8'h14 == io_state_in_9 ? 8'hfa : _GEN_2323; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2325 = 8'h15 == io_state_in_9 ? 8'h59 : _GEN_2324; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2326 = 8'h16 == io_state_in_9 ? 8'h47 : _GEN_2325; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2327 = 8'h17 == io_state_in_9 ? 8'hf0 : _GEN_2326; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2328 = 8'h18 == io_state_in_9 ? 8'had : _GEN_2327; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2329 = 8'h19 == io_state_in_9 ? 8'hd4 : _GEN_2328; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2330 = 8'h1a == io_state_in_9 ? 8'ha2 : _GEN_2329; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2331 = 8'h1b == io_state_in_9 ? 8'haf : _GEN_2330; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2332 = 8'h1c == io_state_in_9 ? 8'h9c : _GEN_2331; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2333 = 8'h1d == io_state_in_9 ? 8'ha4 : _GEN_2332; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2334 = 8'h1e == io_state_in_9 ? 8'h72 : _GEN_2333; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2335 = 8'h1f == io_state_in_9 ? 8'hc0 : _GEN_2334; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2336 = 8'h20 == io_state_in_9 ? 8'hb7 : _GEN_2335; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2337 = 8'h21 == io_state_in_9 ? 8'hfd : _GEN_2336; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2338 = 8'h22 == io_state_in_9 ? 8'h93 : _GEN_2337; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2339 = 8'h23 == io_state_in_9 ? 8'h26 : _GEN_2338; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2340 = 8'h24 == io_state_in_9 ? 8'h36 : _GEN_2339; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2341 = 8'h25 == io_state_in_9 ? 8'h3f : _GEN_2340; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2342 = 8'h26 == io_state_in_9 ? 8'hf7 : _GEN_2341; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2343 = 8'h27 == io_state_in_9 ? 8'hcc : _GEN_2342; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2344 = 8'h28 == io_state_in_9 ? 8'h34 : _GEN_2343; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2345 = 8'h29 == io_state_in_9 ? 8'ha5 : _GEN_2344; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2346 = 8'h2a == io_state_in_9 ? 8'he5 : _GEN_2345; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2347 = 8'h2b == io_state_in_9 ? 8'hf1 : _GEN_2346; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2348 = 8'h2c == io_state_in_9 ? 8'h71 : _GEN_2347; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2349 = 8'h2d == io_state_in_9 ? 8'hd8 : _GEN_2348; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2350 = 8'h2e == io_state_in_9 ? 8'h31 : _GEN_2349; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2351 = 8'h2f == io_state_in_9 ? 8'h15 : _GEN_2350; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2352 = 8'h30 == io_state_in_9 ? 8'h4 : _GEN_2351; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2353 = 8'h31 == io_state_in_9 ? 8'hc7 : _GEN_2352; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2354 = 8'h32 == io_state_in_9 ? 8'h23 : _GEN_2353; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2355 = 8'h33 == io_state_in_9 ? 8'hc3 : _GEN_2354; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2356 = 8'h34 == io_state_in_9 ? 8'h18 : _GEN_2355; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2357 = 8'h35 == io_state_in_9 ? 8'h96 : _GEN_2356; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2358 = 8'h36 == io_state_in_9 ? 8'h5 : _GEN_2357; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2359 = 8'h37 == io_state_in_9 ? 8'h9a : _GEN_2358; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2360 = 8'h38 == io_state_in_9 ? 8'h7 : _GEN_2359; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2361 = 8'h39 == io_state_in_9 ? 8'h12 : _GEN_2360; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2362 = 8'h3a == io_state_in_9 ? 8'h80 : _GEN_2361; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2363 = 8'h3b == io_state_in_9 ? 8'he2 : _GEN_2362; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2364 = 8'h3c == io_state_in_9 ? 8'heb : _GEN_2363; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2365 = 8'h3d == io_state_in_9 ? 8'h27 : _GEN_2364; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2366 = 8'h3e == io_state_in_9 ? 8'hb2 : _GEN_2365; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2367 = 8'h3f == io_state_in_9 ? 8'h75 : _GEN_2366; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2368 = 8'h40 == io_state_in_9 ? 8'h9 : _GEN_2367; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2369 = 8'h41 == io_state_in_9 ? 8'h83 : _GEN_2368; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2370 = 8'h42 == io_state_in_9 ? 8'h2c : _GEN_2369; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2371 = 8'h43 == io_state_in_9 ? 8'h1a : _GEN_2370; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2372 = 8'h44 == io_state_in_9 ? 8'h1b : _GEN_2371; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2373 = 8'h45 == io_state_in_9 ? 8'h6e : _GEN_2372; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2374 = 8'h46 == io_state_in_9 ? 8'h5a : _GEN_2373; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2375 = 8'h47 == io_state_in_9 ? 8'ha0 : _GEN_2374; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2376 = 8'h48 == io_state_in_9 ? 8'h52 : _GEN_2375; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2377 = 8'h49 == io_state_in_9 ? 8'h3b : _GEN_2376; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2378 = 8'h4a == io_state_in_9 ? 8'hd6 : _GEN_2377; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2379 = 8'h4b == io_state_in_9 ? 8'hb3 : _GEN_2378; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2380 = 8'h4c == io_state_in_9 ? 8'h29 : _GEN_2379; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2381 = 8'h4d == io_state_in_9 ? 8'he3 : _GEN_2380; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2382 = 8'h4e == io_state_in_9 ? 8'h2f : _GEN_2381; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2383 = 8'h4f == io_state_in_9 ? 8'h84 : _GEN_2382; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2384 = 8'h50 == io_state_in_9 ? 8'h53 : _GEN_2383; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2385 = 8'h51 == io_state_in_9 ? 8'hd1 : _GEN_2384; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2386 = 8'h52 == io_state_in_9 ? 8'h0 : _GEN_2385; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2387 = 8'h53 == io_state_in_9 ? 8'hed : _GEN_2386; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2388 = 8'h54 == io_state_in_9 ? 8'h20 : _GEN_2387; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2389 = 8'h55 == io_state_in_9 ? 8'hfc : _GEN_2388; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2390 = 8'h56 == io_state_in_9 ? 8'hb1 : _GEN_2389; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2391 = 8'h57 == io_state_in_9 ? 8'h5b : _GEN_2390; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2392 = 8'h58 == io_state_in_9 ? 8'h6a : _GEN_2391; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2393 = 8'h59 == io_state_in_9 ? 8'hcb : _GEN_2392; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2394 = 8'h5a == io_state_in_9 ? 8'hbe : _GEN_2393; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2395 = 8'h5b == io_state_in_9 ? 8'h39 : _GEN_2394; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2396 = 8'h5c == io_state_in_9 ? 8'h4a : _GEN_2395; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2397 = 8'h5d == io_state_in_9 ? 8'h4c : _GEN_2396; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2398 = 8'h5e == io_state_in_9 ? 8'h58 : _GEN_2397; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2399 = 8'h5f == io_state_in_9 ? 8'hcf : _GEN_2398; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2400 = 8'h60 == io_state_in_9 ? 8'hd0 : _GEN_2399; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2401 = 8'h61 == io_state_in_9 ? 8'hef : _GEN_2400; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2402 = 8'h62 == io_state_in_9 ? 8'haa : _GEN_2401; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2403 = 8'h63 == io_state_in_9 ? 8'hfb : _GEN_2402; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2404 = 8'h64 == io_state_in_9 ? 8'h43 : _GEN_2403; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2405 = 8'h65 == io_state_in_9 ? 8'h4d : _GEN_2404; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2406 = 8'h66 == io_state_in_9 ? 8'h33 : _GEN_2405; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2407 = 8'h67 == io_state_in_9 ? 8'h85 : _GEN_2406; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2408 = 8'h68 == io_state_in_9 ? 8'h45 : _GEN_2407; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2409 = 8'h69 == io_state_in_9 ? 8'hf9 : _GEN_2408; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2410 = 8'h6a == io_state_in_9 ? 8'h2 : _GEN_2409; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2411 = 8'h6b == io_state_in_9 ? 8'h7f : _GEN_2410; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2412 = 8'h6c == io_state_in_9 ? 8'h50 : _GEN_2411; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2413 = 8'h6d == io_state_in_9 ? 8'h3c : _GEN_2412; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2414 = 8'h6e == io_state_in_9 ? 8'h9f : _GEN_2413; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2415 = 8'h6f == io_state_in_9 ? 8'ha8 : _GEN_2414; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2416 = 8'h70 == io_state_in_9 ? 8'h51 : _GEN_2415; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2417 = 8'h71 == io_state_in_9 ? 8'ha3 : _GEN_2416; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2418 = 8'h72 == io_state_in_9 ? 8'h40 : _GEN_2417; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2419 = 8'h73 == io_state_in_9 ? 8'h8f : _GEN_2418; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2420 = 8'h74 == io_state_in_9 ? 8'h92 : _GEN_2419; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2421 = 8'h75 == io_state_in_9 ? 8'h9d : _GEN_2420; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2422 = 8'h76 == io_state_in_9 ? 8'h38 : _GEN_2421; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2423 = 8'h77 == io_state_in_9 ? 8'hf5 : _GEN_2422; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2424 = 8'h78 == io_state_in_9 ? 8'hbc : _GEN_2423; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2425 = 8'h79 == io_state_in_9 ? 8'hb6 : _GEN_2424; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2426 = 8'h7a == io_state_in_9 ? 8'hda : _GEN_2425; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2427 = 8'h7b == io_state_in_9 ? 8'h21 : _GEN_2426; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2428 = 8'h7c == io_state_in_9 ? 8'h10 : _GEN_2427; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2429 = 8'h7d == io_state_in_9 ? 8'hff : _GEN_2428; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2430 = 8'h7e == io_state_in_9 ? 8'hf3 : _GEN_2429; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2431 = 8'h7f == io_state_in_9 ? 8'hd2 : _GEN_2430; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2432 = 8'h80 == io_state_in_9 ? 8'hcd : _GEN_2431; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2433 = 8'h81 == io_state_in_9 ? 8'hc : _GEN_2432; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2434 = 8'h82 == io_state_in_9 ? 8'h13 : _GEN_2433; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2435 = 8'h83 == io_state_in_9 ? 8'hec : _GEN_2434; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2436 = 8'h84 == io_state_in_9 ? 8'h5f : _GEN_2435; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2437 = 8'h85 == io_state_in_9 ? 8'h97 : _GEN_2436; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2438 = 8'h86 == io_state_in_9 ? 8'h44 : _GEN_2437; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2439 = 8'h87 == io_state_in_9 ? 8'h17 : _GEN_2438; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2440 = 8'h88 == io_state_in_9 ? 8'hc4 : _GEN_2439; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2441 = 8'h89 == io_state_in_9 ? 8'ha7 : _GEN_2440; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2442 = 8'h8a == io_state_in_9 ? 8'h7e : _GEN_2441; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2443 = 8'h8b == io_state_in_9 ? 8'h3d : _GEN_2442; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2444 = 8'h8c == io_state_in_9 ? 8'h64 : _GEN_2443; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2445 = 8'h8d == io_state_in_9 ? 8'h5d : _GEN_2444; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2446 = 8'h8e == io_state_in_9 ? 8'h19 : _GEN_2445; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2447 = 8'h8f == io_state_in_9 ? 8'h73 : _GEN_2446; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2448 = 8'h90 == io_state_in_9 ? 8'h60 : _GEN_2447; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2449 = 8'h91 == io_state_in_9 ? 8'h81 : _GEN_2448; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2450 = 8'h92 == io_state_in_9 ? 8'h4f : _GEN_2449; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2451 = 8'h93 == io_state_in_9 ? 8'hdc : _GEN_2450; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2452 = 8'h94 == io_state_in_9 ? 8'h22 : _GEN_2451; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2453 = 8'h95 == io_state_in_9 ? 8'h2a : _GEN_2452; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2454 = 8'h96 == io_state_in_9 ? 8'h90 : _GEN_2453; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2455 = 8'h97 == io_state_in_9 ? 8'h88 : _GEN_2454; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2456 = 8'h98 == io_state_in_9 ? 8'h46 : _GEN_2455; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2457 = 8'h99 == io_state_in_9 ? 8'hee : _GEN_2456; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2458 = 8'h9a == io_state_in_9 ? 8'hb8 : _GEN_2457; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2459 = 8'h9b == io_state_in_9 ? 8'h14 : _GEN_2458; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2460 = 8'h9c == io_state_in_9 ? 8'hde : _GEN_2459; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2461 = 8'h9d == io_state_in_9 ? 8'h5e : _GEN_2460; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2462 = 8'h9e == io_state_in_9 ? 8'hb : _GEN_2461; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2463 = 8'h9f == io_state_in_9 ? 8'hdb : _GEN_2462; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2464 = 8'ha0 == io_state_in_9 ? 8'he0 : _GEN_2463; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2465 = 8'ha1 == io_state_in_9 ? 8'h32 : _GEN_2464; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2466 = 8'ha2 == io_state_in_9 ? 8'h3a : _GEN_2465; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2467 = 8'ha3 == io_state_in_9 ? 8'ha : _GEN_2466; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2468 = 8'ha4 == io_state_in_9 ? 8'h49 : _GEN_2467; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2469 = 8'ha5 == io_state_in_9 ? 8'h6 : _GEN_2468; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2470 = 8'ha6 == io_state_in_9 ? 8'h24 : _GEN_2469; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2471 = 8'ha7 == io_state_in_9 ? 8'h5c : _GEN_2470; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2472 = 8'ha8 == io_state_in_9 ? 8'hc2 : _GEN_2471; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2473 = 8'ha9 == io_state_in_9 ? 8'hd3 : _GEN_2472; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2474 = 8'haa == io_state_in_9 ? 8'hac : _GEN_2473; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2475 = 8'hab == io_state_in_9 ? 8'h62 : _GEN_2474; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2476 = 8'hac == io_state_in_9 ? 8'h91 : _GEN_2475; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2477 = 8'had == io_state_in_9 ? 8'h95 : _GEN_2476; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2478 = 8'hae == io_state_in_9 ? 8'he4 : _GEN_2477; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2479 = 8'haf == io_state_in_9 ? 8'h79 : _GEN_2478; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2480 = 8'hb0 == io_state_in_9 ? 8'he7 : _GEN_2479; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2481 = 8'hb1 == io_state_in_9 ? 8'hc8 : _GEN_2480; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2482 = 8'hb2 == io_state_in_9 ? 8'h37 : _GEN_2481; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2483 = 8'hb3 == io_state_in_9 ? 8'h6d : _GEN_2482; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2484 = 8'hb4 == io_state_in_9 ? 8'h8d : _GEN_2483; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2485 = 8'hb5 == io_state_in_9 ? 8'hd5 : _GEN_2484; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2486 = 8'hb6 == io_state_in_9 ? 8'h4e : _GEN_2485; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2487 = 8'hb7 == io_state_in_9 ? 8'ha9 : _GEN_2486; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2488 = 8'hb8 == io_state_in_9 ? 8'h6c : _GEN_2487; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2489 = 8'hb9 == io_state_in_9 ? 8'h56 : _GEN_2488; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2490 = 8'hba == io_state_in_9 ? 8'hf4 : _GEN_2489; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2491 = 8'hbb == io_state_in_9 ? 8'hea : _GEN_2490; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2492 = 8'hbc == io_state_in_9 ? 8'h65 : _GEN_2491; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2493 = 8'hbd == io_state_in_9 ? 8'h7a : _GEN_2492; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2494 = 8'hbe == io_state_in_9 ? 8'hae : _GEN_2493; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2495 = 8'hbf == io_state_in_9 ? 8'h8 : _GEN_2494; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2496 = 8'hc0 == io_state_in_9 ? 8'hba : _GEN_2495; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2497 = 8'hc1 == io_state_in_9 ? 8'h78 : _GEN_2496; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2498 = 8'hc2 == io_state_in_9 ? 8'h25 : _GEN_2497; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2499 = 8'hc3 == io_state_in_9 ? 8'h2e : _GEN_2498; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2500 = 8'hc4 == io_state_in_9 ? 8'h1c : _GEN_2499; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2501 = 8'hc5 == io_state_in_9 ? 8'ha6 : _GEN_2500; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2502 = 8'hc6 == io_state_in_9 ? 8'hb4 : _GEN_2501; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2503 = 8'hc7 == io_state_in_9 ? 8'hc6 : _GEN_2502; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2504 = 8'hc8 == io_state_in_9 ? 8'he8 : _GEN_2503; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2505 = 8'hc9 == io_state_in_9 ? 8'hdd : _GEN_2504; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2506 = 8'hca == io_state_in_9 ? 8'h74 : _GEN_2505; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2507 = 8'hcb == io_state_in_9 ? 8'h1f : _GEN_2506; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2508 = 8'hcc == io_state_in_9 ? 8'h4b : _GEN_2507; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2509 = 8'hcd == io_state_in_9 ? 8'hbd : _GEN_2508; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2510 = 8'hce == io_state_in_9 ? 8'h8b : _GEN_2509; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2511 = 8'hcf == io_state_in_9 ? 8'h8a : _GEN_2510; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2512 = 8'hd0 == io_state_in_9 ? 8'h70 : _GEN_2511; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2513 = 8'hd1 == io_state_in_9 ? 8'h3e : _GEN_2512; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2514 = 8'hd2 == io_state_in_9 ? 8'hb5 : _GEN_2513; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2515 = 8'hd3 == io_state_in_9 ? 8'h66 : _GEN_2514; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2516 = 8'hd4 == io_state_in_9 ? 8'h48 : _GEN_2515; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2517 = 8'hd5 == io_state_in_9 ? 8'h3 : _GEN_2516; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2518 = 8'hd6 == io_state_in_9 ? 8'hf6 : _GEN_2517; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2519 = 8'hd7 == io_state_in_9 ? 8'he : _GEN_2518; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2520 = 8'hd8 == io_state_in_9 ? 8'h61 : _GEN_2519; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2521 = 8'hd9 == io_state_in_9 ? 8'h35 : _GEN_2520; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2522 = 8'hda == io_state_in_9 ? 8'h57 : _GEN_2521; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2523 = 8'hdb == io_state_in_9 ? 8'hb9 : _GEN_2522; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2524 = 8'hdc == io_state_in_9 ? 8'h86 : _GEN_2523; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2525 = 8'hdd == io_state_in_9 ? 8'hc1 : _GEN_2524; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2526 = 8'hde == io_state_in_9 ? 8'h1d : _GEN_2525; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2527 = 8'hdf == io_state_in_9 ? 8'h9e : _GEN_2526; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2528 = 8'he0 == io_state_in_9 ? 8'he1 : _GEN_2527; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2529 = 8'he1 == io_state_in_9 ? 8'hf8 : _GEN_2528; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2530 = 8'he2 == io_state_in_9 ? 8'h98 : _GEN_2529; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2531 = 8'he3 == io_state_in_9 ? 8'h11 : _GEN_2530; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2532 = 8'he4 == io_state_in_9 ? 8'h69 : _GEN_2531; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2533 = 8'he5 == io_state_in_9 ? 8'hd9 : _GEN_2532; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2534 = 8'he6 == io_state_in_9 ? 8'h8e : _GEN_2533; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2535 = 8'he7 == io_state_in_9 ? 8'h94 : _GEN_2534; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2536 = 8'he8 == io_state_in_9 ? 8'h9b : _GEN_2535; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2537 = 8'he9 == io_state_in_9 ? 8'h1e : _GEN_2536; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2538 = 8'hea == io_state_in_9 ? 8'h87 : _GEN_2537; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2539 = 8'heb == io_state_in_9 ? 8'he9 : _GEN_2538; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2540 = 8'hec == io_state_in_9 ? 8'hce : _GEN_2539; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2541 = 8'hed == io_state_in_9 ? 8'h55 : _GEN_2540; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2542 = 8'hee == io_state_in_9 ? 8'h28 : _GEN_2541; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2543 = 8'hef == io_state_in_9 ? 8'hdf : _GEN_2542; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2544 = 8'hf0 == io_state_in_9 ? 8'h8c : _GEN_2543; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2545 = 8'hf1 == io_state_in_9 ? 8'ha1 : _GEN_2544; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2546 = 8'hf2 == io_state_in_9 ? 8'h89 : _GEN_2545; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2547 = 8'hf3 == io_state_in_9 ? 8'hd : _GEN_2546; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2548 = 8'hf4 == io_state_in_9 ? 8'hbf : _GEN_2547; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2549 = 8'hf5 == io_state_in_9 ? 8'he6 : _GEN_2548; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2550 = 8'hf6 == io_state_in_9 ? 8'h42 : _GEN_2549; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2551 = 8'hf7 == io_state_in_9 ? 8'h68 : _GEN_2550; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2552 = 8'hf8 == io_state_in_9 ? 8'h41 : _GEN_2551; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2553 = 8'hf9 == io_state_in_9 ? 8'h99 : _GEN_2552; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2554 = 8'hfa == io_state_in_9 ? 8'h2d : _GEN_2553; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2555 = 8'hfb == io_state_in_9 ? 8'hf : _GEN_2554; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2556 = 8'hfc == io_state_in_9 ? 8'hb0 : _GEN_2555; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2557 = 8'hfd == io_state_in_9 ? 8'h54 : _GEN_2556; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2558 = 8'hfe == io_state_in_9 ? 8'hbb : _GEN_2557; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2561 = 8'h1 == io_state_in_10 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2562 = 8'h2 == io_state_in_10 ? 8'h77 : _GEN_2561; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2563 = 8'h3 == io_state_in_10 ? 8'h7b : _GEN_2562; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2564 = 8'h4 == io_state_in_10 ? 8'hf2 : _GEN_2563; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2565 = 8'h5 == io_state_in_10 ? 8'h6b : _GEN_2564; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2566 = 8'h6 == io_state_in_10 ? 8'h6f : _GEN_2565; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2567 = 8'h7 == io_state_in_10 ? 8'hc5 : _GEN_2566; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2568 = 8'h8 == io_state_in_10 ? 8'h30 : _GEN_2567; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2569 = 8'h9 == io_state_in_10 ? 8'h1 : _GEN_2568; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2570 = 8'ha == io_state_in_10 ? 8'h67 : _GEN_2569; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2571 = 8'hb == io_state_in_10 ? 8'h2b : _GEN_2570; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2572 = 8'hc == io_state_in_10 ? 8'hfe : _GEN_2571; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2573 = 8'hd == io_state_in_10 ? 8'hd7 : _GEN_2572; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2574 = 8'he == io_state_in_10 ? 8'hab : _GEN_2573; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2575 = 8'hf == io_state_in_10 ? 8'h76 : _GEN_2574; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2576 = 8'h10 == io_state_in_10 ? 8'hca : _GEN_2575; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2577 = 8'h11 == io_state_in_10 ? 8'h82 : _GEN_2576; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2578 = 8'h12 == io_state_in_10 ? 8'hc9 : _GEN_2577; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2579 = 8'h13 == io_state_in_10 ? 8'h7d : _GEN_2578; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2580 = 8'h14 == io_state_in_10 ? 8'hfa : _GEN_2579; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2581 = 8'h15 == io_state_in_10 ? 8'h59 : _GEN_2580; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2582 = 8'h16 == io_state_in_10 ? 8'h47 : _GEN_2581; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2583 = 8'h17 == io_state_in_10 ? 8'hf0 : _GEN_2582; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2584 = 8'h18 == io_state_in_10 ? 8'had : _GEN_2583; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2585 = 8'h19 == io_state_in_10 ? 8'hd4 : _GEN_2584; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2586 = 8'h1a == io_state_in_10 ? 8'ha2 : _GEN_2585; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2587 = 8'h1b == io_state_in_10 ? 8'haf : _GEN_2586; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2588 = 8'h1c == io_state_in_10 ? 8'h9c : _GEN_2587; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2589 = 8'h1d == io_state_in_10 ? 8'ha4 : _GEN_2588; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2590 = 8'h1e == io_state_in_10 ? 8'h72 : _GEN_2589; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2591 = 8'h1f == io_state_in_10 ? 8'hc0 : _GEN_2590; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2592 = 8'h20 == io_state_in_10 ? 8'hb7 : _GEN_2591; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2593 = 8'h21 == io_state_in_10 ? 8'hfd : _GEN_2592; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2594 = 8'h22 == io_state_in_10 ? 8'h93 : _GEN_2593; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2595 = 8'h23 == io_state_in_10 ? 8'h26 : _GEN_2594; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2596 = 8'h24 == io_state_in_10 ? 8'h36 : _GEN_2595; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2597 = 8'h25 == io_state_in_10 ? 8'h3f : _GEN_2596; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2598 = 8'h26 == io_state_in_10 ? 8'hf7 : _GEN_2597; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2599 = 8'h27 == io_state_in_10 ? 8'hcc : _GEN_2598; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2600 = 8'h28 == io_state_in_10 ? 8'h34 : _GEN_2599; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2601 = 8'h29 == io_state_in_10 ? 8'ha5 : _GEN_2600; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2602 = 8'h2a == io_state_in_10 ? 8'he5 : _GEN_2601; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2603 = 8'h2b == io_state_in_10 ? 8'hf1 : _GEN_2602; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2604 = 8'h2c == io_state_in_10 ? 8'h71 : _GEN_2603; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2605 = 8'h2d == io_state_in_10 ? 8'hd8 : _GEN_2604; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2606 = 8'h2e == io_state_in_10 ? 8'h31 : _GEN_2605; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2607 = 8'h2f == io_state_in_10 ? 8'h15 : _GEN_2606; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2608 = 8'h30 == io_state_in_10 ? 8'h4 : _GEN_2607; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2609 = 8'h31 == io_state_in_10 ? 8'hc7 : _GEN_2608; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2610 = 8'h32 == io_state_in_10 ? 8'h23 : _GEN_2609; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2611 = 8'h33 == io_state_in_10 ? 8'hc3 : _GEN_2610; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2612 = 8'h34 == io_state_in_10 ? 8'h18 : _GEN_2611; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2613 = 8'h35 == io_state_in_10 ? 8'h96 : _GEN_2612; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2614 = 8'h36 == io_state_in_10 ? 8'h5 : _GEN_2613; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2615 = 8'h37 == io_state_in_10 ? 8'h9a : _GEN_2614; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2616 = 8'h38 == io_state_in_10 ? 8'h7 : _GEN_2615; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2617 = 8'h39 == io_state_in_10 ? 8'h12 : _GEN_2616; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2618 = 8'h3a == io_state_in_10 ? 8'h80 : _GEN_2617; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2619 = 8'h3b == io_state_in_10 ? 8'he2 : _GEN_2618; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2620 = 8'h3c == io_state_in_10 ? 8'heb : _GEN_2619; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2621 = 8'h3d == io_state_in_10 ? 8'h27 : _GEN_2620; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2622 = 8'h3e == io_state_in_10 ? 8'hb2 : _GEN_2621; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2623 = 8'h3f == io_state_in_10 ? 8'h75 : _GEN_2622; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2624 = 8'h40 == io_state_in_10 ? 8'h9 : _GEN_2623; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2625 = 8'h41 == io_state_in_10 ? 8'h83 : _GEN_2624; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2626 = 8'h42 == io_state_in_10 ? 8'h2c : _GEN_2625; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2627 = 8'h43 == io_state_in_10 ? 8'h1a : _GEN_2626; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2628 = 8'h44 == io_state_in_10 ? 8'h1b : _GEN_2627; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2629 = 8'h45 == io_state_in_10 ? 8'h6e : _GEN_2628; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2630 = 8'h46 == io_state_in_10 ? 8'h5a : _GEN_2629; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2631 = 8'h47 == io_state_in_10 ? 8'ha0 : _GEN_2630; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2632 = 8'h48 == io_state_in_10 ? 8'h52 : _GEN_2631; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2633 = 8'h49 == io_state_in_10 ? 8'h3b : _GEN_2632; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2634 = 8'h4a == io_state_in_10 ? 8'hd6 : _GEN_2633; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2635 = 8'h4b == io_state_in_10 ? 8'hb3 : _GEN_2634; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2636 = 8'h4c == io_state_in_10 ? 8'h29 : _GEN_2635; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2637 = 8'h4d == io_state_in_10 ? 8'he3 : _GEN_2636; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2638 = 8'h4e == io_state_in_10 ? 8'h2f : _GEN_2637; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2639 = 8'h4f == io_state_in_10 ? 8'h84 : _GEN_2638; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2640 = 8'h50 == io_state_in_10 ? 8'h53 : _GEN_2639; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2641 = 8'h51 == io_state_in_10 ? 8'hd1 : _GEN_2640; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2642 = 8'h52 == io_state_in_10 ? 8'h0 : _GEN_2641; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2643 = 8'h53 == io_state_in_10 ? 8'hed : _GEN_2642; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2644 = 8'h54 == io_state_in_10 ? 8'h20 : _GEN_2643; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2645 = 8'h55 == io_state_in_10 ? 8'hfc : _GEN_2644; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2646 = 8'h56 == io_state_in_10 ? 8'hb1 : _GEN_2645; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2647 = 8'h57 == io_state_in_10 ? 8'h5b : _GEN_2646; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2648 = 8'h58 == io_state_in_10 ? 8'h6a : _GEN_2647; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2649 = 8'h59 == io_state_in_10 ? 8'hcb : _GEN_2648; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2650 = 8'h5a == io_state_in_10 ? 8'hbe : _GEN_2649; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2651 = 8'h5b == io_state_in_10 ? 8'h39 : _GEN_2650; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2652 = 8'h5c == io_state_in_10 ? 8'h4a : _GEN_2651; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2653 = 8'h5d == io_state_in_10 ? 8'h4c : _GEN_2652; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2654 = 8'h5e == io_state_in_10 ? 8'h58 : _GEN_2653; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2655 = 8'h5f == io_state_in_10 ? 8'hcf : _GEN_2654; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2656 = 8'h60 == io_state_in_10 ? 8'hd0 : _GEN_2655; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2657 = 8'h61 == io_state_in_10 ? 8'hef : _GEN_2656; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2658 = 8'h62 == io_state_in_10 ? 8'haa : _GEN_2657; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2659 = 8'h63 == io_state_in_10 ? 8'hfb : _GEN_2658; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2660 = 8'h64 == io_state_in_10 ? 8'h43 : _GEN_2659; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2661 = 8'h65 == io_state_in_10 ? 8'h4d : _GEN_2660; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2662 = 8'h66 == io_state_in_10 ? 8'h33 : _GEN_2661; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2663 = 8'h67 == io_state_in_10 ? 8'h85 : _GEN_2662; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2664 = 8'h68 == io_state_in_10 ? 8'h45 : _GEN_2663; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2665 = 8'h69 == io_state_in_10 ? 8'hf9 : _GEN_2664; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2666 = 8'h6a == io_state_in_10 ? 8'h2 : _GEN_2665; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2667 = 8'h6b == io_state_in_10 ? 8'h7f : _GEN_2666; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2668 = 8'h6c == io_state_in_10 ? 8'h50 : _GEN_2667; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2669 = 8'h6d == io_state_in_10 ? 8'h3c : _GEN_2668; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2670 = 8'h6e == io_state_in_10 ? 8'h9f : _GEN_2669; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2671 = 8'h6f == io_state_in_10 ? 8'ha8 : _GEN_2670; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2672 = 8'h70 == io_state_in_10 ? 8'h51 : _GEN_2671; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2673 = 8'h71 == io_state_in_10 ? 8'ha3 : _GEN_2672; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2674 = 8'h72 == io_state_in_10 ? 8'h40 : _GEN_2673; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2675 = 8'h73 == io_state_in_10 ? 8'h8f : _GEN_2674; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2676 = 8'h74 == io_state_in_10 ? 8'h92 : _GEN_2675; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2677 = 8'h75 == io_state_in_10 ? 8'h9d : _GEN_2676; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2678 = 8'h76 == io_state_in_10 ? 8'h38 : _GEN_2677; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2679 = 8'h77 == io_state_in_10 ? 8'hf5 : _GEN_2678; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2680 = 8'h78 == io_state_in_10 ? 8'hbc : _GEN_2679; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2681 = 8'h79 == io_state_in_10 ? 8'hb6 : _GEN_2680; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2682 = 8'h7a == io_state_in_10 ? 8'hda : _GEN_2681; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2683 = 8'h7b == io_state_in_10 ? 8'h21 : _GEN_2682; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2684 = 8'h7c == io_state_in_10 ? 8'h10 : _GEN_2683; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2685 = 8'h7d == io_state_in_10 ? 8'hff : _GEN_2684; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2686 = 8'h7e == io_state_in_10 ? 8'hf3 : _GEN_2685; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2687 = 8'h7f == io_state_in_10 ? 8'hd2 : _GEN_2686; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2688 = 8'h80 == io_state_in_10 ? 8'hcd : _GEN_2687; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2689 = 8'h81 == io_state_in_10 ? 8'hc : _GEN_2688; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2690 = 8'h82 == io_state_in_10 ? 8'h13 : _GEN_2689; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2691 = 8'h83 == io_state_in_10 ? 8'hec : _GEN_2690; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2692 = 8'h84 == io_state_in_10 ? 8'h5f : _GEN_2691; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2693 = 8'h85 == io_state_in_10 ? 8'h97 : _GEN_2692; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2694 = 8'h86 == io_state_in_10 ? 8'h44 : _GEN_2693; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2695 = 8'h87 == io_state_in_10 ? 8'h17 : _GEN_2694; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2696 = 8'h88 == io_state_in_10 ? 8'hc4 : _GEN_2695; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2697 = 8'h89 == io_state_in_10 ? 8'ha7 : _GEN_2696; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2698 = 8'h8a == io_state_in_10 ? 8'h7e : _GEN_2697; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2699 = 8'h8b == io_state_in_10 ? 8'h3d : _GEN_2698; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2700 = 8'h8c == io_state_in_10 ? 8'h64 : _GEN_2699; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2701 = 8'h8d == io_state_in_10 ? 8'h5d : _GEN_2700; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2702 = 8'h8e == io_state_in_10 ? 8'h19 : _GEN_2701; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2703 = 8'h8f == io_state_in_10 ? 8'h73 : _GEN_2702; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2704 = 8'h90 == io_state_in_10 ? 8'h60 : _GEN_2703; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2705 = 8'h91 == io_state_in_10 ? 8'h81 : _GEN_2704; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2706 = 8'h92 == io_state_in_10 ? 8'h4f : _GEN_2705; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2707 = 8'h93 == io_state_in_10 ? 8'hdc : _GEN_2706; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2708 = 8'h94 == io_state_in_10 ? 8'h22 : _GEN_2707; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2709 = 8'h95 == io_state_in_10 ? 8'h2a : _GEN_2708; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2710 = 8'h96 == io_state_in_10 ? 8'h90 : _GEN_2709; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2711 = 8'h97 == io_state_in_10 ? 8'h88 : _GEN_2710; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2712 = 8'h98 == io_state_in_10 ? 8'h46 : _GEN_2711; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2713 = 8'h99 == io_state_in_10 ? 8'hee : _GEN_2712; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2714 = 8'h9a == io_state_in_10 ? 8'hb8 : _GEN_2713; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2715 = 8'h9b == io_state_in_10 ? 8'h14 : _GEN_2714; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2716 = 8'h9c == io_state_in_10 ? 8'hde : _GEN_2715; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2717 = 8'h9d == io_state_in_10 ? 8'h5e : _GEN_2716; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2718 = 8'h9e == io_state_in_10 ? 8'hb : _GEN_2717; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2719 = 8'h9f == io_state_in_10 ? 8'hdb : _GEN_2718; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2720 = 8'ha0 == io_state_in_10 ? 8'he0 : _GEN_2719; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2721 = 8'ha1 == io_state_in_10 ? 8'h32 : _GEN_2720; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2722 = 8'ha2 == io_state_in_10 ? 8'h3a : _GEN_2721; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2723 = 8'ha3 == io_state_in_10 ? 8'ha : _GEN_2722; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2724 = 8'ha4 == io_state_in_10 ? 8'h49 : _GEN_2723; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2725 = 8'ha5 == io_state_in_10 ? 8'h6 : _GEN_2724; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2726 = 8'ha6 == io_state_in_10 ? 8'h24 : _GEN_2725; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2727 = 8'ha7 == io_state_in_10 ? 8'h5c : _GEN_2726; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2728 = 8'ha8 == io_state_in_10 ? 8'hc2 : _GEN_2727; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2729 = 8'ha9 == io_state_in_10 ? 8'hd3 : _GEN_2728; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2730 = 8'haa == io_state_in_10 ? 8'hac : _GEN_2729; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2731 = 8'hab == io_state_in_10 ? 8'h62 : _GEN_2730; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2732 = 8'hac == io_state_in_10 ? 8'h91 : _GEN_2731; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2733 = 8'had == io_state_in_10 ? 8'h95 : _GEN_2732; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2734 = 8'hae == io_state_in_10 ? 8'he4 : _GEN_2733; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2735 = 8'haf == io_state_in_10 ? 8'h79 : _GEN_2734; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2736 = 8'hb0 == io_state_in_10 ? 8'he7 : _GEN_2735; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2737 = 8'hb1 == io_state_in_10 ? 8'hc8 : _GEN_2736; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2738 = 8'hb2 == io_state_in_10 ? 8'h37 : _GEN_2737; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2739 = 8'hb3 == io_state_in_10 ? 8'h6d : _GEN_2738; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2740 = 8'hb4 == io_state_in_10 ? 8'h8d : _GEN_2739; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2741 = 8'hb5 == io_state_in_10 ? 8'hd5 : _GEN_2740; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2742 = 8'hb6 == io_state_in_10 ? 8'h4e : _GEN_2741; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2743 = 8'hb7 == io_state_in_10 ? 8'ha9 : _GEN_2742; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2744 = 8'hb8 == io_state_in_10 ? 8'h6c : _GEN_2743; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2745 = 8'hb9 == io_state_in_10 ? 8'h56 : _GEN_2744; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2746 = 8'hba == io_state_in_10 ? 8'hf4 : _GEN_2745; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2747 = 8'hbb == io_state_in_10 ? 8'hea : _GEN_2746; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2748 = 8'hbc == io_state_in_10 ? 8'h65 : _GEN_2747; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2749 = 8'hbd == io_state_in_10 ? 8'h7a : _GEN_2748; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2750 = 8'hbe == io_state_in_10 ? 8'hae : _GEN_2749; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2751 = 8'hbf == io_state_in_10 ? 8'h8 : _GEN_2750; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2752 = 8'hc0 == io_state_in_10 ? 8'hba : _GEN_2751; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2753 = 8'hc1 == io_state_in_10 ? 8'h78 : _GEN_2752; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2754 = 8'hc2 == io_state_in_10 ? 8'h25 : _GEN_2753; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2755 = 8'hc3 == io_state_in_10 ? 8'h2e : _GEN_2754; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2756 = 8'hc4 == io_state_in_10 ? 8'h1c : _GEN_2755; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2757 = 8'hc5 == io_state_in_10 ? 8'ha6 : _GEN_2756; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2758 = 8'hc6 == io_state_in_10 ? 8'hb4 : _GEN_2757; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2759 = 8'hc7 == io_state_in_10 ? 8'hc6 : _GEN_2758; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2760 = 8'hc8 == io_state_in_10 ? 8'he8 : _GEN_2759; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2761 = 8'hc9 == io_state_in_10 ? 8'hdd : _GEN_2760; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2762 = 8'hca == io_state_in_10 ? 8'h74 : _GEN_2761; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2763 = 8'hcb == io_state_in_10 ? 8'h1f : _GEN_2762; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2764 = 8'hcc == io_state_in_10 ? 8'h4b : _GEN_2763; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2765 = 8'hcd == io_state_in_10 ? 8'hbd : _GEN_2764; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2766 = 8'hce == io_state_in_10 ? 8'h8b : _GEN_2765; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2767 = 8'hcf == io_state_in_10 ? 8'h8a : _GEN_2766; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2768 = 8'hd0 == io_state_in_10 ? 8'h70 : _GEN_2767; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2769 = 8'hd1 == io_state_in_10 ? 8'h3e : _GEN_2768; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2770 = 8'hd2 == io_state_in_10 ? 8'hb5 : _GEN_2769; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2771 = 8'hd3 == io_state_in_10 ? 8'h66 : _GEN_2770; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2772 = 8'hd4 == io_state_in_10 ? 8'h48 : _GEN_2771; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2773 = 8'hd5 == io_state_in_10 ? 8'h3 : _GEN_2772; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2774 = 8'hd6 == io_state_in_10 ? 8'hf6 : _GEN_2773; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2775 = 8'hd7 == io_state_in_10 ? 8'he : _GEN_2774; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2776 = 8'hd8 == io_state_in_10 ? 8'h61 : _GEN_2775; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2777 = 8'hd9 == io_state_in_10 ? 8'h35 : _GEN_2776; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2778 = 8'hda == io_state_in_10 ? 8'h57 : _GEN_2777; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2779 = 8'hdb == io_state_in_10 ? 8'hb9 : _GEN_2778; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2780 = 8'hdc == io_state_in_10 ? 8'h86 : _GEN_2779; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2781 = 8'hdd == io_state_in_10 ? 8'hc1 : _GEN_2780; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2782 = 8'hde == io_state_in_10 ? 8'h1d : _GEN_2781; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2783 = 8'hdf == io_state_in_10 ? 8'h9e : _GEN_2782; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2784 = 8'he0 == io_state_in_10 ? 8'he1 : _GEN_2783; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2785 = 8'he1 == io_state_in_10 ? 8'hf8 : _GEN_2784; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2786 = 8'he2 == io_state_in_10 ? 8'h98 : _GEN_2785; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2787 = 8'he3 == io_state_in_10 ? 8'h11 : _GEN_2786; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2788 = 8'he4 == io_state_in_10 ? 8'h69 : _GEN_2787; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2789 = 8'he5 == io_state_in_10 ? 8'hd9 : _GEN_2788; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2790 = 8'he6 == io_state_in_10 ? 8'h8e : _GEN_2789; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2791 = 8'he7 == io_state_in_10 ? 8'h94 : _GEN_2790; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2792 = 8'he8 == io_state_in_10 ? 8'h9b : _GEN_2791; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2793 = 8'he9 == io_state_in_10 ? 8'h1e : _GEN_2792; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2794 = 8'hea == io_state_in_10 ? 8'h87 : _GEN_2793; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2795 = 8'heb == io_state_in_10 ? 8'he9 : _GEN_2794; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2796 = 8'hec == io_state_in_10 ? 8'hce : _GEN_2795; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2797 = 8'hed == io_state_in_10 ? 8'h55 : _GEN_2796; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2798 = 8'hee == io_state_in_10 ? 8'h28 : _GEN_2797; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2799 = 8'hef == io_state_in_10 ? 8'hdf : _GEN_2798; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2800 = 8'hf0 == io_state_in_10 ? 8'h8c : _GEN_2799; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2801 = 8'hf1 == io_state_in_10 ? 8'ha1 : _GEN_2800; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2802 = 8'hf2 == io_state_in_10 ? 8'h89 : _GEN_2801; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2803 = 8'hf3 == io_state_in_10 ? 8'hd : _GEN_2802; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2804 = 8'hf4 == io_state_in_10 ? 8'hbf : _GEN_2803; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2805 = 8'hf5 == io_state_in_10 ? 8'he6 : _GEN_2804; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2806 = 8'hf6 == io_state_in_10 ? 8'h42 : _GEN_2805; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2807 = 8'hf7 == io_state_in_10 ? 8'h68 : _GEN_2806; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2808 = 8'hf8 == io_state_in_10 ? 8'h41 : _GEN_2807; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2809 = 8'hf9 == io_state_in_10 ? 8'h99 : _GEN_2808; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2810 = 8'hfa == io_state_in_10 ? 8'h2d : _GEN_2809; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2811 = 8'hfb == io_state_in_10 ? 8'hf : _GEN_2810; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2812 = 8'hfc == io_state_in_10 ? 8'hb0 : _GEN_2811; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2813 = 8'hfd == io_state_in_10 ? 8'h54 : _GEN_2812; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2814 = 8'hfe == io_state_in_10 ? 8'hbb : _GEN_2813; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2817 = 8'h1 == io_state_in_11 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2818 = 8'h2 == io_state_in_11 ? 8'h77 : _GEN_2817; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2819 = 8'h3 == io_state_in_11 ? 8'h7b : _GEN_2818; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2820 = 8'h4 == io_state_in_11 ? 8'hf2 : _GEN_2819; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2821 = 8'h5 == io_state_in_11 ? 8'h6b : _GEN_2820; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2822 = 8'h6 == io_state_in_11 ? 8'h6f : _GEN_2821; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2823 = 8'h7 == io_state_in_11 ? 8'hc5 : _GEN_2822; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2824 = 8'h8 == io_state_in_11 ? 8'h30 : _GEN_2823; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2825 = 8'h9 == io_state_in_11 ? 8'h1 : _GEN_2824; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2826 = 8'ha == io_state_in_11 ? 8'h67 : _GEN_2825; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2827 = 8'hb == io_state_in_11 ? 8'h2b : _GEN_2826; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2828 = 8'hc == io_state_in_11 ? 8'hfe : _GEN_2827; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2829 = 8'hd == io_state_in_11 ? 8'hd7 : _GEN_2828; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2830 = 8'he == io_state_in_11 ? 8'hab : _GEN_2829; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2831 = 8'hf == io_state_in_11 ? 8'h76 : _GEN_2830; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2832 = 8'h10 == io_state_in_11 ? 8'hca : _GEN_2831; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2833 = 8'h11 == io_state_in_11 ? 8'h82 : _GEN_2832; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2834 = 8'h12 == io_state_in_11 ? 8'hc9 : _GEN_2833; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2835 = 8'h13 == io_state_in_11 ? 8'h7d : _GEN_2834; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2836 = 8'h14 == io_state_in_11 ? 8'hfa : _GEN_2835; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2837 = 8'h15 == io_state_in_11 ? 8'h59 : _GEN_2836; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2838 = 8'h16 == io_state_in_11 ? 8'h47 : _GEN_2837; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2839 = 8'h17 == io_state_in_11 ? 8'hf0 : _GEN_2838; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2840 = 8'h18 == io_state_in_11 ? 8'had : _GEN_2839; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2841 = 8'h19 == io_state_in_11 ? 8'hd4 : _GEN_2840; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2842 = 8'h1a == io_state_in_11 ? 8'ha2 : _GEN_2841; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2843 = 8'h1b == io_state_in_11 ? 8'haf : _GEN_2842; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2844 = 8'h1c == io_state_in_11 ? 8'h9c : _GEN_2843; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2845 = 8'h1d == io_state_in_11 ? 8'ha4 : _GEN_2844; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2846 = 8'h1e == io_state_in_11 ? 8'h72 : _GEN_2845; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2847 = 8'h1f == io_state_in_11 ? 8'hc0 : _GEN_2846; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2848 = 8'h20 == io_state_in_11 ? 8'hb7 : _GEN_2847; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2849 = 8'h21 == io_state_in_11 ? 8'hfd : _GEN_2848; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2850 = 8'h22 == io_state_in_11 ? 8'h93 : _GEN_2849; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2851 = 8'h23 == io_state_in_11 ? 8'h26 : _GEN_2850; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2852 = 8'h24 == io_state_in_11 ? 8'h36 : _GEN_2851; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2853 = 8'h25 == io_state_in_11 ? 8'h3f : _GEN_2852; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2854 = 8'h26 == io_state_in_11 ? 8'hf7 : _GEN_2853; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2855 = 8'h27 == io_state_in_11 ? 8'hcc : _GEN_2854; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2856 = 8'h28 == io_state_in_11 ? 8'h34 : _GEN_2855; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2857 = 8'h29 == io_state_in_11 ? 8'ha5 : _GEN_2856; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2858 = 8'h2a == io_state_in_11 ? 8'he5 : _GEN_2857; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2859 = 8'h2b == io_state_in_11 ? 8'hf1 : _GEN_2858; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2860 = 8'h2c == io_state_in_11 ? 8'h71 : _GEN_2859; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2861 = 8'h2d == io_state_in_11 ? 8'hd8 : _GEN_2860; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2862 = 8'h2e == io_state_in_11 ? 8'h31 : _GEN_2861; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2863 = 8'h2f == io_state_in_11 ? 8'h15 : _GEN_2862; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2864 = 8'h30 == io_state_in_11 ? 8'h4 : _GEN_2863; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2865 = 8'h31 == io_state_in_11 ? 8'hc7 : _GEN_2864; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2866 = 8'h32 == io_state_in_11 ? 8'h23 : _GEN_2865; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2867 = 8'h33 == io_state_in_11 ? 8'hc3 : _GEN_2866; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2868 = 8'h34 == io_state_in_11 ? 8'h18 : _GEN_2867; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2869 = 8'h35 == io_state_in_11 ? 8'h96 : _GEN_2868; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2870 = 8'h36 == io_state_in_11 ? 8'h5 : _GEN_2869; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2871 = 8'h37 == io_state_in_11 ? 8'h9a : _GEN_2870; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2872 = 8'h38 == io_state_in_11 ? 8'h7 : _GEN_2871; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2873 = 8'h39 == io_state_in_11 ? 8'h12 : _GEN_2872; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2874 = 8'h3a == io_state_in_11 ? 8'h80 : _GEN_2873; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2875 = 8'h3b == io_state_in_11 ? 8'he2 : _GEN_2874; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2876 = 8'h3c == io_state_in_11 ? 8'heb : _GEN_2875; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2877 = 8'h3d == io_state_in_11 ? 8'h27 : _GEN_2876; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2878 = 8'h3e == io_state_in_11 ? 8'hb2 : _GEN_2877; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2879 = 8'h3f == io_state_in_11 ? 8'h75 : _GEN_2878; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2880 = 8'h40 == io_state_in_11 ? 8'h9 : _GEN_2879; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2881 = 8'h41 == io_state_in_11 ? 8'h83 : _GEN_2880; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2882 = 8'h42 == io_state_in_11 ? 8'h2c : _GEN_2881; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2883 = 8'h43 == io_state_in_11 ? 8'h1a : _GEN_2882; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2884 = 8'h44 == io_state_in_11 ? 8'h1b : _GEN_2883; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2885 = 8'h45 == io_state_in_11 ? 8'h6e : _GEN_2884; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2886 = 8'h46 == io_state_in_11 ? 8'h5a : _GEN_2885; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2887 = 8'h47 == io_state_in_11 ? 8'ha0 : _GEN_2886; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2888 = 8'h48 == io_state_in_11 ? 8'h52 : _GEN_2887; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2889 = 8'h49 == io_state_in_11 ? 8'h3b : _GEN_2888; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2890 = 8'h4a == io_state_in_11 ? 8'hd6 : _GEN_2889; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2891 = 8'h4b == io_state_in_11 ? 8'hb3 : _GEN_2890; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2892 = 8'h4c == io_state_in_11 ? 8'h29 : _GEN_2891; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2893 = 8'h4d == io_state_in_11 ? 8'he3 : _GEN_2892; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2894 = 8'h4e == io_state_in_11 ? 8'h2f : _GEN_2893; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2895 = 8'h4f == io_state_in_11 ? 8'h84 : _GEN_2894; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2896 = 8'h50 == io_state_in_11 ? 8'h53 : _GEN_2895; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2897 = 8'h51 == io_state_in_11 ? 8'hd1 : _GEN_2896; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2898 = 8'h52 == io_state_in_11 ? 8'h0 : _GEN_2897; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2899 = 8'h53 == io_state_in_11 ? 8'hed : _GEN_2898; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2900 = 8'h54 == io_state_in_11 ? 8'h20 : _GEN_2899; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2901 = 8'h55 == io_state_in_11 ? 8'hfc : _GEN_2900; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2902 = 8'h56 == io_state_in_11 ? 8'hb1 : _GEN_2901; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2903 = 8'h57 == io_state_in_11 ? 8'h5b : _GEN_2902; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2904 = 8'h58 == io_state_in_11 ? 8'h6a : _GEN_2903; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2905 = 8'h59 == io_state_in_11 ? 8'hcb : _GEN_2904; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2906 = 8'h5a == io_state_in_11 ? 8'hbe : _GEN_2905; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2907 = 8'h5b == io_state_in_11 ? 8'h39 : _GEN_2906; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2908 = 8'h5c == io_state_in_11 ? 8'h4a : _GEN_2907; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2909 = 8'h5d == io_state_in_11 ? 8'h4c : _GEN_2908; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2910 = 8'h5e == io_state_in_11 ? 8'h58 : _GEN_2909; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2911 = 8'h5f == io_state_in_11 ? 8'hcf : _GEN_2910; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2912 = 8'h60 == io_state_in_11 ? 8'hd0 : _GEN_2911; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2913 = 8'h61 == io_state_in_11 ? 8'hef : _GEN_2912; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2914 = 8'h62 == io_state_in_11 ? 8'haa : _GEN_2913; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2915 = 8'h63 == io_state_in_11 ? 8'hfb : _GEN_2914; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2916 = 8'h64 == io_state_in_11 ? 8'h43 : _GEN_2915; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2917 = 8'h65 == io_state_in_11 ? 8'h4d : _GEN_2916; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2918 = 8'h66 == io_state_in_11 ? 8'h33 : _GEN_2917; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2919 = 8'h67 == io_state_in_11 ? 8'h85 : _GEN_2918; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2920 = 8'h68 == io_state_in_11 ? 8'h45 : _GEN_2919; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2921 = 8'h69 == io_state_in_11 ? 8'hf9 : _GEN_2920; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2922 = 8'h6a == io_state_in_11 ? 8'h2 : _GEN_2921; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2923 = 8'h6b == io_state_in_11 ? 8'h7f : _GEN_2922; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2924 = 8'h6c == io_state_in_11 ? 8'h50 : _GEN_2923; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2925 = 8'h6d == io_state_in_11 ? 8'h3c : _GEN_2924; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2926 = 8'h6e == io_state_in_11 ? 8'h9f : _GEN_2925; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2927 = 8'h6f == io_state_in_11 ? 8'ha8 : _GEN_2926; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2928 = 8'h70 == io_state_in_11 ? 8'h51 : _GEN_2927; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2929 = 8'h71 == io_state_in_11 ? 8'ha3 : _GEN_2928; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2930 = 8'h72 == io_state_in_11 ? 8'h40 : _GEN_2929; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2931 = 8'h73 == io_state_in_11 ? 8'h8f : _GEN_2930; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2932 = 8'h74 == io_state_in_11 ? 8'h92 : _GEN_2931; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2933 = 8'h75 == io_state_in_11 ? 8'h9d : _GEN_2932; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2934 = 8'h76 == io_state_in_11 ? 8'h38 : _GEN_2933; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2935 = 8'h77 == io_state_in_11 ? 8'hf5 : _GEN_2934; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2936 = 8'h78 == io_state_in_11 ? 8'hbc : _GEN_2935; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2937 = 8'h79 == io_state_in_11 ? 8'hb6 : _GEN_2936; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2938 = 8'h7a == io_state_in_11 ? 8'hda : _GEN_2937; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2939 = 8'h7b == io_state_in_11 ? 8'h21 : _GEN_2938; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2940 = 8'h7c == io_state_in_11 ? 8'h10 : _GEN_2939; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2941 = 8'h7d == io_state_in_11 ? 8'hff : _GEN_2940; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2942 = 8'h7e == io_state_in_11 ? 8'hf3 : _GEN_2941; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2943 = 8'h7f == io_state_in_11 ? 8'hd2 : _GEN_2942; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2944 = 8'h80 == io_state_in_11 ? 8'hcd : _GEN_2943; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2945 = 8'h81 == io_state_in_11 ? 8'hc : _GEN_2944; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2946 = 8'h82 == io_state_in_11 ? 8'h13 : _GEN_2945; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2947 = 8'h83 == io_state_in_11 ? 8'hec : _GEN_2946; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2948 = 8'h84 == io_state_in_11 ? 8'h5f : _GEN_2947; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2949 = 8'h85 == io_state_in_11 ? 8'h97 : _GEN_2948; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2950 = 8'h86 == io_state_in_11 ? 8'h44 : _GEN_2949; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2951 = 8'h87 == io_state_in_11 ? 8'h17 : _GEN_2950; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2952 = 8'h88 == io_state_in_11 ? 8'hc4 : _GEN_2951; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2953 = 8'h89 == io_state_in_11 ? 8'ha7 : _GEN_2952; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2954 = 8'h8a == io_state_in_11 ? 8'h7e : _GEN_2953; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2955 = 8'h8b == io_state_in_11 ? 8'h3d : _GEN_2954; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2956 = 8'h8c == io_state_in_11 ? 8'h64 : _GEN_2955; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2957 = 8'h8d == io_state_in_11 ? 8'h5d : _GEN_2956; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2958 = 8'h8e == io_state_in_11 ? 8'h19 : _GEN_2957; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2959 = 8'h8f == io_state_in_11 ? 8'h73 : _GEN_2958; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2960 = 8'h90 == io_state_in_11 ? 8'h60 : _GEN_2959; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2961 = 8'h91 == io_state_in_11 ? 8'h81 : _GEN_2960; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2962 = 8'h92 == io_state_in_11 ? 8'h4f : _GEN_2961; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2963 = 8'h93 == io_state_in_11 ? 8'hdc : _GEN_2962; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2964 = 8'h94 == io_state_in_11 ? 8'h22 : _GEN_2963; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2965 = 8'h95 == io_state_in_11 ? 8'h2a : _GEN_2964; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2966 = 8'h96 == io_state_in_11 ? 8'h90 : _GEN_2965; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2967 = 8'h97 == io_state_in_11 ? 8'h88 : _GEN_2966; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2968 = 8'h98 == io_state_in_11 ? 8'h46 : _GEN_2967; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2969 = 8'h99 == io_state_in_11 ? 8'hee : _GEN_2968; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2970 = 8'h9a == io_state_in_11 ? 8'hb8 : _GEN_2969; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2971 = 8'h9b == io_state_in_11 ? 8'h14 : _GEN_2970; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2972 = 8'h9c == io_state_in_11 ? 8'hde : _GEN_2971; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2973 = 8'h9d == io_state_in_11 ? 8'h5e : _GEN_2972; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2974 = 8'h9e == io_state_in_11 ? 8'hb : _GEN_2973; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2975 = 8'h9f == io_state_in_11 ? 8'hdb : _GEN_2974; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2976 = 8'ha0 == io_state_in_11 ? 8'he0 : _GEN_2975; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2977 = 8'ha1 == io_state_in_11 ? 8'h32 : _GEN_2976; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2978 = 8'ha2 == io_state_in_11 ? 8'h3a : _GEN_2977; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2979 = 8'ha3 == io_state_in_11 ? 8'ha : _GEN_2978; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2980 = 8'ha4 == io_state_in_11 ? 8'h49 : _GEN_2979; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2981 = 8'ha5 == io_state_in_11 ? 8'h6 : _GEN_2980; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2982 = 8'ha6 == io_state_in_11 ? 8'h24 : _GEN_2981; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2983 = 8'ha7 == io_state_in_11 ? 8'h5c : _GEN_2982; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2984 = 8'ha8 == io_state_in_11 ? 8'hc2 : _GEN_2983; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2985 = 8'ha9 == io_state_in_11 ? 8'hd3 : _GEN_2984; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2986 = 8'haa == io_state_in_11 ? 8'hac : _GEN_2985; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2987 = 8'hab == io_state_in_11 ? 8'h62 : _GEN_2986; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2988 = 8'hac == io_state_in_11 ? 8'h91 : _GEN_2987; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2989 = 8'had == io_state_in_11 ? 8'h95 : _GEN_2988; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2990 = 8'hae == io_state_in_11 ? 8'he4 : _GEN_2989; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2991 = 8'haf == io_state_in_11 ? 8'h79 : _GEN_2990; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2992 = 8'hb0 == io_state_in_11 ? 8'he7 : _GEN_2991; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2993 = 8'hb1 == io_state_in_11 ? 8'hc8 : _GEN_2992; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2994 = 8'hb2 == io_state_in_11 ? 8'h37 : _GEN_2993; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2995 = 8'hb3 == io_state_in_11 ? 8'h6d : _GEN_2994; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2996 = 8'hb4 == io_state_in_11 ? 8'h8d : _GEN_2995; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2997 = 8'hb5 == io_state_in_11 ? 8'hd5 : _GEN_2996; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2998 = 8'hb6 == io_state_in_11 ? 8'h4e : _GEN_2997; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_2999 = 8'hb7 == io_state_in_11 ? 8'ha9 : _GEN_2998; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3000 = 8'hb8 == io_state_in_11 ? 8'h6c : _GEN_2999; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3001 = 8'hb9 == io_state_in_11 ? 8'h56 : _GEN_3000; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3002 = 8'hba == io_state_in_11 ? 8'hf4 : _GEN_3001; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3003 = 8'hbb == io_state_in_11 ? 8'hea : _GEN_3002; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3004 = 8'hbc == io_state_in_11 ? 8'h65 : _GEN_3003; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3005 = 8'hbd == io_state_in_11 ? 8'h7a : _GEN_3004; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3006 = 8'hbe == io_state_in_11 ? 8'hae : _GEN_3005; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3007 = 8'hbf == io_state_in_11 ? 8'h8 : _GEN_3006; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3008 = 8'hc0 == io_state_in_11 ? 8'hba : _GEN_3007; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3009 = 8'hc1 == io_state_in_11 ? 8'h78 : _GEN_3008; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3010 = 8'hc2 == io_state_in_11 ? 8'h25 : _GEN_3009; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3011 = 8'hc3 == io_state_in_11 ? 8'h2e : _GEN_3010; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3012 = 8'hc4 == io_state_in_11 ? 8'h1c : _GEN_3011; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3013 = 8'hc5 == io_state_in_11 ? 8'ha6 : _GEN_3012; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3014 = 8'hc6 == io_state_in_11 ? 8'hb4 : _GEN_3013; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3015 = 8'hc7 == io_state_in_11 ? 8'hc6 : _GEN_3014; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3016 = 8'hc8 == io_state_in_11 ? 8'he8 : _GEN_3015; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3017 = 8'hc9 == io_state_in_11 ? 8'hdd : _GEN_3016; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3018 = 8'hca == io_state_in_11 ? 8'h74 : _GEN_3017; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3019 = 8'hcb == io_state_in_11 ? 8'h1f : _GEN_3018; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3020 = 8'hcc == io_state_in_11 ? 8'h4b : _GEN_3019; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3021 = 8'hcd == io_state_in_11 ? 8'hbd : _GEN_3020; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3022 = 8'hce == io_state_in_11 ? 8'h8b : _GEN_3021; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3023 = 8'hcf == io_state_in_11 ? 8'h8a : _GEN_3022; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3024 = 8'hd0 == io_state_in_11 ? 8'h70 : _GEN_3023; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3025 = 8'hd1 == io_state_in_11 ? 8'h3e : _GEN_3024; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3026 = 8'hd2 == io_state_in_11 ? 8'hb5 : _GEN_3025; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3027 = 8'hd3 == io_state_in_11 ? 8'h66 : _GEN_3026; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3028 = 8'hd4 == io_state_in_11 ? 8'h48 : _GEN_3027; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3029 = 8'hd5 == io_state_in_11 ? 8'h3 : _GEN_3028; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3030 = 8'hd6 == io_state_in_11 ? 8'hf6 : _GEN_3029; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3031 = 8'hd7 == io_state_in_11 ? 8'he : _GEN_3030; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3032 = 8'hd8 == io_state_in_11 ? 8'h61 : _GEN_3031; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3033 = 8'hd9 == io_state_in_11 ? 8'h35 : _GEN_3032; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3034 = 8'hda == io_state_in_11 ? 8'h57 : _GEN_3033; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3035 = 8'hdb == io_state_in_11 ? 8'hb9 : _GEN_3034; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3036 = 8'hdc == io_state_in_11 ? 8'h86 : _GEN_3035; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3037 = 8'hdd == io_state_in_11 ? 8'hc1 : _GEN_3036; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3038 = 8'hde == io_state_in_11 ? 8'h1d : _GEN_3037; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3039 = 8'hdf == io_state_in_11 ? 8'h9e : _GEN_3038; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3040 = 8'he0 == io_state_in_11 ? 8'he1 : _GEN_3039; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3041 = 8'he1 == io_state_in_11 ? 8'hf8 : _GEN_3040; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3042 = 8'he2 == io_state_in_11 ? 8'h98 : _GEN_3041; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3043 = 8'he3 == io_state_in_11 ? 8'h11 : _GEN_3042; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3044 = 8'he4 == io_state_in_11 ? 8'h69 : _GEN_3043; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3045 = 8'he5 == io_state_in_11 ? 8'hd9 : _GEN_3044; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3046 = 8'he6 == io_state_in_11 ? 8'h8e : _GEN_3045; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3047 = 8'he7 == io_state_in_11 ? 8'h94 : _GEN_3046; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3048 = 8'he8 == io_state_in_11 ? 8'h9b : _GEN_3047; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3049 = 8'he9 == io_state_in_11 ? 8'h1e : _GEN_3048; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3050 = 8'hea == io_state_in_11 ? 8'h87 : _GEN_3049; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3051 = 8'heb == io_state_in_11 ? 8'he9 : _GEN_3050; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3052 = 8'hec == io_state_in_11 ? 8'hce : _GEN_3051; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3053 = 8'hed == io_state_in_11 ? 8'h55 : _GEN_3052; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3054 = 8'hee == io_state_in_11 ? 8'h28 : _GEN_3053; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3055 = 8'hef == io_state_in_11 ? 8'hdf : _GEN_3054; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3056 = 8'hf0 == io_state_in_11 ? 8'h8c : _GEN_3055; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3057 = 8'hf1 == io_state_in_11 ? 8'ha1 : _GEN_3056; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3058 = 8'hf2 == io_state_in_11 ? 8'h89 : _GEN_3057; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3059 = 8'hf3 == io_state_in_11 ? 8'hd : _GEN_3058; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3060 = 8'hf4 == io_state_in_11 ? 8'hbf : _GEN_3059; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3061 = 8'hf5 == io_state_in_11 ? 8'he6 : _GEN_3060; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3062 = 8'hf6 == io_state_in_11 ? 8'h42 : _GEN_3061; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3063 = 8'hf7 == io_state_in_11 ? 8'h68 : _GEN_3062; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3064 = 8'hf8 == io_state_in_11 ? 8'h41 : _GEN_3063; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3065 = 8'hf9 == io_state_in_11 ? 8'h99 : _GEN_3064; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3066 = 8'hfa == io_state_in_11 ? 8'h2d : _GEN_3065; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3067 = 8'hfb == io_state_in_11 ? 8'hf : _GEN_3066; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3068 = 8'hfc == io_state_in_11 ? 8'hb0 : _GEN_3067; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3069 = 8'hfd == io_state_in_11 ? 8'h54 : _GEN_3068; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3070 = 8'hfe == io_state_in_11 ? 8'hbb : _GEN_3069; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3073 = 8'h1 == io_state_in_12 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3074 = 8'h2 == io_state_in_12 ? 8'h77 : _GEN_3073; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3075 = 8'h3 == io_state_in_12 ? 8'h7b : _GEN_3074; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3076 = 8'h4 == io_state_in_12 ? 8'hf2 : _GEN_3075; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3077 = 8'h5 == io_state_in_12 ? 8'h6b : _GEN_3076; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3078 = 8'h6 == io_state_in_12 ? 8'h6f : _GEN_3077; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3079 = 8'h7 == io_state_in_12 ? 8'hc5 : _GEN_3078; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3080 = 8'h8 == io_state_in_12 ? 8'h30 : _GEN_3079; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3081 = 8'h9 == io_state_in_12 ? 8'h1 : _GEN_3080; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3082 = 8'ha == io_state_in_12 ? 8'h67 : _GEN_3081; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3083 = 8'hb == io_state_in_12 ? 8'h2b : _GEN_3082; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3084 = 8'hc == io_state_in_12 ? 8'hfe : _GEN_3083; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3085 = 8'hd == io_state_in_12 ? 8'hd7 : _GEN_3084; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3086 = 8'he == io_state_in_12 ? 8'hab : _GEN_3085; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3087 = 8'hf == io_state_in_12 ? 8'h76 : _GEN_3086; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3088 = 8'h10 == io_state_in_12 ? 8'hca : _GEN_3087; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3089 = 8'h11 == io_state_in_12 ? 8'h82 : _GEN_3088; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3090 = 8'h12 == io_state_in_12 ? 8'hc9 : _GEN_3089; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3091 = 8'h13 == io_state_in_12 ? 8'h7d : _GEN_3090; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3092 = 8'h14 == io_state_in_12 ? 8'hfa : _GEN_3091; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3093 = 8'h15 == io_state_in_12 ? 8'h59 : _GEN_3092; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3094 = 8'h16 == io_state_in_12 ? 8'h47 : _GEN_3093; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3095 = 8'h17 == io_state_in_12 ? 8'hf0 : _GEN_3094; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3096 = 8'h18 == io_state_in_12 ? 8'had : _GEN_3095; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3097 = 8'h19 == io_state_in_12 ? 8'hd4 : _GEN_3096; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3098 = 8'h1a == io_state_in_12 ? 8'ha2 : _GEN_3097; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3099 = 8'h1b == io_state_in_12 ? 8'haf : _GEN_3098; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3100 = 8'h1c == io_state_in_12 ? 8'h9c : _GEN_3099; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3101 = 8'h1d == io_state_in_12 ? 8'ha4 : _GEN_3100; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3102 = 8'h1e == io_state_in_12 ? 8'h72 : _GEN_3101; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3103 = 8'h1f == io_state_in_12 ? 8'hc0 : _GEN_3102; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3104 = 8'h20 == io_state_in_12 ? 8'hb7 : _GEN_3103; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3105 = 8'h21 == io_state_in_12 ? 8'hfd : _GEN_3104; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3106 = 8'h22 == io_state_in_12 ? 8'h93 : _GEN_3105; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3107 = 8'h23 == io_state_in_12 ? 8'h26 : _GEN_3106; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3108 = 8'h24 == io_state_in_12 ? 8'h36 : _GEN_3107; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3109 = 8'h25 == io_state_in_12 ? 8'h3f : _GEN_3108; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3110 = 8'h26 == io_state_in_12 ? 8'hf7 : _GEN_3109; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3111 = 8'h27 == io_state_in_12 ? 8'hcc : _GEN_3110; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3112 = 8'h28 == io_state_in_12 ? 8'h34 : _GEN_3111; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3113 = 8'h29 == io_state_in_12 ? 8'ha5 : _GEN_3112; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3114 = 8'h2a == io_state_in_12 ? 8'he5 : _GEN_3113; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3115 = 8'h2b == io_state_in_12 ? 8'hf1 : _GEN_3114; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3116 = 8'h2c == io_state_in_12 ? 8'h71 : _GEN_3115; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3117 = 8'h2d == io_state_in_12 ? 8'hd8 : _GEN_3116; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3118 = 8'h2e == io_state_in_12 ? 8'h31 : _GEN_3117; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3119 = 8'h2f == io_state_in_12 ? 8'h15 : _GEN_3118; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3120 = 8'h30 == io_state_in_12 ? 8'h4 : _GEN_3119; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3121 = 8'h31 == io_state_in_12 ? 8'hc7 : _GEN_3120; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3122 = 8'h32 == io_state_in_12 ? 8'h23 : _GEN_3121; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3123 = 8'h33 == io_state_in_12 ? 8'hc3 : _GEN_3122; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3124 = 8'h34 == io_state_in_12 ? 8'h18 : _GEN_3123; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3125 = 8'h35 == io_state_in_12 ? 8'h96 : _GEN_3124; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3126 = 8'h36 == io_state_in_12 ? 8'h5 : _GEN_3125; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3127 = 8'h37 == io_state_in_12 ? 8'h9a : _GEN_3126; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3128 = 8'h38 == io_state_in_12 ? 8'h7 : _GEN_3127; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3129 = 8'h39 == io_state_in_12 ? 8'h12 : _GEN_3128; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3130 = 8'h3a == io_state_in_12 ? 8'h80 : _GEN_3129; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3131 = 8'h3b == io_state_in_12 ? 8'he2 : _GEN_3130; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3132 = 8'h3c == io_state_in_12 ? 8'heb : _GEN_3131; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3133 = 8'h3d == io_state_in_12 ? 8'h27 : _GEN_3132; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3134 = 8'h3e == io_state_in_12 ? 8'hb2 : _GEN_3133; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3135 = 8'h3f == io_state_in_12 ? 8'h75 : _GEN_3134; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3136 = 8'h40 == io_state_in_12 ? 8'h9 : _GEN_3135; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3137 = 8'h41 == io_state_in_12 ? 8'h83 : _GEN_3136; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3138 = 8'h42 == io_state_in_12 ? 8'h2c : _GEN_3137; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3139 = 8'h43 == io_state_in_12 ? 8'h1a : _GEN_3138; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3140 = 8'h44 == io_state_in_12 ? 8'h1b : _GEN_3139; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3141 = 8'h45 == io_state_in_12 ? 8'h6e : _GEN_3140; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3142 = 8'h46 == io_state_in_12 ? 8'h5a : _GEN_3141; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3143 = 8'h47 == io_state_in_12 ? 8'ha0 : _GEN_3142; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3144 = 8'h48 == io_state_in_12 ? 8'h52 : _GEN_3143; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3145 = 8'h49 == io_state_in_12 ? 8'h3b : _GEN_3144; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3146 = 8'h4a == io_state_in_12 ? 8'hd6 : _GEN_3145; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3147 = 8'h4b == io_state_in_12 ? 8'hb3 : _GEN_3146; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3148 = 8'h4c == io_state_in_12 ? 8'h29 : _GEN_3147; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3149 = 8'h4d == io_state_in_12 ? 8'he3 : _GEN_3148; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3150 = 8'h4e == io_state_in_12 ? 8'h2f : _GEN_3149; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3151 = 8'h4f == io_state_in_12 ? 8'h84 : _GEN_3150; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3152 = 8'h50 == io_state_in_12 ? 8'h53 : _GEN_3151; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3153 = 8'h51 == io_state_in_12 ? 8'hd1 : _GEN_3152; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3154 = 8'h52 == io_state_in_12 ? 8'h0 : _GEN_3153; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3155 = 8'h53 == io_state_in_12 ? 8'hed : _GEN_3154; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3156 = 8'h54 == io_state_in_12 ? 8'h20 : _GEN_3155; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3157 = 8'h55 == io_state_in_12 ? 8'hfc : _GEN_3156; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3158 = 8'h56 == io_state_in_12 ? 8'hb1 : _GEN_3157; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3159 = 8'h57 == io_state_in_12 ? 8'h5b : _GEN_3158; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3160 = 8'h58 == io_state_in_12 ? 8'h6a : _GEN_3159; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3161 = 8'h59 == io_state_in_12 ? 8'hcb : _GEN_3160; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3162 = 8'h5a == io_state_in_12 ? 8'hbe : _GEN_3161; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3163 = 8'h5b == io_state_in_12 ? 8'h39 : _GEN_3162; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3164 = 8'h5c == io_state_in_12 ? 8'h4a : _GEN_3163; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3165 = 8'h5d == io_state_in_12 ? 8'h4c : _GEN_3164; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3166 = 8'h5e == io_state_in_12 ? 8'h58 : _GEN_3165; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3167 = 8'h5f == io_state_in_12 ? 8'hcf : _GEN_3166; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3168 = 8'h60 == io_state_in_12 ? 8'hd0 : _GEN_3167; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3169 = 8'h61 == io_state_in_12 ? 8'hef : _GEN_3168; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3170 = 8'h62 == io_state_in_12 ? 8'haa : _GEN_3169; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3171 = 8'h63 == io_state_in_12 ? 8'hfb : _GEN_3170; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3172 = 8'h64 == io_state_in_12 ? 8'h43 : _GEN_3171; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3173 = 8'h65 == io_state_in_12 ? 8'h4d : _GEN_3172; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3174 = 8'h66 == io_state_in_12 ? 8'h33 : _GEN_3173; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3175 = 8'h67 == io_state_in_12 ? 8'h85 : _GEN_3174; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3176 = 8'h68 == io_state_in_12 ? 8'h45 : _GEN_3175; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3177 = 8'h69 == io_state_in_12 ? 8'hf9 : _GEN_3176; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3178 = 8'h6a == io_state_in_12 ? 8'h2 : _GEN_3177; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3179 = 8'h6b == io_state_in_12 ? 8'h7f : _GEN_3178; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3180 = 8'h6c == io_state_in_12 ? 8'h50 : _GEN_3179; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3181 = 8'h6d == io_state_in_12 ? 8'h3c : _GEN_3180; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3182 = 8'h6e == io_state_in_12 ? 8'h9f : _GEN_3181; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3183 = 8'h6f == io_state_in_12 ? 8'ha8 : _GEN_3182; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3184 = 8'h70 == io_state_in_12 ? 8'h51 : _GEN_3183; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3185 = 8'h71 == io_state_in_12 ? 8'ha3 : _GEN_3184; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3186 = 8'h72 == io_state_in_12 ? 8'h40 : _GEN_3185; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3187 = 8'h73 == io_state_in_12 ? 8'h8f : _GEN_3186; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3188 = 8'h74 == io_state_in_12 ? 8'h92 : _GEN_3187; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3189 = 8'h75 == io_state_in_12 ? 8'h9d : _GEN_3188; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3190 = 8'h76 == io_state_in_12 ? 8'h38 : _GEN_3189; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3191 = 8'h77 == io_state_in_12 ? 8'hf5 : _GEN_3190; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3192 = 8'h78 == io_state_in_12 ? 8'hbc : _GEN_3191; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3193 = 8'h79 == io_state_in_12 ? 8'hb6 : _GEN_3192; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3194 = 8'h7a == io_state_in_12 ? 8'hda : _GEN_3193; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3195 = 8'h7b == io_state_in_12 ? 8'h21 : _GEN_3194; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3196 = 8'h7c == io_state_in_12 ? 8'h10 : _GEN_3195; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3197 = 8'h7d == io_state_in_12 ? 8'hff : _GEN_3196; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3198 = 8'h7e == io_state_in_12 ? 8'hf3 : _GEN_3197; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3199 = 8'h7f == io_state_in_12 ? 8'hd2 : _GEN_3198; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3200 = 8'h80 == io_state_in_12 ? 8'hcd : _GEN_3199; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3201 = 8'h81 == io_state_in_12 ? 8'hc : _GEN_3200; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3202 = 8'h82 == io_state_in_12 ? 8'h13 : _GEN_3201; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3203 = 8'h83 == io_state_in_12 ? 8'hec : _GEN_3202; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3204 = 8'h84 == io_state_in_12 ? 8'h5f : _GEN_3203; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3205 = 8'h85 == io_state_in_12 ? 8'h97 : _GEN_3204; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3206 = 8'h86 == io_state_in_12 ? 8'h44 : _GEN_3205; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3207 = 8'h87 == io_state_in_12 ? 8'h17 : _GEN_3206; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3208 = 8'h88 == io_state_in_12 ? 8'hc4 : _GEN_3207; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3209 = 8'h89 == io_state_in_12 ? 8'ha7 : _GEN_3208; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3210 = 8'h8a == io_state_in_12 ? 8'h7e : _GEN_3209; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3211 = 8'h8b == io_state_in_12 ? 8'h3d : _GEN_3210; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3212 = 8'h8c == io_state_in_12 ? 8'h64 : _GEN_3211; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3213 = 8'h8d == io_state_in_12 ? 8'h5d : _GEN_3212; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3214 = 8'h8e == io_state_in_12 ? 8'h19 : _GEN_3213; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3215 = 8'h8f == io_state_in_12 ? 8'h73 : _GEN_3214; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3216 = 8'h90 == io_state_in_12 ? 8'h60 : _GEN_3215; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3217 = 8'h91 == io_state_in_12 ? 8'h81 : _GEN_3216; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3218 = 8'h92 == io_state_in_12 ? 8'h4f : _GEN_3217; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3219 = 8'h93 == io_state_in_12 ? 8'hdc : _GEN_3218; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3220 = 8'h94 == io_state_in_12 ? 8'h22 : _GEN_3219; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3221 = 8'h95 == io_state_in_12 ? 8'h2a : _GEN_3220; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3222 = 8'h96 == io_state_in_12 ? 8'h90 : _GEN_3221; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3223 = 8'h97 == io_state_in_12 ? 8'h88 : _GEN_3222; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3224 = 8'h98 == io_state_in_12 ? 8'h46 : _GEN_3223; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3225 = 8'h99 == io_state_in_12 ? 8'hee : _GEN_3224; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3226 = 8'h9a == io_state_in_12 ? 8'hb8 : _GEN_3225; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3227 = 8'h9b == io_state_in_12 ? 8'h14 : _GEN_3226; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3228 = 8'h9c == io_state_in_12 ? 8'hde : _GEN_3227; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3229 = 8'h9d == io_state_in_12 ? 8'h5e : _GEN_3228; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3230 = 8'h9e == io_state_in_12 ? 8'hb : _GEN_3229; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3231 = 8'h9f == io_state_in_12 ? 8'hdb : _GEN_3230; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3232 = 8'ha0 == io_state_in_12 ? 8'he0 : _GEN_3231; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3233 = 8'ha1 == io_state_in_12 ? 8'h32 : _GEN_3232; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3234 = 8'ha2 == io_state_in_12 ? 8'h3a : _GEN_3233; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3235 = 8'ha3 == io_state_in_12 ? 8'ha : _GEN_3234; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3236 = 8'ha4 == io_state_in_12 ? 8'h49 : _GEN_3235; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3237 = 8'ha5 == io_state_in_12 ? 8'h6 : _GEN_3236; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3238 = 8'ha6 == io_state_in_12 ? 8'h24 : _GEN_3237; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3239 = 8'ha7 == io_state_in_12 ? 8'h5c : _GEN_3238; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3240 = 8'ha8 == io_state_in_12 ? 8'hc2 : _GEN_3239; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3241 = 8'ha9 == io_state_in_12 ? 8'hd3 : _GEN_3240; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3242 = 8'haa == io_state_in_12 ? 8'hac : _GEN_3241; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3243 = 8'hab == io_state_in_12 ? 8'h62 : _GEN_3242; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3244 = 8'hac == io_state_in_12 ? 8'h91 : _GEN_3243; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3245 = 8'had == io_state_in_12 ? 8'h95 : _GEN_3244; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3246 = 8'hae == io_state_in_12 ? 8'he4 : _GEN_3245; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3247 = 8'haf == io_state_in_12 ? 8'h79 : _GEN_3246; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3248 = 8'hb0 == io_state_in_12 ? 8'he7 : _GEN_3247; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3249 = 8'hb1 == io_state_in_12 ? 8'hc8 : _GEN_3248; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3250 = 8'hb2 == io_state_in_12 ? 8'h37 : _GEN_3249; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3251 = 8'hb3 == io_state_in_12 ? 8'h6d : _GEN_3250; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3252 = 8'hb4 == io_state_in_12 ? 8'h8d : _GEN_3251; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3253 = 8'hb5 == io_state_in_12 ? 8'hd5 : _GEN_3252; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3254 = 8'hb6 == io_state_in_12 ? 8'h4e : _GEN_3253; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3255 = 8'hb7 == io_state_in_12 ? 8'ha9 : _GEN_3254; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3256 = 8'hb8 == io_state_in_12 ? 8'h6c : _GEN_3255; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3257 = 8'hb9 == io_state_in_12 ? 8'h56 : _GEN_3256; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3258 = 8'hba == io_state_in_12 ? 8'hf4 : _GEN_3257; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3259 = 8'hbb == io_state_in_12 ? 8'hea : _GEN_3258; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3260 = 8'hbc == io_state_in_12 ? 8'h65 : _GEN_3259; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3261 = 8'hbd == io_state_in_12 ? 8'h7a : _GEN_3260; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3262 = 8'hbe == io_state_in_12 ? 8'hae : _GEN_3261; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3263 = 8'hbf == io_state_in_12 ? 8'h8 : _GEN_3262; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3264 = 8'hc0 == io_state_in_12 ? 8'hba : _GEN_3263; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3265 = 8'hc1 == io_state_in_12 ? 8'h78 : _GEN_3264; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3266 = 8'hc2 == io_state_in_12 ? 8'h25 : _GEN_3265; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3267 = 8'hc3 == io_state_in_12 ? 8'h2e : _GEN_3266; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3268 = 8'hc4 == io_state_in_12 ? 8'h1c : _GEN_3267; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3269 = 8'hc5 == io_state_in_12 ? 8'ha6 : _GEN_3268; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3270 = 8'hc6 == io_state_in_12 ? 8'hb4 : _GEN_3269; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3271 = 8'hc7 == io_state_in_12 ? 8'hc6 : _GEN_3270; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3272 = 8'hc8 == io_state_in_12 ? 8'he8 : _GEN_3271; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3273 = 8'hc9 == io_state_in_12 ? 8'hdd : _GEN_3272; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3274 = 8'hca == io_state_in_12 ? 8'h74 : _GEN_3273; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3275 = 8'hcb == io_state_in_12 ? 8'h1f : _GEN_3274; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3276 = 8'hcc == io_state_in_12 ? 8'h4b : _GEN_3275; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3277 = 8'hcd == io_state_in_12 ? 8'hbd : _GEN_3276; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3278 = 8'hce == io_state_in_12 ? 8'h8b : _GEN_3277; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3279 = 8'hcf == io_state_in_12 ? 8'h8a : _GEN_3278; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3280 = 8'hd0 == io_state_in_12 ? 8'h70 : _GEN_3279; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3281 = 8'hd1 == io_state_in_12 ? 8'h3e : _GEN_3280; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3282 = 8'hd2 == io_state_in_12 ? 8'hb5 : _GEN_3281; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3283 = 8'hd3 == io_state_in_12 ? 8'h66 : _GEN_3282; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3284 = 8'hd4 == io_state_in_12 ? 8'h48 : _GEN_3283; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3285 = 8'hd5 == io_state_in_12 ? 8'h3 : _GEN_3284; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3286 = 8'hd6 == io_state_in_12 ? 8'hf6 : _GEN_3285; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3287 = 8'hd7 == io_state_in_12 ? 8'he : _GEN_3286; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3288 = 8'hd8 == io_state_in_12 ? 8'h61 : _GEN_3287; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3289 = 8'hd9 == io_state_in_12 ? 8'h35 : _GEN_3288; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3290 = 8'hda == io_state_in_12 ? 8'h57 : _GEN_3289; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3291 = 8'hdb == io_state_in_12 ? 8'hb9 : _GEN_3290; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3292 = 8'hdc == io_state_in_12 ? 8'h86 : _GEN_3291; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3293 = 8'hdd == io_state_in_12 ? 8'hc1 : _GEN_3292; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3294 = 8'hde == io_state_in_12 ? 8'h1d : _GEN_3293; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3295 = 8'hdf == io_state_in_12 ? 8'h9e : _GEN_3294; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3296 = 8'he0 == io_state_in_12 ? 8'he1 : _GEN_3295; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3297 = 8'he1 == io_state_in_12 ? 8'hf8 : _GEN_3296; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3298 = 8'he2 == io_state_in_12 ? 8'h98 : _GEN_3297; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3299 = 8'he3 == io_state_in_12 ? 8'h11 : _GEN_3298; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3300 = 8'he4 == io_state_in_12 ? 8'h69 : _GEN_3299; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3301 = 8'he5 == io_state_in_12 ? 8'hd9 : _GEN_3300; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3302 = 8'he6 == io_state_in_12 ? 8'h8e : _GEN_3301; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3303 = 8'he7 == io_state_in_12 ? 8'h94 : _GEN_3302; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3304 = 8'he8 == io_state_in_12 ? 8'h9b : _GEN_3303; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3305 = 8'he9 == io_state_in_12 ? 8'h1e : _GEN_3304; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3306 = 8'hea == io_state_in_12 ? 8'h87 : _GEN_3305; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3307 = 8'heb == io_state_in_12 ? 8'he9 : _GEN_3306; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3308 = 8'hec == io_state_in_12 ? 8'hce : _GEN_3307; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3309 = 8'hed == io_state_in_12 ? 8'h55 : _GEN_3308; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3310 = 8'hee == io_state_in_12 ? 8'h28 : _GEN_3309; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3311 = 8'hef == io_state_in_12 ? 8'hdf : _GEN_3310; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3312 = 8'hf0 == io_state_in_12 ? 8'h8c : _GEN_3311; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3313 = 8'hf1 == io_state_in_12 ? 8'ha1 : _GEN_3312; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3314 = 8'hf2 == io_state_in_12 ? 8'h89 : _GEN_3313; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3315 = 8'hf3 == io_state_in_12 ? 8'hd : _GEN_3314; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3316 = 8'hf4 == io_state_in_12 ? 8'hbf : _GEN_3315; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3317 = 8'hf5 == io_state_in_12 ? 8'he6 : _GEN_3316; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3318 = 8'hf6 == io_state_in_12 ? 8'h42 : _GEN_3317; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3319 = 8'hf7 == io_state_in_12 ? 8'h68 : _GEN_3318; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3320 = 8'hf8 == io_state_in_12 ? 8'h41 : _GEN_3319; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3321 = 8'hf9 == io_state_in_12 ? 8'h99 : _GEN_3320; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3322 = 8'hfa == io_state_in_12 ? 8'h2d : _GEN_3321; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3323 = 8'hfb == io_state_in_12 ? 8'hf : _GEN_3322; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3324 = 8'hfc == io_state_in_12 ? 8'hb0 : _GEN_3323; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3325 = 8'hfd == io_state_in_12 ? 8'h54 : _GEN_3324; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3326 = 8'hfe == io_state_in_12 ? 8'hbb : _GEN_3325; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3329 = 8'h1 == io_state_in_13 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3330 = 8'h2 == io_state_in_13 ? 8'h77 : _GEN_3329; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3331 = 8'h3 == io_state_in_13 ? 8'h7b : _GEN_3330; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3332 = 8'h4 == io_state_in_13 ? 8'hf2 : _GEN_3331; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3333 = 8'h5 == io_state_in_13 ? 8'h6b : _GEN_3332; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3334 = 8'h6 == io_state_in_13 ? 8'h6f : _GEN_3333; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3335 = 8'h7 == io_state_in_13 ? 8'hc5 : _GEN_3334; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3336 = 8'h8 == io_state_in_13 ? 8'h30 : _GEN_3335; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3337 = 8'h9 == io_state_in_13 ? 8'h1 : _GEN_3336; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3338 = 8'ha == io_state_in_13 ? 8'h67 : _GEN_3337; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3339 = 8'hb == io_state_in_13 ? 8'h2b : _GEN_3338; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3340 = 8'hc == io_state_in_13 ? 8'hfe : _GEN_3339; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3341 = 8'hd == io_state_in_13 ? 8'hd7 : _GEN_3340; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3342 = 8'he == io_state_in_13 ? 8'hab : _GEN_3341; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3343 = 8'hf == io_state_in_13 ? 8'h76 : _GEN_3342; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3344 = 8'h10 == io_state_in_13 ? 8'hca : _GEN_3343; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3345 = 8'h11 == io_state_in_13 ? 8'h82 : _GEN_3344; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3346 = 8'h12 == io_state_in_13 ? 8'hc9 : _GEN_3345; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3347 = 8'h13 == io_state_in_13 ? 8'h7d : _GEN_3346; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3348 = 8'h14 == io_state_in_13 ? 8'hfa : _GEN_3347; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3349 = 8'h15 == io_state_in_13 ? 8'h59 : _GEN_3348; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3350 = 8'h16 == io_state_in_13 ? 8'h47 : _GEN_3349; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3351 = 8'h17 == io_state_in_13 ? 8'hf0 : _GEN_3350; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3352 = 8'h18 == io_state_in_13 ? 8'had : _GEN_3351; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3353 = 8'h19 == io_state_in_13 ? 8'hd4 : _GEN_3352; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3354 = 8'h1a == io_state_in_13 ? 8'ha2 : _GEN_3353; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3355 = 8'h1b == io_state_in_13 ? 8'haf : _GEN_3354; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3356 = 8'h1c == io_state_in_13 ? 8'h9c : _GEN_3355; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3357 = 8'h1d == io_state_in_13 ? 8'ha4 : _GEN_3356; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3358 = 8'h1e == io_state_in_13 ? 8'h72 : _GEN_3357; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3359 = 8'h1f == io_state_in_13 ? 8'hc0 : _GEN_3358; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3360 = 8'h20 == io_state_in_13 ? 8'hb7 : _GEN_3359; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3361 = 8'h21 == io_state_in_13 ? 8'hfd : _GEN_3360; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3362 = 8'h22 == io_state_in_13 ? 8'h93 : _GEN_3361; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3363 = 8'h23 == io_state_in_13 ? 8'h26 : _GEN_3362; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3364 = 8'h24 == io_state_in_13 ? 8'h36 : _GEN_3363; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3365 = 8'h25 == io_state_in_13 ? 8'h3f : _GEN_3364; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3366 = 8'h26 == io_state_in_13 ? 8'hf7 : _GEN_3365; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3367 = 8'h27 == io_state_in_13 ? 8'hcc : _GEN_3366; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3368 = 8'h28 == io_state_in_13 ? 8'h34 : _GEN_3367; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3369 = 8'h29 == io_state_in_13 ? 8'ha5 : _GEN_3368; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3370 = 8'h2a == io_state_in_13 ? 8'he5 : _GEN_3369; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3371 = 8'h2b == io_state_in_13 ? 8'hf1 : _GEN_3370; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3372 = 8'h2c == io_state_in_13 ? 8'h71 : _GEN_3371; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3373 = 8'h2d == io_state_in_13 ? 8'hd8 : _GEN_3372; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3374 = 8'h2e == io_state_in_13 ? 8'h31 : _GEN_3373; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3375 = 8'h2f == io_state_in_13 ? 8'h15 : _GEN_3374; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3376 = 8'h30 == io_state_in_13 ? 8'h4 : _GEN_3375; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3377 = 8'h31 == io_state_in_13 ? 8'hc7 : _GEN_3376; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3378 = 8'h32 == io_state_in_13 ? 8'h23 : _GEN_3377; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3379 = 8'h33 == io_state_in_13 ? 8'hc3 : _GEN_3378; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3380 = 8'h34 == io_state_in_13 ? 8'h18 : _GEN_3379; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3381 = 8'h35 == io_state_in_13 ? 8'h96 : _GEN_3380; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3382 = 8'h36 == io_state_in_13 ? 8'h5 : _GEN_3381; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3383 = 8'h37 == io_state_in_13 ? 8'h9a : _GEN_3382; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3384 = 8'h38 == io_state_in_13 ? 8'h7 : _GEN_3383; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3385 = 8'h39 == io_state_in_13 ? 8'h12 : _GEN_3384; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3386 = 8'h3a == io_state_in_13 ? 8'h80 : _GEN_3385; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3387 = 8'h3b == io_state_in_13 ? 8'he2 : _GEN_3386; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3388 = 8'h3c == io_state_in_13 ? 8'heb : _GEN_3387; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3389 = 8'h3d == io_state_in_13 ? 8'h27 : _GEN_3388; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3390 = 8'h3e == io_state_in_13 ? 8'hb2 : _GEN_3389; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3391 = 8'h3f == io_state_in_13 ? 8'h75 : _GEN_3390; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3392 = 8'h40 == io_state_in_13 ? 8'h9 : _GEN_3391; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3393 = 8'h41 == io_state_in_13 ? 8'h83 : _GEN_3392; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3394 = 8'h42 == io_state_in_13 ? 8'h2c : _GEN_3393; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3395 = 8'h43 == io_state_in_13 ? 8'h1a : _GEN_3394; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3396 = 8'h44 == io_state_in_13 ? 8'h1b : _GEN_3395; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3397 = 8'h45 == io_state_in_13 ? 8'h6e : _GEN_3396; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3398 = 8'h46 == io_state_in_13 ? 8'h5a : _GEN_3397; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3399 = 8'h47 == io_state_in_13 ? 8'ha0 : _GEN_3398; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3400 = 8'h48 == io_state_in_13 ? 8'h52 : _GEN_3399; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3401 = 8'h49 == io_state_in_13 ? 8'h3b : _GEN_3400; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3402 = 8'h4a == io_state_in_13 ? 8'hd6 : _GEN_3401; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3403 = 8'h4b == io_state_in_13 ? 8'hb3 : _GEN_3402; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3404 = 8'h4c == io_state_in_13 ? 8'h29 : _GEN_3403; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3405 = 8'h4d == io_state_in_13 ? 8'he3 : _GEN_3404; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3406 = 8'h4e == io_state_in_13 ? 8'h2f : _GEN_3405; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3407 = 8'h4f == io_state_in_13 ? 8'h84 : _GEN_3406; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3408 = 8'h50 == io_state_in_13 ? 8'h53 : _GEN_3407; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3409 = 8'h51 == io_state_in_13 ? 8'hd1 : _GEN_3408; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3410 = 8'h52 == io_state_in_13 ? 8'h0 : _GEN_3409; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3411 = 8'h53 == io_state_in_13 ? 8'hed : _GEN_3410; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3412 = 8'h54 == io_state_in_13 ? 8'h20 : _GEN_3411; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3413 = 8'h55 == io_state_in_13 ? 8'hfc : _GEN_3412; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3414 = 8'h56 == io_state_in_13 ? 8'hb1 : _GEN_3413; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3415 = 8'h57 == io_state_in_13 ? 8'h5b : _GEN_3414; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3416 = 8'h58 == io_state_in_13 ? 8'h6a : _GEN_3415; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3417 = 8'h59 == io_state_in_13 ? 8'hcb : _GEN_3416; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3418 = 8'h5a == io_state_in_13 ? 8'hbe : _GEN_3417; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3419 = 8'h5b == io_state_in_13 ? 8'h39 : _GEN_3418; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3420 = 8'h5c == io_state_in_13 ? 8'h4a : _GEN_3419; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3421 = 8'h5d == io_state_in_13 ? 8'h4c : _GEN_3420; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3422 = 8'h5e == io_state_in_13 ? 8'h58 : _GEN_3421; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3423 = 8'h5f == io_state_in_13 ? 8'hcf : _GEN_3422; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3424 = 8'h60 == io_state_in_13 ? 8'hd0 : _GEN_3423; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3425 = 8'h61 == io_state_in_13 ? 8'hef : _GEN_3424; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3426 = 8'h62 == io_state_in_13 ? 8'haa : _GEN_3425; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3427 = 8'h63 == io_state_in_13 ? 8'hfb : _GEN_3426; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3428 = 8'h64 == io_state_in_13 ? 8'h43 : _GEN_3427; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3429 = 8'h65 == io_state_in_13 ? 8'h4d : _GEN_3428; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3430 = 8'h66 == io_state_in_13 ? 8'h33 : _GEN_3429; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3431 = 8'h67 == io_state_in_13 ? 8'h85 : _GEN_3430; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3432 = 8'h68 == io_state_in_13 ? 8'h45 : _GEN_3431; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3433 = 8'h69 == io_state_in_13 ? 8'hf9 : _GEN_3432; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3434 = 8'h6a == io_state_in_13 ? 8'h2 : _GEN_3433; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3435 = 8'h6b == io_state_in_13 ? 8'h7f : _GEN_3434; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3436 = 8'h6c == io_state_in_13 ? 8'h50 : _GEN_3435; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3437 = 8'h6d == io_state_in_13 ? 8'h3c : _GEN_3436; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3438 = 8'h6e == io_state_in_13 ? 8'h9f : _GEN_3437; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3439 = 8'h6f == io_state_in_13 ? 8'ha8 : _GEN_3438; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3440 = 8'h70 == io_state_in_13 ? 8'h51 : _GEN_3439; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3441 = 8'h71 == io_state_in_13 ? 8'ha3 : _GEN_3440; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3442 = 8'h72 == io_state_in_13 ? 8'h40 : _GEN_3441; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3443 = 8'h73 == io_state_in_13 ? 8'h8f : _GEN_3442; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3444 = 8'h74 == io_state_in_13 ? 8'h92 : _GEN_3443; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3445 = 8'h75 == io_state_in_13 ? 8'h9d : _GEN_3444; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3446 = 8'h76 == io_state_in_13 ? 8'h38 : _GEN_3445; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3447 = 8'h77 == io_state_in_13 ? 8'hf5 : _GEN_3446; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3448 = 8'h78 == io_state_in_13 ? 8'hbc : _GEN_3447; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3449 = 8'h79 == io_state_in_13 ? 8'hb6 : _GEN_3448; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3450 = 8'h7a == io_state_in_13 ? 8'hda : _GEN_3449; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3451 = 8'h7b == io_state_in_13 ? 8'h21 : _GEN_3450; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3452 = 8'h7c == io_state_in_13 ? 8'h10 : _GEN_3451; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3453 = 8'h7d == io_state_in_13 ? 8'hff : _GEN_3452; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3454 = 8'h7e == io_state_in_13 ? 8'hf3 : _GEN_3453; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3455 = 8'h7f == io_state_in_13 ? 8'hd2 : _GEN_3454; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3456 = 8'h80 == io_state_in_13 ? 8'hcd : _GEN_3455; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3457 = 8'h81 == io_state_in_13 ? 8'hc : _GEN_3456; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3458 = 8'h82 == io_state_in_13 ? 8'h13 : _GEN_3457; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3459 = 8'h83 == io_state_in_13 ? 8'hec : _GEN_3458; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3460 = 8'h84 == io_state_in_13 ? 8'h5f : _GEN_3459; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3461 = 8'h85 == io_state_in_13 ? 8'h97 : _GEN_3460; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3462 = 8'h86 == io_state_in_13 ? 8'h44 : _GEN_3461; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3463 = 8'h87 == io_state_in_13 ? 8'h17 : _GEN_3462; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3464 = 8'h88 == io_state_in_13 ? 8'hc4 : _GEN_3463; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3465 = 8'h89 == io_state_in_13 ? 8'ha7 : _GEN_3464; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3466 = 8'h8a == io_state_in_13 ? 8'h7e : _GEN_3465; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3467 = 8'h8b == io_state_in_13 ? 8'h3d : _GEN_3466; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3468 = 8'h8c == io_state_in_13 ? 8'h64 : _GEN_3467; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3469 = 8'h8d == io_state_in_13 ? 8'h5d : _GEN_3468; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3470 = 8'h8e == io_state_in_13 ? 8'h19 : _GEN_3469; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3471 = 8'h8f == io_state_in_13 ? 8'h73 : _GEN_3470; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3472 = 8'h90 == io_state_in_13 ? 8'h60 : _GEN_3471; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3473 = 8'h91 == io_state_in_13 ? 8'h81 : _GEN_3472; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3474 = 8'h92 == io_state_in_13 ? 8'h4f : _GEN_3473; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3475 = 8'h93 == io_state_in_13 ? 8'hdc : _GEN_3474; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3476 = 8'h94 == io_state_in_13 ? 8'h22 : _GEN_3475; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3477 = 8'h95 == io_state_in_13 ? 8'h2a : _GEN_3476; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3478 = 8'h96 == io_state_in_13 ? 8'h90 : _GEN_3477; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3479 = 8'h97 == io_state_in_13 ? 8'h88 : _GEN_3478; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3480 = 8'h98 == io_state_in_13 ? 8'h46 : _GEN_3479; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3481 = 8'h99 == io_state_in_13 ? 8'hee : _GEN_3480; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3482 = 8'h9a == io_state_in_13 ? 8'hb8 : _GEN_3481; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3483 = 8'h9b == io_state_in_13 ? 8'h14 : _GEN_3482; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3484 = 8'h9c == io_state_in_13 ? 8'hde : _GEN_3483; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3485 = 8'h9d == io_state_in_13 ? 8'h5e : _GEN_3484; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3486 = 8'h9e == io_state_in_13 ? 8'hb : _GEN_3485; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3487 = 8'h9f == io_state_in_13 ? 8'hdb : _GEN_3486; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3488 = 8'ha0 == io_state_in_13 ? 8'he0 : _GEN_3487; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3489 = 8'ha1 == io_state_in_13 ? 8'h32 : _GEN_3488; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3490 = 8'ha2 == io_state_in_13 ? 8'h3a : _GEN_3489; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3491 = 8'ha3 == io_state_in_13 ? 8'ha : _GEN_3490; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3492 = 8'ha4 == io_state_in_13 ? 8'h49 : _GEN_3491; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3493 = 8'ha5 == io_state_in_13 ? 8'h6 : _GEN_3492; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3494 = 8'ha6 == io_state_in_13 ? 8'h24 : _GEN_3493; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3495 = 8'ha7 == io_state_in_13 ? 8'h5c : _GEN_3494; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3496 = 8'ha8 == io_state_in_13 ? 8'hc2 : _GEN_3495; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3497 = 8'ha9 == io_state_in_13 ? 8'hd3 : _GEN_3496; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3498 = 8'haa == io_state_in_13 ? 8'hac : _GEN_3497; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3499 = 8'hab == io_state_in_13 ? 8'h62 : _GEN_3498; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3500 = 8'hac == io_state_in_13 ? 8'h91 : _GEN_3499; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3501 = 8'had == io_state_in_13 ? 8'h95 : _GEN_3500; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3502 = 8'hae == io_state_in_13 ? 8'he4 : _GEN_3501; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3503 = 8'haf == io_state_in_13 ? 8'h79 : _GEN_3502; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3504 = 8'hb0 == io_state_in_13 ? 8'he7 : _GEN_3503; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3505 = 8'hb1 == io_state_in_13 ? 8'hc8 : _GEN_3504; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3506 = 8'hb2 == io_state_in_13 ? 8'h37 : _GEN_3505; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3507 = 8'hb3 == io_state_in_13 ? 8'h6d : _GEN_3506; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3508 = 8'hb4 == io_state_in_13 ? 8'h8d : _GEN_3507; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3509 = 8'hb5 == io_state_in_13 ? 8'hd5 : _GEN_3508; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3510 = 8'hb6 == io_state_in_13 ? 8'h4e : _GEN_3509; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3511 = 8'hb7 == io_state_in_13 ? 8'ha9 : _GEN_3510; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3512 = 8'hb8 == io_state_in_13 ? 8'h6c : _GEN_3511; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3513 = 8'hb9 == io_state_in_13 ? 8'h56 : _GEN_3512; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3514 = 8'hba == io_state_in_13 ? 8'hf4 : _GEN_3513; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3515 = 8'hbb == io_state_in_13 ? 8'hea : _GEN_3514; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3516 = 8'hbc == io_state_in_13 ? 8'h65 : _GEN_3515; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3517 = 8'hbd == io_state_in_13 ? 8'h7a : _GEN_3516; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3518 = 8'hbe == io_state_in_13 ? 8'hae : _GEN_3517; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3519 = 8'hbf == io_state_in_13 ? 8'h8 : _GEN_3518; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3520 = 8'hc0 == io_state_in_13 ? 8'hba : _GEN_3519; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3521 = 8'hc1 == io_state_in_13 ? 8'h78 : _GEN_3520; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3522 = 8'hc2 == io_state_in_13 ? 8'h25 : _GEN_3521; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3523 = 8'hc3 == io_state_in_13 ? 8'h2e : _GEN_3522; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3524 = 8'hc4 == io_state_in_13 ? 8'h1c : _GEN_3523; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3525 = 8'hc5 == io_state_in_13 ? 8'ha6 : _GEN_3524; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3526 = 8'hc6 == io_state_in_13 ? 8'hb4 : _GEN_3525; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3527 = 8'hc7 == io_state_in_13 ? 8'hc6 : _GEN_3526; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3528 = 8'hc8 == io_state_in_13 ? 8'he8 : _GEN_3527; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3529 = 8'hc9 == io_state_in_13 ? 8'hdd : _GEN_3528; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3530 = 8'hca == io_state_in_13 ? 8'h74 : _GEN_3529; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3531 = 8'hcb == io_state_in_13 ? 8'h1f : _GEN_3530; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3532 = 8'hcc == io_state_in_13 ? 8'h4b : _GEN_3531; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3533 = 8'hcd == io_state_in_13 ? 8'hbd : _GEN_3532; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3534 = 8'hce == io_state_in_13 ? 8'h8b : _GEN_3533; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3535 = 8'hcf == io_state_in_13 ? 8'h8a : _GEN_3534; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3536 = 8'hd0 == io_state_in_13 ? 8'h70 : _GEN_3535; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3537 = 8'hd1 == io_state_in_13 ? 8'h3e : _GEN_3536; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3538 = 8'hd2 == io_state_in_13 ? 8'hb5 : _GEN_3537; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3539 = 8'hd3 == io_state_in_13 ? 8'h66 : _GEN_3538; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3540 = 8'hd4 == io_state_in_13 ? 8'h48 : _GEN_3539; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3541 = 8'hd5 == io_state_in_13 ? 8'h3 : _GEN_3540; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3542 = 8'hd6 == io_state_in_13 ? 8'hf6 : _GEN_3541; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3543 = 8'hd7 == io_state_in_13 ? 8'he : _GEN_3542; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3544 = 8'hd8 == io_state_in_13 ? 8'h61 : _GEN_3543; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3545 = 8'hd9 == io_state_in_13 ? 8'h35 : _GEN_3544; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3546 = 8'hda == io_state_in_13 ? 8'h57 : _GEN_3545; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3547 = 8'hdb == io_state_in_13 ? 8'hb9 : _GEN_3546; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3548 = 8'hdc == io_state_in_13 ? 8'h86 : _GEN_3547; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3549 = 8'hdd == io_state_in_13 ? 8'hc1 : _GEN_3548; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3550 = 8'hde == io_state_in_13 ? 8'h1d : _GEN_3549; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3551 = 8'hdf == io_state_in_13 ? 8'h9e : _GEN_3550; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3552 = 8'he0 == io_state_in_13 ? 8'he1 : _GEN_3551; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3553 = 8'he1 == io_state_in_13 ? 8'hf8 : _GEN_3552; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3554 = 8'he2 == io_state_in_13 ? 8'h98 : _GEN_3553; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3555 = 8'he3 == io_state_in_13 ? 8'h11 : _GEN_3554; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3556 = 8'he4 == io_state_in_13 ? 8'h69 : _GEN_3555; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3557 = 8'he5 == io_state_in_13 ? 8'hd9 : _GEN_3556; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3558 = 8'he6 == io_state_in_13 ? 8'h8e : _GEN_3557; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3559 = 8'he7 == io_state_in_13 ? 8'h94 : _GEN_3558; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3560 = 8'he8 == io_state_in_13 ? 8'h9b : _GEN_3559; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3561 = 8'he9 == io_state_in_13 ? 8'h1e : _GEN_3560; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3562 = 8'hea == io_state_in_13 ? 8'h87 : _GEN_3561; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3563 = 8'heb == io_state_in_13 ? 8'he9 : _GEN_3562; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3564 = 8'hec == io_state_in_13 ? 8'hce : _GEN_3563; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3565 = 8'hed == io_state_in_13 ? 8'h55 : _GEN_3564; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3566 = 8'hee == io_state_in_13 ? 8'h28 : _GEN_3565; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3567 = 8'hef == io_state_in_13 ? 8'hdf : _GEN_3566; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3568 = 8'hf0 == io_state_in_13 ? 8'h8c : _GEN_3567; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3569 = 8'hf1 == io_state_in_13 ? 8'ha1 : _GEN_3568; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3570 = 8'hf2 == io_state_in_13 ? 8'h89 : _GEN_3569; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3571 = 8'hf3 == io_state_in_13 ? 8'hd : _GEN_3570; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3572 = 8'hf4 == io_state_in_13 ? 8'hbf : _GEN_3571; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3573 = 8'hf5 == io_state_in_13 ? 8'he6 : _GEN_3572; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3574 = 8'hf6 == io_state_in_13 ? 8'h42 : _GEN_3573; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3575 = 8'hf7 == io_state_in_13 ? 8'h68 : _GEN_3574; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3576 = 8'hf8 == io_state_in_13 ? 8'h41 : _GEN_3575; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3577 = 8'hf9 == io_state_in_13 ? 8'h99 : _GEN_3576; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3578 = 8'hfa == io_state_in_13 ? 8'h2d : _GEN_3577; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3579 = 8'hfb == io_state_in_13 ? 8'hf : _GEN_3578; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3580 = 8'hfc == io_state_in_13 ? 8'hb0 : _GEN_3579; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3581 = 8'hfd == io_state_in_13 ? 8'h54 : _GEN_3580; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3582 = 8'hfe == io_state_in_13 ? 8'hbb : _GEN_3581; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3585 = 8'h1 == io_state_in_14 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3586 = 8'h2 == io_state_in_14 ? 8'h77 : _GEN_3585; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3587 = 8'h3 == io_state_in_14 ? 8'h7b : _GEN_3586; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3588 = 8'h4 == io_state_in_14 ? 8'hf2 : _GEN_3587; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3589 = 8'h5 == io_state_in_14 ? 8'h6b : _GEN_3588; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3590 = 8'h6 == io_state_in_14 ? 8'h6f : _GEN_3589; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3591 = 8'h7 == io_state_in_14 ? 8'hc5 : _GEN_3590; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3592 = 8'h8 == io_state_in_14 ? 8'h30 : _GEN_3591; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3593 = 8'h9 == io_state_in_14 ? 8'h1 : _GEN_3592; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3594 = 8'ha == io_state_in_14 ? 8'h67 : _GEN_3593; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3595 = 8'hb == io_state_in_14 ? 8'h2b : _GEN_3594; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3596 = 8'hc == io_state_in_14 ? 8'hfe : _GEN_3595; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3597 = 8'hd == io_state_in_14 ? 8'hd7 : _GEN_3596; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3598 = 8'he == io_state_in_14 ? 8'hab : _GEN_3597; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3599 = 8'hf == io_state_in_14 ? 8'h76 : _GEN_3598; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3600 = 8'h10 == io_state_in_14 ? 8'hca : _GEN_3599; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3601 = 8'h11 == io_state_in_14 ? 8'h82 : _GEN_3600; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3602 = 8'h12 == io_state_in_14 ? 8'hc9 : _GEN_3601; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3603 = 8'h13 == io_state_in_14 ? 8'h7d : _GEN_3602; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3604 = 8'h14 == io_state_in_14 ? 8'hfa : _GEN_3603; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3605 = 8'h15 == io_state_in_14 ? 8'h59 : _GEN_3604; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3606 = 8'h16 == io_state_in_14 ? 8'h47 : _GEN_3605; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3607 = 8'h17 == io_state_in_14 ? 8'hf0 : _GEN_3606; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3608 = 8'h18 == io_state_in_14 ? 8'had : _GEN_3607; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3609 = 8'h19 == io_state_in_14 ? 8'hd4 : _GEN_3608; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3610 = 8'h1a == io_state_in_14 ? 8'ha2 : _GEN_3609; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3611 = 8'h1b == io_state_in_14 ? 8'haf : _GEN_3610; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3612 = 8'h1c == io_state_in_14 ? 8'h9c : _GEN_3611; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3613 = 8'h1d == io_state_in_14 ? 8'ha4 : _GEN_3612; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3614 = 8'h1e == io_state_in_14 ? 8'h72 : _GEN_3613; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3615 = 8'h1f == io_state_in_14 ? 8'hc0 : _GEN_3614; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3616 = 8'h20 == io_state_in_14 ? 8'hb7 : _GEN_3615; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3617 = 8'h21 == io_state_in_14 ? 8'hfd : _GEN_3616; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3618 = 8'h22 == io_state_in_14 ? 8'h93 : _GEN_3617; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3619 = 8'h23 == io_state_in_14 ? 8'h26 : _GEN_3618; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3620 = 8'h24 == io_state_in_14 ? 8'h36 : _GEN_3619; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3621 = 8'h25 == io_state_in_14 ? 8'h3f : _GEN_3620; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3622 = 8'h26 == io_state_in_14 ? 8'hf7 : _GEN_3621; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3623 = 8'h27 == io_state_in_14 ? 8'hcc : _GEN_3622; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3624 = 8'h28 == io_state_in_14 ? 8'h34 : _GEN_3623; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3625 = 8'h29 == io_state_in_14 ? 8'ha5 : _GEN_3624; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3626 = 8'h2a == io_state_in_14 ? 8'he5 : _GEN_3625; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3627 = 8'h2b == io_state_in_14 ? 8'hf1 : _GEN_3626; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3628 = 8'h2c == io_state_in_14 ? 8'h71 : _GEN_3627; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3629 = 8'h2d == io_state_in_14 ? 8'hd8 : _GEN_3628; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3630 = 8'h2e == io_state_in_14 ? 8'h31 : _GEN_3629; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3631 = 8'h2f == io_state_in_14 ? 8'h15 : _GEN_3630; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3632 = 8'h30 == io_state_in_14 ? 8'h4 : _GEN_3631; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3633 = 8'h31 == io_state_in_14 ? 8'hc7 : _GEN_3632; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3634 = 8'h32 == io_state_in_14 ? 8'h23 : _GEN_3633; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3635 = 8'h33 == io_state_in_14 ? 8'hc3 : _GEN_3634; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3636 = 8'h34 == io_state_in_14 ? 8'h18 : _GEN_3635; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3637 = 8'h35 == io_state_in_14 ? 8'h96 : _GEN_3636; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3638 = 8'h36 == io_state_in_14 ? 8'h5 : _GEN_3637; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3639 = 8'h37 == io_state_in_14 ? 8'h9a : _GEN_3638; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3640 = 8'h38 == io_state_in_14 ? 8'h7 : _GEN_3639; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3641 = 8'h39 == io_state_in_14 ? 8'h12 : _GEN_3640; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3642 = 8'h3a == io_state_in_14 ? 8'h80 : _GEN_3641; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3643 = 8'h3b == io_state_in_14 ? 8'he2 : _GEN_3642; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3644 = 8'h3c == io_state_in_14 ? 8'heb : _GEN_3643; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3645 = 8'h3d == io_state_in_14 ? 8'h27 : _GEN_3644; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3646 = 8'h3e == io_state_in_14 ? 8'hb2 : _GEN_3645; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3647 = 8'h3f == io_state_in_14 ? 8'h75 : _GEN_3646; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3648 = 8'h40 == io_state_in_14 ? 8'h9 : _GEN_3647; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3649 = 8'h41 == io_state_in_14 ? 8'h83 : _GEN_3648; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3650 = 8'h42 == io_state_in_14 ? 8'h2c : _GEN_3649; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3651 = 8'h43 == io_state_in_14 ? 8'h1a : _GEN_3650; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3652 = 8'h44 == io_state_in_14 ? 8'h1b : _GEN_3651; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3653 = 8'h45 == io_state_in_14 ? 8'h6e : _GEN_3652; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3654 = 8'h46 == io_state_in_14 ? 8'h5a : _GEN_3653; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3655 = 8'h47 == io_state_in_14 ? 8'ha0 : _GEN_3654; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3656 = 8'h48 == io_state_in_14 ? 8'h52 : _GEN_3655; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3657 = 8'h49 == io_state_in_14 ? 8'h3b : _GEN_3656; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3658 = 8'h4a == io_state_in_14 ? 8'hd6 : _GEN_3657; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3659 = 8'h4b == io_state_in_14 ? 8'hb3 : _GEN_3658; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3660 = 8'h4c == io_state_in_14 ? 8'h29 : _GEN_3659; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3661 = 8'h4d == io_state_in_14 ? 8'he3 : _GEN_3660; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3662 = 8'h4e == io_state_in_14 ? 8'h2f : _GEN_3661; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3663 = 8'h4f == io_state_in_14 ? 8'h84 : _GEN_3662; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3664 = 8'h50 == io_state_in_14 ? 8'h53 : _GEN_3663; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3665 = 8'h51 == io_state_in_14 ? 8'hd1 : _GEN_3664; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3666 = 8'h52 == io_state_in_14 ? 8'h0 : _GEN_3665; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3667 = 8'h53 == io_state_in_14 ? 8'hed : _GEN_3666; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3668 = 8'h54 == io_state_in_14 ? 8'h20 : _GEN_3667; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3669 = 8'h55 == io_state_in_14 ? 8'hfc : _GEN_3668; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3670 = 8'h56 == io_state_in_14 ? 8'hb1 : _GEN_3669; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3671 = 8'h57 == io_state_in_14 ? 8'h5b : _GEN_3670; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3672 = 8'h58 == io_state_in_14 ? 8'h6a : _GEN_3671; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3673 = 8'h59 == io_state_in_14 ? 8'hcb : _GEN_3672; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3674 = 8'h5a == io_state_in_14 ? 8'hbe : _GEN_3673; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3675 = 8'h5b == io_state_in_14 ? 8'h39 : _GEN_3674; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3676 = 8'h5c == io_state_in_14 ? 8'h4a : _GEN_3675; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3677 = 8'h5d == io_state_in_14 ? 8'h4c : _GEN_3676; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3678 = 8'h5e == io_state_in_14 ? 8'h58 : _GEN_3677; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3679 = 8'h5f == io_state_in_14 ? 8'hcf : _GEN_3678; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3680 = 8'h60 == io_state_in_14 ? 8'hd0 : _GEN_3679; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3681 = 8'h61 == io_state_in_14 ? 8'hef : _GEN_3680; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3682 = 8'h62 == io_state_in_14 ? 8'haa : _GEN_3681; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3683 = 8'h63 == io_state_in_14 ? 8'hfb : _GEN_3682; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3684 = 8'h64 == io_state_in_14 ? 8'h43 : _GEN_3683; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3685 = 8'h65 == io_state_in_14 ? 8'h4d : _GEN_3684; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3686 = 8'h66 == io_state_in_14 ? 8'h33 : _GEN_3685; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3687 = 8'h67 == io_state_in_14 ? 8'h85 : _GEN_3686; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3688 = 8'h68 == io_state_in_14 ? 8'h45 : _GEN_3687; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3689 = 8'h69 == io_state_in_14 ? 8'hf9 : _GEN_3688; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3690 = 8'h6a == io_state_in_14 ? 8'h2 : _GEN_3689; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3691 = 8'h6b == io_state_in_14 ? 8'h7f : _GEN_3690; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3692 = 8'h6c == io_state_in_14 ? 8'h50 : _GEN_3691; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3693 = 8'h6d == io_state_in_14 ? 8'h3c : _GEN_3692; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3694 = 8'h6e == io_state_in_14 ? 8'h9f : _GEN_3693; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3695 = 8'h6f == io_state_in_14 ? 8'ha8 : _GEN_3694; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3696 = 8'h70 == io_state_in_14 ? 8'h51 : _GEN_3695; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3697 = 8'h71 == io_state_in_14 ? 8'ha3 : _GEN_3696; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3698 = 8'h72 == io_state_in_14 ? 8'h40 : _GEN_3697; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3699 = 8'h73 == io_state_in_14 ? 8'h8f : _GEN_3698; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3700 = 8'h74 == io_state_in_14 ? 8'h92 : _GEN_3699; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3701 = 8'h75 == io_state_in_14 ? 8'h9d : _GEN_3700; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3702 = 8'h76 == io_state_in_14 ? 8'h38 : _GEN_3701; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3703 = 8'h77 == io_state_in_14 ? 8'hf5 : _GEN_3702; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3704 = 8'h78 == io_state_in_14 ? 8'hbc : _GEN_3703; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3705 = 8'h79 == io_state_in_14 ? 8'hb6 : _GEN_3704; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3706 = 8'h7a == io_state_in_14 ? 8'hda : _GEN_3705; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3707 = 8'h7b == io_state_in_14 ? 8'h21 : _GEN_3706; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3708 = 8'h7c == io_state_in_14 ? 8'h10 : _GEN_3707; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3709 = 8'h7d == io_state_in_14 ? 8'hff : _GEN_3708; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3710 = 8'h7e == io_state_in_14 ? 8'hf3 : _GEN_3709; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3711 = 8'h7f == io_state_in_14 ? 8'hd2 : _GEN_3710; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3712 = 8'h80 == io_state_in_14 ? 8'hcd : _GEN_3711; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3713 = 8'h81 == io_state_in_14 ? 8'hc : _GEN_3712; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3714 = 8'h82 == io_state_in_14 ? 8'h13 : _GEN_3713; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3715 = 8'h83 == io_state_in_14 ? 8'hec : _GEN_3714; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3716 = 8'h84 == io_state_in_14 ? 8'h5f : _GEN_3715; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3717 = 8'h85 == io_state_in_14 ? 8'h97 : _GEN_3716; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3718 = 8'h86 == io_state_in_14 ? 8'h44 : _GEN_3717; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3719 = 8'h87 == io_state_in_14 ? 8'h17 : _GEN_3718; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3720 = 8'h88 == io_state_in_14 ? 8'hc4 : _GEN_3719; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3721 = 8'h89 == io_state_in_14 ? 8'ha7 : _GEN_3720; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3722 = 8'h8a == io_state_in_14 ? 8'h7e : _GEN_3721; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3723 = 8'h8b == io_state_in_14 ? 8'h3d : _GEN_3722; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3724 = 8'h8c == io_state_in_14 ? 8'h64 : _GEN_3723; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3725 = 8'h8d == io_state_in_14 ? 8'h5d : _GEN_3724; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3726 = 8'h8e == io_state_in_14 ? 8'h19 : _GEN_3725; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3727 = 8'h8f == io_state_in_14 ? 8'h73 : _GEN_3726; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3728 = 8'h90 == io_state_in_14 ? 8'h60 : _GEN_3727; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3729 = 8'h91 == io_state_in_14 ? 8'h81 : _GEN_3728; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3730 = 8'h92 == io_state_in_14 ? 8'h4f : _GEN_3729; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3731 = 8'h93 == io_state_in_14 ? 8'hdc : _GEN_3730; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3732 = 8'h94 == io_state_in_14 ? 8'h22 : _GEN_3731; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3733 = 8'h95 == io_state_in_14 ? 8'h2a : _GEN_3732; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3734 = 8'h96 == io_state_in_14 ? 8'h90 : _GEN_3733; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3735 = 8'h97 == io_state_in_14 ? 8'h88 : _GEN_3734; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3736 = 8'h98 == io_state_in_14 ? 8'h46 : _GEN_3735; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3737 = 8'h99 == io_state_in_14 ? 8'hee : _GEN_3736; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3738 = 8'h9a == io_state_in_14 ? 8'hb8 : _GEN_3737; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3739 = 8'h9b == io_state_in_14 ? 8'h14 : _GEN_3738; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3740 = 8'h9c == io_state_in_14 ? 8'hde : _GEN_3739; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3741 = 8'h9d == io_state_in_14 ? 8'h5e : _GEN_3740; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3742 = 8'h9e == io_state_in_14 ? 8'hb : _GEN_3741; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3743 = 8'h9f == io_state_in_14 ? 8'hdb : _GEN_3742; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3744 = 8'ha0 == io_state_in_14 ? 8'he0 : _GEN_3743; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3745 = 8'ha1 == io_state_in_14 ? 8'h32 : _GEN_3744; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3746 = 8'ha2 == io_state_in_14 ? 8'h3a : _GEN_3745; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3747 = 8'ha3 == io_state_in_14 ? 8'ha : _GEN_3746; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3748 = 8'ha4 == io_state_in_14 ? 8'h49 : _GEN_3747; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3749 = 8'ha5 == io_state_in_14 ? 8'h6 : _GEN_3748; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3750 = 8'ha6 == io_state_in_14 ? 8'h24 : _GEN_3749; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3751 = 8'ha7 == io_state_in_14 ? 8'h5c : _GEN_3750; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3752 = 8'ha8 == io_state_in_14 ? 8'hc2 : _GEN_3751; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3753 = 8'ha9 == io_state_in_14 ? 8'hd3 : _GEN_3752; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3754 = 8'haa == io_state_in_14 ? 8'hac : _GEN_3753; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3755 = 8'hab == io_state_in_14 ? 8'h62 : _GEN_3754; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3756 = 8'hac == io_state_in_14 ? 8'h91 : _GEN_3755; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3757 = 8'had == io_state_in_14 ? 8'h95 : _GEN_3756; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3758 = 8'hae == io_state_in_14 ? 8'he4 : _GEN_3757; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3759 = 8'haf == io_state_in_14 ? 8'h79 : _GEN_3758; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3760 = 8'hb0 == io_state_in_14 ? 8'he7 : _GEN_3759; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3761 = 8'hb1 == io_state_in_14 ? 8'hc8 : _GEN_3760; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3762 = 8'hb2 == io_state_in_14 ? 8'h37 : _GEN_3761; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3763 = 8'hb3 == io_state_in_14 ? 8'h6d : _GEN_3762; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3764 = 8'hb4 == io_state_in_14 ? 8'h8d : _GEN_3763; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3765 = 8'hb5 == io_state_in_14 ? 8'hd5 : _GEN_3764; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3766 = 8'hb6 == io_state_in_14 ? 8'h4e : _GEN_3765; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3767 = 8'hb7 == io_state_in_14 ? 8'ha9 : _GEN_3766; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3768 = 8'hb8 == io_state_in_14 ? 8'h6c : _GEN_3767; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3769 = 8'hb9 == io_state_in_14 ? 8'h56 : _GEN_3768; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3770 = 8'hba == io_state_in_14 ? 8'hf4 : _GEN_3769; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3771 = 8'hbb == io_state_in_14 ? 8'hea : _GEN_3770; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3772 = 8'hbc == io_state_in_14 ? 8'h65 : _GEN_3771; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3773 = 8'hbd == io_state_in_14 ? 8'h7a : _GEN_3772; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3774 = 8'hbe == io_state_in_14 ? 8'hae : _GEN_3773; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3775 = 8'hbf == io_state_in_14 ? 8'h8 : _GEN_3774; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3776 = 8'hc0 == io_state_in_14 ? 8'hba : _GEN_3775; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3777 = 8'hc1 == io_state_in_14 ? 8'h78 : _GEN_3776; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3778 = 8'hc2 == io_state_in_14 ? 8'h25 : _GEN_3777; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3779 = 8'hc3 == io_state_in_14 ? 8'h2e : _GEN_3778; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3780 = 8'hc4 == io_state_in_14 ? 8'h1c : _GEN_3779; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3781 = 8'hc5 == io_state_in_14 ? 8'ha6 : _GEN_3780; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3782 = 8'hc6 == io_state_in_14 ? 8'hb4 : _GEN_3781; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3783 = 8'hc7 == io_state_in_14 ? 8'hc6 : _GEN_3782; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3784 = 8'hc8 == io_state_in_14 ? 8'he8 : _GEN_3783; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3785 = 8'hc9 == io_state_in_14 ? 8'hdd : _GEN_3784; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3786 = 8'hca == io_state_in_14 ? 8'h74 : _GEN_3785; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3787 = 8'hcb == io_state_in_14 ? 8'h1f : _GEN_3786; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3788 = 8'hcc == io_state_in_14 ? 8'h4b : _GEN_3787; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3789 = 8'hcd == io_state_in_14 ? 8'hbd : _GEN_3788; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3790 = 8'hce == io_state_in_14 ? 8'h8b : _GEN_3789; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3791 = 8'hcf == io_state_in_14 ? 8'h8a : _GEN_3790; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3792 = 8'hd0 == io_state_in_14 ? 8'h70 : _GEN_3791; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3793 = 8'hd1 == io_state_in_14 ? 8'h3e : _GEN_3792; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3794 = 8'hd2 == io_state_in_14 ? 8'hb5 : _GEN_3793; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3795 = 8'hd3 == io_state_in_14 ? 8'h66 : _GEN_3794; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3796 = 8'hd4 == io_state_in_14 ? 8'h48 : _GEN_3795; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3797 = 8'hd5 == io_state_in_14 ? 8'h3 : _GEN_3796; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3798 = 8'hd6 == io_state_in_14 ? 8'hf6 : _GEN_3797; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3799 = 8'hd7 == io_state_in_14 ? 8'he : _GEN_3798; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3800 = 8'hd8 == io_state_in_14 ? 8'h61 : _GEN_3799; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3801 = 8'hd9 == io_state_in_14 ? 8'h35 : _GEN_3800; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3802 = 8'hda == io_state_in_14 ? 8'h57 : _GEN_3801; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3803 = 8'hdb == io_state_in_14 ? 8'hb9 : _GEN_3802; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3804 = 8'hdc == io_state_in_14 ? 8'h86 : _GEN_3803; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3805 = 8'hdd == io_state_in_14 ? 8'hc1 : _GEN_3804; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3806 = 8'hde == io_state_in_14 ? 8'h1d : _GEN_3805; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3807 = 8'hdf == io_state_in_14 ? 8'h9e : _GEN_3806; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3808 = 8'he0 == io_state_in_14 ? 8'he1 : _GEN_3807; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3809 = 8'he1 == io_state_in_14 ? 8'hf8 : _GEN_3808; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3810 = 8'he2 == io_state_in_14 ? 8'h98 : _GEN_3809; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3811 = 8'he3 == io_state_in_14 ? 8'h11 : _GEN_3810; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3812 = 8'he4 == io_state_in_14 ? 8'h69 : _GEN_3811; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3813 = 8'he5 == io_state_in_14 ? 8'hd9 : _GEN_3812; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3814 = 8'he6 == io_state_in_14 ? 8'h8e : _GEN_3813; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3815 = 8'he7 == io_state_in_14 ? 8'h94 : _GEN_3814; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3816 = 8'he8 == io_state_in_14 ? 8'h9b : _GEN_3815; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3817 = 8'he9 == io_state_in_14 ? 8'h1e : _GEN_3816; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3818 = 8'hea == io_state_in_14 ? 8'h87 : _GEN_3817; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3819 = 8'heb == io_state_in_14 ? 8'he9 : _GEN_3818; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3820 = 8'hec == io_state_in_14 ? 8'hce : _GEN_3819; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3821 = 8'hed == io_state_in_14 ? 8'h55 : _GEN_3820; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3822 = 8'hee == io_state_in_14 ? 8'h28 : _GEN_3821; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3823 = 8'hef == io_state_in_14 ? 8'hdf : _GEN_3822; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3824 = 8'hf0 == io_state_in_14 ? 8'h8c : _GEN_3823; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3825 = 8'hf1 == io_state_in_14 ? 8'ha1 : _GEN_3824; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3826 = 8'hf2 == io_state_in_14 ? 8'h89 : _GEN_3825; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3827 = 8'hf3 == io_state_in_14 ? 8'hd : _GEN_3826; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3828 = 8'hf4 == io_state_in_14 ? 8'hbf : _GEN_3827; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3829 = 8'hf5 == io_state_in_14 ? 8'he6 : _GEN_3828; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3830 = 8'hf6 == io_state_in_14 ? 8'h42 : _GEN_3829; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3831 = 8'hf7 == io_state_in_14 ? 8'h68 : _GEN_3830; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3832 = 8'hf8 == io_state_in_14 ? 8'h41 : _GEN_3831; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3833 = 8'hf9 == io_state_in_14 ? 8'h99 : _GEN_3832; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3834 = 8'hfa == io_state_in_14 ? 8'h2d : _GEN_3833; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3835 = 8'hfb == io_state_in_14 ? 8'hf : _GEN_3834; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3836 = 8'hfc == io_state_in_14 ? 8'hb0 : _GEN_3835; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3837 = 8'hfd == io_state_in_14 ? 8'h54 : _GEN_3836; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3838 = 8'hfe == io_state_in_14 ? 8'hbb : _GEN_3837; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3841 = 8'h1 == io_state_in_15 ? 8'h7c : 8'h63; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3842 = 8'h2 == io_state_in_15 ? 8'h77 : _GEN_3841; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3843 = 8'h3 == io_state_in_15 ? 8'h7b : _GEN_3842; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3844 = 8'h4 == io_state_in_15 ? 8'hf2 : _GEN_3843; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3845 = 8'h5 == io_state_in_15 ? 8'h6b : _GEN_3844; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3846 = 8'h6 == io_state_in_15 ? 8'h6f : _GEN_3845; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3847 = 8'h7 == io_state_in_15 ? 8'hc5 : _GEN_3846; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3848 = 8'h8 == io_state_in_15 ? 8'h30 : _GEN_3847; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3849 = 8'h9 == io_state_in_15 ? 8'h1 : _GEN_3848; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3850 = 8'ha == io_state_in_15 ? 8'h67 : _GEN_3849; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3851 = 8'hb == io_state_in_15 ? 8'h2b : _GEN_3850; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3852 = 8'hc == io_state_in_15 ? 8'hfe : _GEN_3851; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3853 = 8'hd == io_state_in_15 ? 8'hd7 : _GEN_3852; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3854 = 8'he == io_state_in_15 ? 8'hab : _GEN_3853; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3855 = 8'hf == io_state_in_15 ? 8'h76 : _GEN_3854; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3856 = 8'h10 == io_state_in_15 ? 8'hca : _GEN_3855; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3857 = 8'h11 == io_state_in_15 ? 8'h82 : _GEN_3856; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3858 = 8'h12 == io_state_in_15 ? 8'hc9 : _GEN_3857; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3859 = 8'h13 == io_state_in_15 ? 8'h7d : _GEN_3858; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3860 = 8'h14 == io_state_in_15 ? 8'hfa : _GEN_3859; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3861 = 8'h15 == io_state_in_15 ? 8'h59 : _GEN_3860; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3862 = 8'h16 == io_state_in_15 ? 8'h47 : _GEN_3861; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3863 = 8'h17 == io_state_in_15 ? 8'hf0 : _GEN_3862; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3864 = 8'h18 == io_state_in_15 ? 8'had : _GEN_3863; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3865 = 8'h19 == io_state_in_15 ? 8'hd4 : _GEN_3864; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3866 = 8'h1a == io_state_in_15 ? 8'ha2 : _GEN_3865; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3867 = 8'h1b == io_state_in_15 ? 8'haf : _GEN_3866; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3868 = 8'h1c == io_state_in_15 ? 8'h9c : _GEN_3867; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3869 = 8'h1d == io_state_in_15 ? 8'ha4 : _GEN_3868; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3870 = 8'h1e == io_state_in_15 ? 8'h72 : _GEN_3869; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3871 = 8'h1f == io_state_in_15 ? 8'hc0 : _GEN_3870; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3872 = 8'h20 == io_state_in_15 ? 8'hb7 : _GEN_3871; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3873 = 8'h21 == io_state_in_15 ? 8'hfd : _GEN_3872; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3874 = 8'h22 == io_state_in_15 ? 8'h93 : _GEN_3873; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3875 = 8'h23 == io_state_in_15 ? 8'h26 : _GEN_3874; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3876 = 8'h24 == io_state_in_15 ? 8'h36 : _GEN_3875; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3877 = 8'h25 == io_state_in_15 ? 8'h3f : _GEN_3876; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3878 = 8'h26 == io_state_in_15 ? 8'hf7 : _GEN_3877; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3879 = 8'h27 == io_state_in_15 ? 8'hcc : _GEN_3878; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3880 = 8'h28 == io_state_in_15 ? 8'h34 : _GEN_3879; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3881 = 8'h29 == io_state_in_15 ? 8'ha5 : _GEN_3880; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3882 = 8'h2a == io_state_in_15 ? 8'he5 : _GEN_3881; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3883 = 8'h2b == io_state_in_15 ? 8'hf1 : _GEN_3882; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3884 = 8'h2c == io_state_in_15 ? 8'h71 : _GEN_3883; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3885 = 8'h2d == io_state_in_15 ? 8'hd8 : _GEN_3884; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3886 = 8'h2e == io_state_in_15 ? 8'h31 : _GEN_3885; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3887 = 8'h2f == io_state_in_15 ? 8'h15 : _GEN_3886; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3888 = 8'h30 == io_state_in_15 ? 8'h4 : _GEN_3887; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3889 = 8'h31 == io_state_in_15 ? 8'hc7 : _GEN_3888; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3890 = 8'h32 == io_state_in_15 ? 8'h23 : _GEN_3889; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3891 = 8'h33 == io_state_in_15 ? 8'hc3 : _GEN_3890; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3892 = 8'h34 == io_state_in_15 ? 8'h18 : _GEN_3891; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3893 = 8'h35 == io_state_in_15 ? 8'h96 : _GEN_3892; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3894 = 8'h36 == io_state_in_15 ? 8'h5 : _GEN_3893; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3895 = 8'h37 == io_state_in_15 ? 8'h9a : _GEN_3894; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3896 = 8'h38 == io_state_in_15 ? 8'h7 : _GEN_3895; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3897 = 8'h39 == io_state_in_15 ? 8'h12 : _GEN_3896; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3898 = 8'h3a == io_state_in_15 ? 8'h80 : _GEN_3897; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3899 = 8'h3b == io_state_in_15 ? 8'he2 : _GEN_3898; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3900 = 8'h3c == io_state_in_15 ? 8'heb : _GEN_3899; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3901 = 8'h3d == io_state_in_15 ? 8'h27 : _GEN_3900; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3902 = 8'h3e == io_state_in_15 ? 8'hb2 : _GEN_3901; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3903 = 8'h3f == io_state_in_15 ? 8'h75 : _GEN_3902; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3904 = 8'h40 == io_state_in_15 ? 8'h9 : _GEN_3903; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3905 = 8'h41 == io_state_in_15 ? 8'h83 : _GEN_3904; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3906 = 8'h42 == io_state_in_15 ? 8'h2c : _GEN_3905; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3907 = 8'h43 == io_state_in_15 ? 8'h1a : _GEN_3906; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3908 = 8'h44 == io_state_in_15 ? 8'h1b : _GEN_3907; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3909 = 8'h45 == io_state_in_15 ? 8'h6e : _GEN_3908; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3910 = 8'h46 == io_state_in_15 ? 8'h5a : _GEN_3909; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3911 = 8'h47 == io_state_in_15 ? 8'ha0 : _GEN_3910; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3912 = 8'h48 == io_state_in_15 ? 8'h52 : _GEN_3911; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3913 = 8'h49 == io_state_in_15 ? 8'h3b : _GEN_3912; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3914 = 8'h4a == io_state_in_15 ? 8'hd6 : _GEN_3913; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3915 = 8'h4b == io_state_in_15 ? 8'hb3 : _GEN_3914; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3916 = 8'h4c == io_state_in_15 ? 8'h29 : _GEN_3915; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3917 = 8'h4d == io_state_in_15 ? 8'he3 : _GEN_3916; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3918 = 8'h4e == io_state_in_15 ? 8'h2f : _GEN_3917; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3919 = 8'h4f == io_state_in_15 ? 8'h84 : _GEN_3918; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3920 = 8'h50 == io_state_in_15 ? 8'h53 : _GEN_3919; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3921 = 8'h51 == io_state_in_15 ? 8'hd1 : _GEN_3920; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3922 = 8'h52 == io_state_in_15 ? 8'h0 : _GEN_3921; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3923 = 8'h53 == io_state_in_15 ? 8'hed : _GEN_3922; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3924 = 8'h54 == io_state_in_15 ? 8'h20 : _GEN_3923; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3925 = 8'h55 == io_state_in_15 ? 8'hfc : _GEN_3924; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3926 = 8'h56 == io_state_in_15 ? 8'hb1 : _GEN_3925; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3927 = 8'h57 == io_state_in_15 ? 8'h5b : _GEN_3926; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3928 = 8'h58 == io_state_in_15 ? 8'h6a : _GEN_3927; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3929 = 8'h59 == io_state_in_15 ? 8'hcb : _GEN_3928; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3930 = 8'h5a == io_state_in_15 ? 8'hbe : _GEN_3929; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3931 = 8'h5b == io_state_in_15 ? 8'h39 : _GEN_3930; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3932 = 8'h5c == io_state_in_15 ? 8'h4a : _GEN_3931; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3933 = 8'h5d == io_state_in_15 ? 8'h4c : _GEN_3932; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3934 = 8'h5e == io_state_in_15 ? 8'h58 : _GEN_3933; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3935 = 8'h5f == io_state_in_15 ? 8'hcf : _GEN_3934; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3936 = 8'h60 == io_state_in_15 ? 8'hd0 : _GEN_3935; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3937 = 8'h61 == io_state_in_15 ? 8'hef : _GEN_3936; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3938 = 8'h62 == io_state_in_15 ? 8'haa : _GEN_3937; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3939 = 8'h63 == io_state_in_15 ? 8'hfb : _GEN_3938; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3940 = 8'h64 == io_state_in_15 ? 8'h43 : _GEN_3939; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3941 = 8'h65 == io_state_in_15 ? 8'h4d : _GEN_3940; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3942 = 8'h66 == io_state_in_15 ? 8'h33 : _GEN_3941; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3943 = 8'h67 == io_state_in_15 ? 8'h85 : _GEN_3942; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3944 = 8'h68 == io_state_in_15 ? 8'h45 : _GEN_3943; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3945 = 8'h69 == io_state_in_15 ? 8'hf9 : _GEN_3944; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3946 = 8'h6a == io_state_in_15 ? 8'h2 : _GEN_3945; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3947 = 8'h6b == io_state_in_15 ? 8'h7f : _GEN_3946; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3948 = 8'h6c == io_state_in_15 ? 8'h50 : _GEN_3947; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3949 = 8'h6d == io_state_in_15 ? 8'h3c : _GEN_3948; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3950 = 8'h6e == io_state_in_15 ? 8'h9f : _GEN_3949; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3951 = 8'h6f == io_state_in_15 ? 8'ha8 : _GEN_3950; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3952 = 8'h70 == io_state_in_15 ? 8'h51 : _GEN_3951; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3953 = 8'h71 == io_state_in_15 ? 8'ha3 : _GEN_3952; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3954 = 8'h72 == io_state_in_15 ? 8'h40 : _GEN_3953; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3955 = 8'h73 == io_state_in_15 ? 8'h8f : _GEN_3954; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3956 = 8'h74 == io_state_in_15 ? 8'h92 : _GEN_3955; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3957 = 8'h75 == io_state_in_15 ? 8'h9d : _GEN_3956; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3958 = 8'h76 == io_state_in_15 ? 8'h38 : _GEN_3957; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3959 = 8'h77 == io_state_in_15 ? 8'hf5 : _GEN_3958; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3960 = 8'h78 == io_state_in_15 ? 8'hbc : _GEN_3959; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3961 = 8'h79 == io_state_in_15 ? 8'hb6 : _GEN_3960; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3962 = 8'h7a == io_state_in_15 ? 8'hda : _GEN_3961; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3963 = 8'h7b == io_state_in_15 ? 8'h21 : _GEN_3962; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3964 = 8'h7c == io_state_in_15 ? 8'h10 : _GEN_3963; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3965 = 8'h7d == io_state_in_15 ? 8'hff : _GEN_3964; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3966 = 8'h7e == io_state_in_15 ? 8'hf3 : _GEN_3965; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3967 = 8'h7f == io_state_in_15 ? 8'hd2 : _GEN_3966; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3968 = 8'h80 == io_state_in_15 ? 8'hcd : _GEN_3967; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3969 = 8'h81 == io_state_in_15 ? 8'hc : _GEN_3968; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3970 = 8'h82 == io_state_in_15 ? 8'h13 : _GEN_3969; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3971 = 8'h83 == io_state_in_15 ? 8'hec : _GEN_3970; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3972 = 8'h84 == io_state_in_15 ? 8'h5f : _GEN_3971; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3973 = 8'h85 == io_state_in_15 ? 8'h97 : _GEN_3972; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3974 = 8'h86 == io_state_in_15 ? 8'h44 : _GEN_3973; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3975 = 8'h87 == io_state_in_15 ? 8'h17 : _GEN_3974; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3976 = 8'h88 == io_state_in_15 ? 8'hc4 : _GEN_3975; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3977 = 8'h89 == io_state_in_15 ? 8'ha7 : _GEN_3976; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3978 = 8'h8a == io_state_in_15 ? 8'h7e : _GEN_3977; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3979 = 8'h8b == io_state_in_15 ? 8'h3d : _GEN_3978; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3980 = 8'h8c == io_state_in_15 ? 8'h64 : _GEN_3979; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3981 = 8'h8d == io_state_in_15 ? 8'h5d : _GEN_3980; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3982 = 8'h8e == io_state_in_15 ? 8'h19 : _GEN_3981; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3983 = 8'h8f == io_state_in_15 ? 8'h73 : _GEN_3982; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3984 = 8'h90 == io_state_in_15 ? 8'h60 : _GEN_3983; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3985 = 8'h91 == io_state_in_15 ? 8'h81 : _GEN_3984; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3986 = 8'h92 == io_state_in_15 ? 8'h4f : _GEN_3985; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3987 = 8'h93 == io_state_in_15 ? 8'hdc : _GEN_3986; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3988 = 8'h94 == io_state_in_15 ? 8'h22 : _GEN_3987; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3989 = 8'h95 == io_state_in_15 ? 8'h2a : _GEN_3988; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3990 = 8'h96 == io_state_in_15 ? 8'h90 : _GEN_3989; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3991 = 8'h97 == io_state_in_15 ? 8'h88 : _GEN_3990; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3992 = 8'h98 == io_state_in_15 ? 8'h46 : _GEN_3991; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3993 = 8'h99 == io_state_in_15 ? 8'hee : _GEN_3992; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3994 = 8'h9a == io_state_in_15 ? 8'hb8 : _GEN_3993; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3995 = 8'h9b == io_state_in_15 ? 8'h14 : _GEN_3994; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3996 = 8'h9c == io_state_in_15 ? 8'hde : _GEN_3995; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3997 = 8'h9d == io_state_in_15 ? 8'h5e : _GEN_3996; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3998 = 8'h9e == io_state_in_15 ? 8'hb : _GEN_3997; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_3999 = 8'h9f == io_state_in_15 ? 8'hdb : _GEN_3998; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4000 = 8'ha0 == io_state_in_15 ? 8'he0 : _GEN_3999; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4001 = 8'ha1 == io_state_in_15 ? 8'h32 : _GEN_4000; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4002 = 8'ha2 == io_state_in_15 ? 8'h3a : _GEN_4001; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4003 = 8'ha3 == io_state_in_15 ? 8'ha : _GEN_4002; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4004 = 8'ha4 == io_state_in_15 ? 8'h49 : _GEN_4003; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4005 = 8'ha5 == io_state_in_15 ? 8'h6 : _GEN_4004; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4006 = 8'ha6 == io_state_in_15 ? 8'h24 : _GEN_4005; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4007 = 8'ha7 == io_state_in_15 ? 8'h5c : _GEN_4006; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4008 = 8'ha8 == io_state_in_15 ? 8'hc2 : _GEN_4007; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4009 = 8'ha9 == io_state_in_15 ? 8'hd3 : _GEN_4008; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4010 = 8'haa == io_state_in_15 ? 8'hac : _GEN_4009; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4011 = 8'hab == io_state_in_15 ? 8'h62 : _GEN_4010; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4012 = 8'hac == io_state_in_15 ? 8'h91 : _GEN_4011; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4013 = 8'had == io_state_in_15 ? 8'h95 : _GEN_4012; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4014 = 8'hae == io_state_in_15 ? 8'he4 : _GEN_4013; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4015 = 8'haf == io_state_in_15 ? 8'h79 : _GEN_4014; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4016 = 8'hb0 == io_state_in_15 ? 8'he7 : _GEN_4015; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4017 = 8'hb1 == io_state_in_15 ? 8'hc8 : _GEN_4016; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4018 = 8'hb2 == io_state_in_15 ? 8'h37 : _GEN_4017; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4019 = 8'hb3 == io_state_in_15 ? 8'h6d : _GEN_4018; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4020 = 8'hb4 == io_state_in_15 ? 8'h8d : _GEN_4019; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4021 = 8'hb5 == io_state_in_15 ? 8'hd5 : _GEN_4020; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4022 = 8'hb6 == io_state_in_15 ? 8'h4e : _GEN_4021; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4023 = 8'hb7 == io_state_in_15 ? 8'ha9 : _GEN_4022; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4024 = 8'hb8 == io_state_in_15 ? 8'h6c : _GEN_4023; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4025 = 8'hb9 == io_state_in_15 ? 8'h56 : _GEN_4024; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4026 = 8'hba == io_state_in_15 ? 8'hf4 : _GEN_4025; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4027 = 8'hbb == io_state_in_15 ? 8'hea : _GEN_4026; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4028 = 8'hbc == io_state_in_15 ? 8'h65 : _GEN_4027; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4029 = 8'hbd == io_state_in_15 ? 8'h7a : _GEN_4028; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4030 = 8'hbe == io_state_in_15 ? 8'hae : _GEN_4029; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4031 = 8'hbf == io_state_in_15 ? 8'h8 : _GEN_4030; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4032 = 8'hc0 == io_state_in_15 ? 8'hba : _GEN_4031; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4033 = 8'hc1 == io_state_in_15 ? 8'h78 : _GEN_4032; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4034 = 8'hc2 == io_state_in_15 ? 8'h25 : _GEN_4033; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4035 = 8'hc3 == io_state_in_15 ? 8'h2e : _GEN_4034; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4036 = 8'hc4 == io_state_in_15 ? 8'h1c : _GEN_4035; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4037 = 8'hc5 == io_state_in_15 ? 8'ha6 : _GEN_4036; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4038 = 8'hc6 == io_state_in_15 ? 8'hb4 : _GEN_4037; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4039 = 8'hc7 == io_state_in_15 ? 8'hc6 : _GEN_4038; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4040 = 8'hc8 == io_state_in_15 ? 8'he8 : _GEN_4039; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4041 = 8'hc9 == io_state_in_15 ? 8'hdd : _GEN_4040; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4042 = 8'hca == io_state_in_15 ? 8'h74 : _GEN_4041; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4043 = 8'hcb == io_state_in_15 ? 8'h1f : _GEN_4042; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4044 = 8'hcc == io_state_in_15 ? 8'h4b : _GEN_4043; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4045 = 8'hcd == io_state_in_15 ? 8'hbd : _GEN_4044; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4046 = 8'hce == io_state_in_15 ? 8'h8b : _GEN_4045; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4047 = 8'hcf == io_state_in_15 ? 8'h8a : _GEN_4046; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4048 = 8'hd0 == io_state_in_15 ? 8'h70 : _GEN_4047; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4049 = 8'hd1 == io_state_in_15 ? 8'h3e : _GEN_4048; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4050 = 8'hd2 == io_state_in_15 ? 8'hb5 : _GEN_4049; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4051 = 8'hd3 == io_state_in_15 ? 8'h66 : _GEN_4050; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4052 = 8'hd4 == io_state_in_15 ? 8'h48 : _GEN_4051; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4053 = 8'hd5 == io_state_in_15 ? 8'h3 : _GEN_4052; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4054 = 8'hd6 == io_state_in_15 ? 8'hf6 : _GEN_4053; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4055 = 8'hd7 == io_state_in_15 ? 8'he : _GEN_4054; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4056 = 8'hd8 == io_state_in_15 ? 8'h61 : _GEN_4055; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4057 = 8'hd9 == io_state_in_15 ? 8'h35 : _GEN_4056; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4058 = 8'hda == io_state_in_15 ? 8'h57 : _GEN_4057; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4059 = 8'hdb == io_state_in_15 ? 8'hb9 : _GEN_4058; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4060 = 8'hdc == io_state_in_15 ? 8'h86 : _GEN_4059; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4061 = 8'hdd == io_state_in_15 ? 8'hc1 : _GEN_4060; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4062 = 8'hde == io_state_in_15 ? 8'h1d : _GEN_4061; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4063 = 8'hdf == io_state_in_15 ? 8'h9e : _GEN_4062; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4064 = 8'he0 == io_state_in_15 ? 8'he1 : _GEN_4063; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4065 = 8'he1 == io_state_in_15 ? 8'hf8 : _GEN_4064; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4066 = 8'he2 == io_state_in_15 ? 8'h98 : _GEN_4065; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4067 = 8'he3 == io_state_in_15 ? 8'h11 : _GEN_4066; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4068 = 8'he4 == io_state_in_15 ? 8'h69 : _GEN_4067; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4069 = 8'he5 == io_state_in_15 ? 8'hd9 : _GEN_4068; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4070 = 8'he6 == io_state_in_15 ? 8'h8e : _GEN_4069; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4071 = 8'he7 == io_state_in_15 ? 8'h94 : _GEN_4070; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4072 = 8'he8 == io_state_in_15 ? 8'h9b : _GEN_4071; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4073 = 8'he9 == io_state_in_15 ? 8'h1e : _GEN_4072; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4074 = 8'hea == io_state_in_15 ? 8'h87 : _GEN_4073; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4075 = 8'heb == io_state_in_15 ? 8'he9 : _GEN_4074; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4076 = 8'hec == io_state_in_15 ? 8'hce : _GEN_4075; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4077 = 8'hed == io_state_in_15 ? 8'h55 : _GEN_4076; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4078 = 8'hee == io_state_in_15 ? 8'h28 : _GEN_4077; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4079 = 8'hef == io_state_in_15 ? 8'hdf : _GEN_4078; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4080 = 8'hf0 == io_state_in_15 ? 8'h8c : _GEN_4079; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4081 = 8'hf1 == io_state_in_15 ? 8'ha1 : _GEN_4080; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4082 = 8'hf2 == io_state_in_15 ? 8'h89 : _GEN_4081; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4083 = 8'hf3 == io_state_in_15 ? 8'hd : _GEN_4082; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4084 = 8'hf4 == io_state_in_15 ? 8'hbf : _GEN_4083; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4085 = 8'hf5 == io_state_in_15 ? 8'he6 : _GEN_4084; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4086 = 8'hf6 == io_state_in_15 ? 8'h42 : _GEN_4085; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4087 = 8'hf7 == io_state_in_15 ? 8'h68 : _GEN_4086; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4088 = 8'hf8 == io_state_in_15 ? 8'h41 : _GEN_4087; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4089 = 8'hf9 == io_state_in_15 ? 8'h99 : _GEN_4088; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4090 = 8'hfa == io_state_in_15 ? 8'h2d : _GEN_4089; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4091 = 8'hfb == io_state_in_15 ? 8'hf : _GEN_4090; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4092 = 8'hfc == io_state_in_15 ? 8'hb0 : _GEN_4091; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4093 = 8'hfd == io_state_in_15 ? 8'h54 : _GEN_4092; // @[SubBytes.scala 35:{23,23}]
  wire [7:0] _GEN_4094 = 8'hfe == io_state_in_15 ? 8'hbb : _GEN_4093; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_0 = 8'hff == io_state_in_0 ? 8'h16 : _GEN_254; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_1 = 8'hff == io_state_in_1 ? 8'h16 : _GEN_510; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_2 = 8'hff == io_state_in_2 ? 8'h16 : _GEN_766; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_3 = 8'hff == io_state_in_3 ? 8'h16 : _GEN_1022; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_4 = 8'hff == io_state_in_4 ? 8'h16 : _GEN_1278; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_5 = 8'hff == io_state_in_5 ? 8'h16 : _GEN_1534; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_6 = 8'hff == io_state_in_6 ? 8'h16 : _GEN_1790; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_7 = 8'hff == io_state_in_7 ? 8'h16 : _GEN_2046; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_8 = 8'hff == io_state_in_8 ? 8'h16 : _GEN_2302; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_9 = 8'hff == io_state_in_9 ? 8'h16 : _GEN_2558; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_10 = 8'hff == io_state_in_10 ? 8'h16 : _GEN_2814; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_11 = 8'hff == io_state_in_11 ? 8'h16 : _GEN_3070; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_12 = 8'hff == io_state_in_12 ? 8'h16 : _GEN_3326; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_13 = 8'hff == io_state_in_13 ? 8'h16 : _GEN_3582; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_14 = 8'hff == io_state_in_14 ? 8'h16 : _GEN_3838; // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_15 = 8'hff == io_state_in_15 ? 8'h16 : _GEN_4094; // @[SubBytes.scala 35:{23,23}]
endmodule
module ShiftRows(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  assign io_state_out_0 = io_state_in_0; // @[ShiftRows.scala 13:19]
  assign io_state_out_1 = io_state_in_5; // @[ShiftRows.scala 14:19]
  assign io_state_out_2 = io_state_in_10; // @[ShiftRows.scala 15:19]
  assign io_state_out_3 = io_state_in_15; // @[ShiftRows.scala 16:19]
  assign io_state_out_4 = io_state_in_4; // @[ShiftRows.scala 18:19]
  assign io_state_out_5 = io_state_in_9; // @[ShiftRows.scala 19:19]
  assign io_state_out_6 = io_state_in_14; // @[ShiftRows.scala 20:19]
  assign io_state_out_7 = io_state_in_3; // @[ShiftRows.scala 21:19]
  assign io_state_out_8 = io_state_in_8; // @[ShiftRows.scala 23:19]
  assign io_state_out_9 = io_state_in_13; // @[ShiftRows.scala 24:19]
  assign io_state_out_10 = io_state_in_2; // @[ShiftRows.scala 25:20]
  assign io_state_out_11 = io_state_in_7; // @[ShiftRows.scala 26:20]
  assign io_state_out_12 = io_state_in_12; // @[ShiftRows.scala 28:20]
  assign io_state_out_13 = io_state_in_1; // @[ShiftRows.scala 29:20]
  assign io_state_out_14 = io_state_in_6; // @[ShiftRows.scala 30:20]
  assign io_state_out_15 = io_state_in_11; // @[ShiftRows.scala 31:20]
endmodule
module MixColumns(
  input  [7:0] io_state_in_0,
  input  [7:0] io_state_in_1,
  input  [7:0] io_state_in_2,
  input  [7:0] io_state_in_3,
  input  [7:0] io_state_in_4,
  input  [7:0] io_state_in_5,
  input  [7:0] io_state_in_6,
  input  [7:0] io_state_in_7,
  input  [7:0] io_state_in_8,
  input  [7:0] io_state_in_9,
  input  [7:0] io_state_in_10,
  input  [7:0] io_state_in_11,
  input  [7:0] io_state_in_12,
  input  [7:0] io_state_in_13,
  input  [7:0] io_state_in_14,
  input  [7:0] io_state_in_15,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15
);
  wire [7:0] _GEN_1 = 8'h1 == io_state_in_0 ? 8'h2 : 8'h0; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_2 = 8'h2 == io_state_in_0 ? 8'h4 : _GEN_1; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_3 = 8'h3 == io_state_in_0 ? 8'h6 : _GEN_2; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_4 = 8'h4 == io_state_in_0 ? 8'h8 : _GEN_3; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_5 = 8'h5 == io_state_in_0 ? 8'ha : _GEN_4; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_6 = 8'h6 == io_state_in_0 ? 8'hc : _GEN_5; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_7 = 8'h7 == io_state_in_0 ? 8'he : _GEN_6; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_8 = 8'h8 == io_state_in_0 ? 8'h10 : _GEN_7; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_9 = 8'h9 == io_state_in_0 ? 8'h12 : _GEN_8; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_10 = 8'ha == io_state_in_0 ? 8'h14 : _GEN_9; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_11 = 8'hb == io_state_in_0 ? 8'h16 : _GEN_10; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_12 = 8'hc == io_state_in_0 ? 8'h18 : _GEN_11; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_13 = 8'hd == io_state_in_0 ? 8'h1a : _GEN_12; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_14 = 8'he == io_state_in_0 ? 8'h1c : _GEN_13; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_15 = 8'hf == io_state_in_0 ? 8'h1e : _GEN_14; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_16 = 8'h10 == io_state_in_0 ? 8'h20 : _GEN_15; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_17 = 8'h11 == io_state_in_0 ? 8'h22 : _GEN_16; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_18 = 8'h12 == io_state_in_0 ? 8'h24 : _GEN_17; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_19 = 8'h13 == io_state_in_0 ? 8'h26 : _GEN_18; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_20 = 8'h14 == io_state_in_0 ? 8'h28 : _GEN_19; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_21 = 8'h15 == io_state_in_0 ? 8'h2a : _GEN_20; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_22 = 8'h16 == io_state_in_0 ? 8'h2c : _GEN_21; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_23 = 8'h17 == io_state_in_0 ? 8'h2e : _GEN_22; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_24 = 8'h18 == io_state_in_0 ? 8'h30 : _GEN_23; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_25 = 8'h19 == io_state_in_0 ? 8'h32 : _GEN_24; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_26 = 8'h1a == io_state_in_0 ? 8'h34 : _GEN_25; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_27 = 8'h1b == io_state_in_0 ? 8'h36 : _GEN_26; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_28 = 8'h1c == io_state_in_0 ? 8'h38 : _GEN_27; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_29 = 8'h1d == io_state_in_0 ? 8'h3a : _GEN_28; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_30 = 8'h1e == io_state_in_0 ? 8'h3c : _GEN_29; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_31 = 8'h1f == io_state_in_0 ? 8'h3e : _GEN_30; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_32 = 8'h20 == io_state_in_0 ? 8'h40 : _GEN_31; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_33 = 8'h21 == io_state_in_0 ? 8'h42 : _GEN_32; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_34 = 8'h22 == io_state_in_0 ? 8'h44 : _GEN_33; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_35 = 8'h23 == io_state_in_0 ? 8'h46 : _GEN_34; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_36 = 8'h24 == io_state_in_0 ? 8'h48 : _GEN_35; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_37 = 8'h25 == io_state_in_0 ? 8'h4a : _GEN_36; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_38 = 8'h26 == io_state_in_0 ? 8'h4c : _GEN_37; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_39 = 8'h27 == io_state_in_0 ? 8'h4e : _GEN_38; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_40 = 8'h28 == io_state_in_0 ? 8'h50 : _GEN_39; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_41 = 8'h29 == io_state_in_0 ? 8'h52 : _GEN_40; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_42 = 8'h2a == io_state_in_0 ? 8'h54 : _GEN_41; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_43 = 8'h2b == io_state_in_0 ? 8'h56 : _GEN_42; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_44 = 8'h2c == io_state_in_0 ? 8'h58 : _GEN_43; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_45 = 8'h2d == io_state_in_0 ? 8'h5a : _GEN_44; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_46 = 8'h2e == io_state_in_0 ? 8'h5c : _GEN_45; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_47 = 8'h2f == io_state_in_0 ? 8'h5e : _GEN_46; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_48 = 8'h30 == io_state_in_0 ? 8'h60 : _GEN_47; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_49 = 8'h31 == io_state_in_0 ? 8'h62 : _GEN_48; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_50 = 8'h32 == io_state_in_0 ? 8'h64 : _GEN_49; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_51 = 8'h33 == io_state_in_0 ? 8'h66 : _GEN_50; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_52 = 8'h34 == io_state_in_0 ? 8'h68 : _GEN_51; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_53 = 8'h35 == io_state_in_0 ? 8'h6a : _GEN_52; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_54 = 8'h36 == io_state_in_0 ? 8'h6c : _GEN_53; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_55 = 8'h37 == io_state_in_0 ? 8'h6e : _GEN_54; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_56 = 8'h38 == io_state_in_0 ? 8'h70 : _GEN_55; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_57 = 8'h39 == io_state_in_0 ? 8'h72 : _GEN_56; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_58 = 8'h3a == io_state_in_0 ? 8'h74 : _GEN_57; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_59 = 8'h3b == io_state_in_0 ? 8'h76 : _GEN_58; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_60 = 8'h3c == io_state_in_0 ? 8'h78 : _GEN_59; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_61 = 8'h3d == io_state_in_0 ? 8'h7a : _GEN_60; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_62 = 8'h3e == io_state_in_0 ? 8'h7c : _GEN_61; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_63 = 8'h3f == io_state_in_0 ? 8'h7e : _GEN_62; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_64 = 8'h40 == io_state_in_0 ? 8'h80 : _GEN_63; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_65 = 8'h41 == io_state_in_0 ? 8'h82 : _GEN_64; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_66 = 8'h42 == io_state_in_0 ? 8'h84 : _GEN_65; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_67 = 8'h43 == io_state_in_0 ? 8'h86 : _GEN_66; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_68 = 8'h44 == io_state_in_0 ? 8'h88 : _GEN_67; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_69 = 8'h45 == io_state_in_0 ? 8'h8a : _GEN_68; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_70 = 8'h46 == io_state_in_0 ? 8'h8c : _GEN_69; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_71 = 8'h47 == io_state_in_0 ? 8'h8e : _GEN_70; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_72 = 8'h48 == io_state_in_0 ? 8'h90 : _GEN_71; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_73 = 8'h49 == io_state_in_0 ? 8'h92 : _GEN_72; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_74 = 8'h4a == io_state_in_0 ? 8'h94 : _GEN_73; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_75 = 8'h4b == io_state_in_0 ? 8'h96 : _GEN_74; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_76 = 8'h4c == io_state_in_0 ? 8'h98 : _GEN_75; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_77 = 8'h4d == io_state_in_0 ? 8'h9a : _GEN_76; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_78 = 8'h4e == io_state_in_0 ? 8'h9c : _GEN_77; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_79 = 8'h4f == io_state_in_0 ? 8'h9e : _GEN_78; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_80 = 8'h50 == io_state_in_0 ? 8'ha0 : _GEN_79; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_81 = 8'h51 == io_state_in_0 ? 8'ha2 : _GEN_80; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_82 = 8'h52 == io_state_in_0 ? 8'ha4 : _GEN_81; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_83 = 8'h53 == io_state_in_0 ? 8'ha6 : _GEN_82; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_84 = 8'h54 == io_state_in_0 ? 8'ha8 : _GEN_83; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_85 = 8'h55 == io_state_in_0 ? 8'haa : _GEN_84; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_86 = 8'h56 == io_state_in_0 ? 8'hac : _GEN_85; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_87 = 8'h57 == io_state_in_0 ? 8'hae : _GEN_86; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_88 = 8'h58 == io_state_in_0 ? 8'hb0 : _GEN_87; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_89 = 8'h59 == io_state_in_0 ? 8'hb2 : _GEN_88; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_90 = 8'h5a == io_state_in_0 ? 8'hb4 : _GEN_89; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_91 = 8'h5b == io_state_in_0 ? 8'hb6 : _GEN_90; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_92 = 8'h5c == io_state_in_0 ? 8'hb8 : _GEN_91; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_93 = 8'h5d == io_state_in_0 ? 8'hba : _GEN_92; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_94 = 8'h5e == io_state_in_0 ? 8'hbc : _GEN_93; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_95 = 8'h5f == io_state_in_0 ? 8'hbe : _GEN_94; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_96 = 8'h60 == io_state_in_0 ? 8'hc0 : _GEN_95; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_97 = 8'h61 == io_state_in_0 ? 8'hc2 : _GEN_96; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_98 = 8'h62 == io_state_in_0 ? 8'hc4 : _GEN_97; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_99 = 8'h63 == io_state_in_0 ? 8'hc6 : _GEN_98; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_100 = 8'h64 == io_state_in_0 ? 8'hc8 : _GEN_99; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_101 = 8'h65 == io_state_in_0 ? 8'hca : _GEN_100; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_102 = 8'h66 == io_state_in_0 ? 8'hcc : _GEN_101; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_103 = 8'h67 == io_state_in_0 ? 8'hce : _GEN_102; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_104 = 8'h68 == io_state_in_0 ? 8'hd0 : _GEN_103; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_105 = 8'h69 == io_state_in_0 ? 8'hd2 : _GEN_104; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_106 = 8'h6a == io_state_in_0 ? 8'hd4 : _GEN_105; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_107 = 8'h6b == io_state_in_0 ? 8'hd6 : _GEN_106; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_108 = 8'h6c == io_state_in_0 ? 8'hd8 : _GEN_107; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_109 = 8'h6d == io_state_in_0 ? 8'hda : _GEN_108; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_110 = 8'h6e == io_state_in_0 ? 8'hdc : _GEN_109; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_111 = 8'h6f == io_state_in_0 ? 8'hde : _GEN_110; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_112 = 8'h70 == io_state_in_0 ? 8'he0 : _GEN_111; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_113 = 8'h71 == io_state_in_0 ? 8'he2 : _GEN_112; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_114 = 8'h72 == io_state_in_0 ? 8'he4 : _GEN_113; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_115 = 8'h73 == io_state_in_0 ? 8'he6 : _GEN_114; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_116 = 8'h74 == io_state_in_0 ? 8'he8 : _GEN_115; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_117 = 8'h75 == io_state_in_0 ? 8'hea : _GEN_116; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_118 = 8'h76 == io_state_in_0 ? 8'hec : _GEN_117; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_119 = 8'h77 == io_state_in_0 ? 8'hee : _GEN_118; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_120 = 8'h78 == io_state_in_0 ? 8'hf0 : _GEN_119; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_121 = 8'h79 == io_state_in_0 ? 8'hf2 : _GEN_120; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_122 = 8'h7a == io_state_in_0 ? 8'hf4 : _GEN_121; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_123 = 8'h7b == io_state_in_0 ? 8'hf6 : _GEN_122; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_124 = 8'h7c == io_state_in_0 ? 8'hf8 : _GEN_123; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_125 = 8'h7d == io_state_in_0 ? 8'hfa : _GEN_124; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_126 = 8'h7e == io_state_in_0 ? 8'hfc : _GEN_125; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_127 = 8'h7f == io_state_in_0 ? 8'hfe : _GEN_126; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_128 = 8'h80 == io_state_in_0 ? 8'h1b : _GEN_127; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_129 = 8'h81 == io_state_in_0 ? 8'h19 : _GEN_128; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_130 = 8'h82 == io_state_in_0 ? 8'h1f : _GEN_129; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_131 = 8'h83 == io_state_in_0 ? 8'h1d : _GEN_130; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_132 = 8'h84 == io_state_in_0 ? 8'h13 : _GEN_131; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_133 = 8'h85 == io_state_in_0 ? 8'h11 : _GEN_132; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_134 = 8'h86 == io_state_in_0 ? 8'h17 : _GEN_133; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_135 = 8'h87 == io_state_in_0 ? 8'h15 : _GEN_134; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_136 = 8'h88 == io_state_in_0 ? 8'hb : _GEN_135; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_137 = 8'h89 == io_state_in_0 ? 8'h9 : _GEN_136; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_138 = 8'h8a == io_state_in_0 ? 8'hf : _GEN_137; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_139 = 8'h8b == io_state_in_0 ? 8'hd : _GEN_138; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_140 = 8'h8c == io_state_in_0 ? 8'h3 : _GEN_139; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_141 = 8'h8d == io_state_in_0 ? 8'h1 : _GEN_140; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_142 = 8'h8e == io_state_in_0 ? 8'h7 : _GEN_141; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_143 = 8'h8f == io_state_in_0 ? 8'h5 : _GEN_142; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_144 = 8'h90 == io_state_in_0 ? 8'h3b : _GEN_143; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_145 = 8'h91 == io_state_in_0 ? 8'h39 : _GEN_144; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_146 = 8'h92 == io_state_in_0 ? 8'h3f : _GEN_145; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_147 = 8'h93 == io_state_in_0 ? 8'h3d : _GEN_146; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_148 = 8'h94 == io_state_in_0 ? 8'h33 : _GEN_147; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_149 = 8'h95 == io_state_in_0 ? 8'h31 : _GEN_148; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_150 = 8'h96 == io_state_in_0 ? 8'h37 : _GEN_149; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_151 = 8'h97 == io_state_in_0 ? 8'h35 : _GEN_150; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_152 = 8'h98 == io_state_in_0 ? 8'h2b : _GEN_151; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_153 = 8'h99 == io_state_in_0 ? 8'h29 : _GEN_152; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_154 = 8'h9a == io_state_in_0 ? 8'h2f : _GEN_153; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_155 = 8'h9b == io_state_in_0 ? 8'h2d : _GEN_154; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_156 = 8'h9c == io_state_in_0 ? 8'h23 : _GEN_155; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_157 = 8'h9d == io_state_in_0 ? 8'h21 : _GEN_156; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_158 = 8'h9e == io_state_in_0 ? 8'h27 : _GEN_157; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_159 = 8'h9f == io_state_in_0 ? 8'h25 : _GEN_158; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_160 = 8'ha0 == io_state_in_0 ? 8'h5b : _GEN_159; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_161 = 8'ha1 == io_state_in_0 ? 8'h59 : _GEN_160; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_162 = 8'ha2 == io_state_in_0 ? 8'h5f : _GEN_161; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_163 = 8'ha3 == io_state_in_0 ? 8'h5d : _GEN_162; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_164 = 8'ha4 == io_state_in_0 ? 8'h53 : _GEN_163; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_165 = 8'ha5 == io_state_in_0 ? 8'h51 : _GEN_164; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_166 = 8'ha6 == io_state_in_0 ? 8'h57 : _GEN_165; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_167 = 8'ha7 == io_state_in_0 ? 8'h55 : _GEN_166; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_168 = 8'ha8 == io_state_in_0 ? 8'h4b : _GEN_167; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_169 = 8'ha9 == io_state_in_0 ? 8'h49 : _GEN_168; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_170 = 8'haa == io_state_in_0 ? 8'h4f : _GEN_169; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_171 = 8'hab == io_state_in_0 ? 8'h4d : _GEN_170; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_172 = 8'hac == io_state_in_0 ? 8'h43 : _GEN_171; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_173 = 8'had == io_state_in_0 ? 8'h41 : _GEN_172; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_174 = 8'hae == io_state_in_0 ? 8'h47 : _GEN_173; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_175 = 8'haf == io_state_in_0 ? 8'h45 : _GEN_174; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_176 = 8'hb0 == io_state_in_0 ? 8'h7b : _GEN_175; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_177 = 8'hb1 == io_state_in_0 ? 8'h79 : _GEN_176; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_178 = 8'hb2 == io_state_in_0 ? 8'h7f : _GEN_177; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_179 = 8'hb3 == io_state_in_0 ? 8'h7d : _GEN_178; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_180 = 8'hb4 == io_state_in_0 ? 8'h73 : _GEN_179; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_181 = 8'hb5 == io_state_in_0 ? 8'h71 : _GEN_180; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_182 = 8'hb6 == io_state_in_0 ? 8'h77 : _GEN_181; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_183 = 8'hb7 == io_state_in_0 ? 8'h75 : _GEN_182; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_184 = 8'hb8 == io_state_in_0 ? 8'h6b : _GEN_183; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_185 = 8'hb9 == io_state_in_0 ? 8'h69 : _GEN_184; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_186 = 8'hba == io_state_in_0 ? 8'h6f : _GEN_185; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_187 = 8'hbb == io_state_in_0 ? 8'h6d : _GEN_186; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_188 = 8'hbc == io_state_in_0 ? 8'h63 : _GEN_187; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_189 = 8'hbd == io_state_in_0 ? 8'h61 : _GEN_188; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_190 = 8'hbe == io_state_in_0 ? 8'h67 : _GEN_189; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_191 = 8'hbf == io_state_in_0 ? 8'h65 : _GEN_190; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_192 = 8'hc0 == io_state_in_0 ? 8'h9b : _GEN_191; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_193 = 8'hc1 == io_state_in_0 ? 8'h99 : _GEN_192; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_194 = 8'hc2 == io_state_in_0 ? 8'h9f : _GEN_193; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_195 = 8'hc3 == io_state_in_0 ? 8'h9d : _GEN_194; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_196 = 8'hc4 == io_state_in_0 ? 8'h93 : _GEN_195; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_197 = 8'hc5 == io_state_in_0 ? 8'h91 : _GEN_196; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_198 = 8'hc6 == io_state_in_0 ? 8'h97 : _GEN_197; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_199 = 8'hc7 == io_state_in_0 ? 8'h95 : _GEN_198; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_200 = 8'hc8 == io_state_in_0 ? 8'h8b : _GEN_199; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_201 = 8'hc9 == io_state_in_0 ? 8'h89 : _GEN_200; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_202 = 8'hca == io_state_in_0 ? 8'h8f : _GEN_201; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_203 = 8'hcb == io_state_in_0 ? 8'h8d : _GEN_202; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_204 = 8'hcc == io_state_in_0 ? 8'h83 : _GEN_203; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_205 = 8'hcd == io_state_in_0 ? 8'h81 : _GEN_204; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_206 = 8'hce == io_state_in_0 ? 8'h87 : _GEN_205; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_207 = 8'hcf == io_state_in_0 ? 8'h85 : _GEN_206; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_208 = 8'hd0 == io_state_in_0 ? 8'hbb : _GEN_207; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_209 = 8'hd1 == io_state_in_0 ? 8'hb9 : _GEN_208; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_210 = 8'hd2 == io_state_in_0 ? 8'hbf : _GEN_209; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_211 = 8'hd3 == io_state_in_0 ? 8'hbd : _GEN_210; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_212 = 8'hd4 == io_state_in_0 ? 8'hb3 : _GEN_211; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_213 = 8'hd5 == io_state_in_0 ? 8'hb1 : _GEN_212; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_214 = 8'hd6 == io_state_in_0 ? 8'hb7 : _GEN_213; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_215 = 8'hd7 == io_state_in_0 ? 8'hb5 : _GEN_214; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_216 = 8'hd8 == io_state_in_0 ? 8'hab : _GEN_215; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_217 = 8'hd9 == io_state_in_0 ? 8'ha9 : _GEN_216; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_218 = 8'hda == io_state_in_0 ? 8'haf : _GEN_217; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_219 = 8'hdb == io_state_in_0 ? 8'had : _GEN_218; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_220 = 8'hdc == io_state_in_0 ? 8'ha3 : _GEN_219; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_221 = 8'hdd == io_state_in_0 ? 8'ha1 : _GEN_220; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_222 = 8'hde == io_state_in_0 ? 8'ha7 : _GEN_221; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_223 = 8'hdf == io_state_in_0 ? 8'ha5 : _GEN_222; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_224 = 8'he0 == io_state_in_0 ? 8'hdb : _GEN_223; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_225 = 8'he1 == io_state_in_0 ? 8'hd9 : _GEN_224; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_226 = 8'he2 == io_state_in_0 ? 8'hdf : _GEN_225; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_227 = 8'he3 == io_state_in_0 ? 8'hdd : _GEN_226; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_228 = 8'he4 == io_state_in_0 ? 8'hd3 : _GEN_227; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_229 = 8'he5 == io_state_in_0 ? 8'hd1 : _GEN_228; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_230 = 8'he6 == io_state_in_0 ? 8'hd7 : _GEN_229; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_231 = 8'he7 == io_state_in_0 ? 8'hd5 : _GEN_230; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_232 = 8'he8 == io_state_in_0 ? 8'hcb : _GEN_231; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_233 = 8'he9 == io_state_in_0 ? 8'hc9 : _GEN_232; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_234 = 8'hea == io_state_in_0 ? 8'hcf : _GEN_233; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_235 = 8'heb == io_state_in_0 ? 8'hcd : _GEN_234; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_236 = 8'hec == io_state_in_0 ? 8'hc3 : _GEN_235; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_237 = 8'hed == io_state_in_0 ? 8'hc1 : _GEN_236; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_238 = 8'hee == io_state_in_0 ? 8'hc7 : _GEN_237; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_239 = 8'hef == io_state_in_0 ? 8'hc5 : _GEN_238; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_240 = 8'hf0 == io_state_in_0 ? 8'hfb : _GEN_239; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_241 = 8'hf1 == io_state_in_0 ? 8'hf9 : _GEN_240; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_242 = 8'hf2 == io_state_in_0 ? 8'hff : _GEN_241; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_243 = 8'hf3 == io_state_in_0 ? 8'hfd : _GEN_242; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_244 = 8'hf4 == io_state_in_0 ? 8'hf3 : _GEN_243; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_245 = 8'hf5 == io_state_in_0 ? 8'hf1 : _GEN_244; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_246 = 8'hf6 == io_state_in_0 ? 8'hf7 : _GEN_245; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_247 = 8'hf7 == io_state_in_0 ? 8'hf5 : _GEN_246; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_248 = 8'hf8 == io_state_in_0 ? 8'heb : _GEN_247; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_249 = 8'hf9 == io_state_in_0 ? 8'he9 : _GEN_248; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_250 = 8'hfa == io_state_in_0 ? 8'hef : _GEN_249; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_251 = 8'hfb == io_state_in_0 ? 8'hed : _GEN_250; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_252 = 8'hfc == io_state_in_0 ? 8'he3 : _GEN_251; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_253 = 8'hfd == io_state_in_0 ? 8'he1 : _GEN_252; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_254 = 8'hfe == io_state_in_0 ? 8'he7 : _GEN_253; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_255 = 8'hff == io_state_in_0 ? 8'he5 : _GEN_254; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_257 = 8'h1 == io_state_in_1 ? 8'h3 : 8'h0; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_258 = 8'h2 == io_state_in_1 ? 8'h6 : _GEN_257; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_259 = 8'h3 == io_state_in_1 ? 8'h5 : _GEN_258; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_260 = 8'h4 == io_state_in_1 ? 8'hc : _GEN_259; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_261 = 8'h5 == io_state_in_1 ? 8'hf : _GEN_260; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_262 = 8'h6 == io_state_in_1 ? 8'ha : _GEN_261; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_263 = 8'h7 == io_state_in_1 ? 8'h9 : _GEN_262; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_264 = 8'h8 == io_state_in_1 ? 8'h18 : _GEN_263; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_265 = 8'h9 == io_state_in_1 ? 8'h1b : _GEN_264; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_266 = 8'ha == io_state_in_1 ? 8'h1e : _GEN_265; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_267 = 8'hb == io_state_in_1 ? 8'h1d : _GEN_266; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_268 = 8'hc == io_state_in_1 ? 8'h14 : _GEN_267; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_269 = 8'hd == io_state_in_1 ? 8'h17 : _GEN_268; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_270 = 8'he == io_state_in_1 ? 8'h12 : _GEN_269; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_271 = 8'hf == io_state_in_1 ? 8'h11 : _GEN_270; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_272 = 8'h10 == io_state_in_1 ? 8'h30 : _GEN_271; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_273 = 8'h11 == io_state_in_1 ? 8'h33 : _GEN_272; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_274 = 8'h12 == io_state_in_1 ? 8'h36 : _GEN_273; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_275 = 8'h13 == io_state_in_1 ? 8'h35 : _GEN_274; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_276 = 8'h14 == io_state_in_1 ? 8'h3c : _GEN_275; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_277 = 8'h15 == io_state_in_1 ? 8'h3f : _GEN_276; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_278 = 8'h16 == io_state_in_1 ? 8'h3a : _GEN_277; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_279 = 8'h17 == io_state_in_1 ? 8'h39 : _GEN_278; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_280 = 8'h18 == io_state_in_1 ? 8'h28 : _GEN_279; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_281 = 8'h19 == io_state_in_1 ? 8'h2b : _GEN_280; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_282 = 8'h1a == io_state_in_1 ? 8'h2e : _GEN_281; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_283 = 8'h1b == io_state_in_1 ? 8'h2d : _GEN_282; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_284 = 8'h1c == io_state_in_1 ? 8'h24 : _GEN_283; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_285 = 8'h1d == io_state_in_1 ? 8'h27 : _GEN_284; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_286 = 8'h1e == io_state_in_1 ? 8'h22 : _GEN_285; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_287 = 8'h1f == io_state_in_1 ? 8'h21 : _GEN_286; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_288 = 8'h20 == io_state_in_1 ? 8'h60 : _GEN_287; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_289 = 8'h21 == io_state_in_1 ? 8'h63 : _GEN_288; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_290 = 8'h22 == io_state_in_1 ? 8'h66 : _GEN_289; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_291 = 8'h23 == io_state_in_1 ? 8'h65 : _GEN_290; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_292 = 8'h24 == io_state_in_1 ? 8'h6c : _GEN_291; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_293 = 8'h25 == io_state_in_1 ? 8'h6f : _GEN_292; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_294 = 8'h26 == io_state_in_1 ? 8'h6a : _GEN_293; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_295 = 8'h27 == io_state_in_1 ? 8'h69 : _GEN_294; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_296 = 8'h28 == io_state_in_1 ? 8'h78 : _GEN_295; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_297 = 8'h29 == io_state_in_1 ? 8'h7b : _GEN_296; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_298 = 8'h2a == io_state_in_1 ? 8'h7e : _GEN_297; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_299 = 8'h2b == io_state_in_1 ? 8'h7d : _GEN_298; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_300 = 8'h2c == io_state_in_1 ? 8'h74 : _GEN_299; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_301 = 8'h2d == io_state_in_1 ? 8'h77 : _GEN_300; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_302 = 8'h2e == io_state_in_1 ? 8'h72 : _GEN_301; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_303 = 8'h2f == io_state_in_1 ? 8'h71 : _GEN_302; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_304 = 8'h30 == io_state_in_1 ? 8'h50 : _GEN_303; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_305 = 8'h31 == io_state_in_1 ? 8'h53 : _GEN_304; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_306 = 8'h32 == io_state_in_1 ? 8'h56 : _GEN_305; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_307 = 8'h33 == io_state_in_1 ? 8'h55 : _GEN_306; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_308 = 8'h34 == io_state_in_1 ? 8'h5c : _GEN_307; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_309 = 8'h35 == io_state_in_1 ? 8'h5f : _GEN_308; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_310 = 8'h36 == io_state_in_1 ? 8'h5a : _GEN_309; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_311 = 8'h37 == io_state_in_1 ? 8'h59 : _GEN_310; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_312 = 8'h38 == io_state_in_1 ? 8'h48 : _GEN_311; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_313 = 8'h39 == io_state_in_1 ? 8'h4b : _GEN_312; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_314 = 8'h3a == io_state_in_1 ? 8'h4e : _GEN_313; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_315 = 8'h3b == io_state_in_1 ? 8'h4d : _GEN_314; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_316 = 8'h3c == io_state_in_1 ? 8'h44 : _GEN_315; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_317 = 8'h3d == io_state_in_1 ? 8'h47 : _GEN_316; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_318 = 8'h3e == io_state_in_1 ? 8'h42 : _GEN_317; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_319 = 8'h3f == io_state_in_1 ? 8'h41 : _GEN_318; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_320 = 8'h40 == io_state_in_1 ? 8'hc0 : _GEN_319; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_321 = 8'h41 == io_state_in_1 ? 8'hc3 : _GEN_320; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_322 = 8'h42 == io_state_in_1 ? 8'hc6 : _GEN_321; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_323 = 8'h43 == io_state_in_1 ? 8'hc5 : _GEN_322; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_324 = 8'h44 == io_state_in_1 ? 8'hcc : _GEN_323; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_325 = 8'h45 == io_state_in_1 ? 8'hcf : _GEN_324; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_326 = 8'h46 == io_state_in_1 ? 8'hca : _GEN_325; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_327 = 8'h47 == io_state_in_1 ? 8'hc9 : _GEN_326; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_328 = 8'h48 == io_state_in_1 ? 8'hd8 : _GEN_327; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_329 = 8'h49 == io_state_in_1 ? 8'hdb : _GEN_328; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_330 = 8'h4a == io_state_in_1 ? 8'hde : _GEN_329; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_331 = 8'h4b == io_state_in_1 ? 8'hdd : _GEN_330; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_332 = 8'h4c == io_state_in_1 ? 8'hd4 : _GEN_331; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_333 = 8'h4d == io_state_in_1 ? 8'hd7 : _GEN_332; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_334 = 8'h4e == io_state_in_1 ? 8'hd2 : _GEN_333; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_335 = 8'h4f == io_state_in_1 ? 8'hd1 : _GEN_334; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_336 = 8'h50 == io_state_in_1 ? 8'hf0 : _GEN_335; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_337 = 8'h51 == io_state_in_1 ? 8'hf3 : _GEN_336; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_338 = 8'h52 == io_state_in_1 ? 8'hf6 : _GEN_337; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_339 = 8'h53 == io_state_in_1 ? 8'hf5 : _GEN_338; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_340 = 8'h54 == io_state_in_1 ? 8'hfc : _GEN_339; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_341 = 8'h55 == io_state_in_1 ? 8'hff : _GEN_340; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_342 = 8'h56 == io_state_in_1 ? 8'hfa : _GEN_341; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_343 = 8'h57 == io_state_in_1 ? 8'hf9 : _GEN_342; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_344 = 8'h58 == io_state_in_1 ? 8'he8 : _GEN_343; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_345 = 8'h59 == io_state_in_1 ? 8'heb : _GEN_344; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_346 = 8'h5a == io_state_in_1 ? 8'hee : _GEN_345; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_347 = 8'h5b == io_state_in_1 ? 8'hed : _GEN_346; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_348 = 8'h5c == io_state_in_1 ? 8'he4 : _GEN_347; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_349 = 8'h5d == io_state_in_1 ? 8'he7 : _GEN_348; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_350 = 8'h5e == io_state_in_1 ? 8'he2 : _GEN_349; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_351 = 8'h5f == io_state_in_1 ? 8'he1 : _GEN_350; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_352 = 8'h60 == io_state_in_1 ? 8'ha0 : _GEN_351; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_353 = 8'h61 == io_state_in_1 ? 8'ha3 : _GEN_352; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_354 = 8'h62 == io_state_in_1 ? 8'ha6 : _GEN_353; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_355 = 8'h63 == io_state_in_1 ? 8'ha5 : _GEN_354; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_356 = 8'h64 == io_state_in_1 ? 8'hac : _GEN_355; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_357 = 8'h65 == io_state_in_1 ? 8'haf : _GEN_356; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_358 = 8'h66 == io_state_in_1 ? 8'haa : _GEN_357; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_359 = 8'h67 == io_state_in_1 ? 8'ha9 : _GEN_358; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_360 = 8'h68 == io_state_in_1 ? 8'hb8 : _GEN_359; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_361 = 8'h69 == io_state_in_1 ? 8'hbb : _GEN_360; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_362 = 8'h6a == io_state_in_1 ? 8'hbe : _GEN_361; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_363 = 8'h6b == io_state_in_1 ? 8'hbd : _GEN_362; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_364 = 8'h6c == io_state_in_1 ? 8'hb4 : _GEN_363; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_365 = 8'h6d == io_state_in_1 ? 8'hb7 : _GEN_364; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_366 = 8'h6e == io_state_in_1 ? 8'hb2 : _GEN_365; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_367 = 8'h6f == io_state_in_1 ? 8'hb1 : _GEN_366; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_368 = 8'h70 == io_state_in_1 ? 8'h90 : _GEN_367; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_369 = 8'h71 == io_state_in_1 ? 8'h93 : _GEN_368; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_370 = 8'h72 == io_state_in_1 ? 8'h96 : _GEN_369; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_371 = 8'h73 == io_state_in_1 ? 8'h95 : _GEN_370; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_372 = 8'h74 == io_state_in_1 ? 8'h9c : _GEN_371; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_373 = 8'h75 == io_state_in_1 ? 8'h9f : _GEN_372; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_374 = 8'h76 == io_state_in_1 ? 8'h9a : _GEN_373; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_375 = 8'h77 == io_state_in_1 ? 8'h99 : _GEN_374; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_376 = 8'h78 == io_state_in_1 ? 8'h88 : _GEN_375; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_377 = 8'h79 == io_state_in_1 ? 8'h8b : _GEN_376; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_378 = 8'h7a == io_state_in_1 ? 8'h8e : _GEN_377; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_379 = 8'h7b == io_state_in_1 ? 8'h8d : _GEN_378; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_380 = 8'h7c == io_state_in_1 ? 8'h84 : _GEN_379; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_381 = 8'h7d == io_state_in_1 ? 8'h87 : _GEN_380; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_382 = 8'h7e == io_state_in_1 ? 8'h82 : _GEN_381; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_383 = 8'h7f == io_state_in_1 ? 8'h81 : _GEN_382; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_384 = 8'h80 == io_state_in_1 ? 8'h9b : _GEN_383; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_385 = 8'h81 == io_state_in_1 ? 8'h98 : _GEN_384; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_386 = 8'h82 == io_state_in_1 ? 8'h9d : _GEN_385; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_387 = 8'h83 == io_state_in_1 ? 8'h9e : _GEN_386; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_388 = 8'h84 == io_state_in_1 ? 8'h97 : _GEN_387; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_389 = 8'h85 == io_state_in_1 ? 8'h94 : _GEN_388; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_390 = 8'h86 == io_state_in_1 ? 8'h91 : _GEN_389; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_391 = 8'h87 == io_state_in_1 ? 8'h92 : _GEN_390; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_392 = 8'h88 == io_state_in_1 ? 8'h83 : _GEN_391; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_393 = 8'h89 == io_state_in_1 ? 8'h80 : _GEN_392; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_394 = 8'h8a == io_state_in_1 ? 8'h85 : _GEN_393; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_395 = 8'h8b == io_state_in_1 ? 8'h86 : _GEN_394; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_396 = 8'h8c == io_state_in_1 ? 8'h8f : _GEN_395; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_397 = 8'h8d == io_state_in_1 ? 8'h8c : _GEN_396; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_398 = 8'h8e == io_state_in_1 ? 8'h89 : _GEN_397; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_399 = 8'h8f == io_state_in_1 ? 8'h8a : _GEN_398; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_400 = 8'h90 == io_state_in_1 ? 8'hab : _GEN_399; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_401 = 8'h91 == io_state_in_1 ? 8'ha8 : _GEN_400; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_402 = 8'h92 == io_state_in_1 ? 8'had : _GEN_401; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_403 = 8'h93 == io_state_in_1 ? 8'hae : _GEN_402; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_404 = 8'h94 == io_state_in_1 ? 8'ha7 : _GEN_403; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_405 = 8'h95 == io_state_in_1 ? 8'ha4 : _GEN_404; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_406 = 8'h96 == io_state_in_1 ? 8'ha1 : _GEN_405; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_407 = 8'h97 == io_state_in_1 ? 8'ha2 : _GEN_406; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_408 = 8'h98 == io_state_in_1 ? 8'hb3 : _GEN_407; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_409 = 8'h99 == io_state_in_1 ? 8'hb0 : _GEN_408; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_410 = 8'h9a == io_state_in_1 ? 8'hb5 : _GEN_409; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_411 = 8'h9b == io_state_in_1 ? 8'hb6 : _GEN_410; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_412 = 8'h9c == io_state_in_1 ? 8'hbf : _GEN_411; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_413 = 8'h9d == io_state_in_1 ? 8'hbc : _GEN_412; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_414 = 8'h9e == io_state_in_1 ? 8'hb9 : _GEN_413; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_415 = 8'h9f == io_state_in_1 ? 8'hba : _GEN_414; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_416 = 8'ha0 == io_state_in_1 ? 8'hfb : _GEN_415; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_417 = 8'ha1 == io_state_in_1 ? 8'hf8 : _GEN_416; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_418 = 8'ha2 == io_state_in_1 ? 8'hfd : _GEN_417; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_419 = 8'ha3 == io_state_in_1 ? 8'hfe : _GEN_418; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_420 = 8'ha4 == io_state_in_1 ? 8'hf7 : _GEN_419; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_421 = 8'ha5 == io_state_in_1 ? 8'hf4 : _GEN_420; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_422 = 8'ha6 == io_state_in_1 ? 8'hf1 : _GEN_421; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_423 = 8'ha7 == io_state_in_1 ? 8'hf2 : _GEN_422; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_424 = 8'ha8 == io_state_in_1 ? 8'he3 : _GEN_423; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_425 = 8'ha9 == io_state_in_1 ? 8'he0 : _GEN_424; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_426 = 8'haa == io_state_in_1 ? 8'he5 : _GEN_425; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_427 = 8'hab == io_state_in_1 ? 8'he6 : _GEN_426; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_428 = 8'hac == io_state_in_1 ? 8'hef : _GEN_427; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_429 = 8'had == io_state_in_1 ? 8'hec : _GEN_428; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_430 = 8'hae == io_state_in_1 ? 8'he9 : _GEN_429; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_431 = 8'haf == io_state_in_1 ? 8'hea : _GEN_430; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_432 = 8'hb0 == io_state_in_1 ? 8'hcb : _GEN_431; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_433 = 8'hb1 == io_state_in_1 ? 8'hc8 : _GEN_432; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_434 = 8'hb2 == io_state_in_1 ? 8'hcd : _GEN_433; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_435 = 8'hb3 == io_state_in_1 ? 8'hce : _GEN_434; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_436 = 8'hb4 == io_state_in_1 ? 8'hc7 : _GEN_435; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_437 = 8'hb5 == io_state_in_1 ? 8'hc4 : _GEN_436; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_438 = 8'hb6 == io_state_in_1 ? 8'hc1 : _GEN_437; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_439 = 8'hb7 == io_state_in_1 ? 8'hc2 : _GEN_438; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_440 = 8'hb8 == io_state_in_1 ? 8'hd3 : _GEN_439; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_441 = 8'hb9 == io_state_in_1 ? 8'hd0 : _GEN_440; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_442 = 8'hba == io_state_in_1 ? 8'hd5 : _GEN_441; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_443 = 8'hbb == io_state_in_1 ? 8'hd6 : _GEN_442; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_444 = 8'hbc == io_state_in_1 ? 8'hdf : _GEN_443; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_445 = 8'hbd == io_state_in_1 ? 8'hdc : _GEN_444; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_446 = 8'hbe == io_state_in_1 ? 8'hd9 : _GEN_445; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_447 = 8'hbf == io_state_in_1 ? 8'hda : _GEN_446; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_448 = 8'hc0 == io_state_in_1 ? 8'h5b : _GEN_447; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_449 = 8'hc1 == io_state_in_1 ? 8'h58 : _GEN_448; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_450 = 8'hc2 == io_state_in_1 ? 8'h5d : _GEN_449; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_451 = 8'hc3 == io_state_in_1 ? 8'h5e : _GEN_450; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_452 = 8'hc4 == io_state_in_1 ? 8'h57 : _GEN_451; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_453 = 8'hc5 == io_state_in_1 ? 8'h54 : _GEN_452; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_454 = 8'hc6 == io_state_in_1 ? 8'h51 : _GEN_453; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_455 = 8'hc7 == io_state_in_1 ? 8'h52 : _GEN_454; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_456 = 8'hc8 == io_state_in_1 ? 8'h43 : _GEN_455; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_457 = 8'hc9 == io_state_in_1 ? 8'h40 : _GEN_456; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_458 = 8'hca == io_state_in_1 ? 8'h45 : _GEN_457; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_459 = 8'hcb == io_state_in_1 ? 8'h46 : _GEN_458; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_460 = 8'hcc == io_state_in_1 ? 8'h4f : _GEN_459; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_461 = 8'hcd == io_state_in_1 ? 8'h4c : _GEN_460; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_462 = 8'hce == io_state_in_1 ? 8'h49 : _GEN_461; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_463 = 8'hcf == io_state_in_1 ? 8'h4a : _GEN_462; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_464 = 8'hd0 == io_state_in_1 ? 8'h6b : _GEN_463; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_465 = 8'hd1 == io_state_in_1 ? 8'h68 : _GEN_464; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_466 = 8'hd2 == io_state_in_1 ? 8'h6d : _GEN_465; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_467 = 8'hd3 == io_state_in_1 ? 8'h6e : _GEN_466; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_468 = 8'hd4 == io_state_in_1 ? 8'h67 : _GEN_467; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_469 = 8'hd5 == io_state_in_1 ? 8'h64 : _GEN_468; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_470 = 8'hd6 == io_state_in_1 ? 8'h61 : _GEN_469; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_471 = 8'hd7 == io_state_in_1 ? 8'h62 : _GEN_470; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_472 = 8'hd8 == io_state_in_1 ? 8'h73 : _GEN_471; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_473 = 8'hd9 == io_state_in_1 ? 8'h70 : _GEN_472; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_474 = 8'hda == io_state_in_1 ? 8'h75 : _GEN_473; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_475 = 8'hdb == io_state_in_1 ? 8'h76 : _GEN_474; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_476 = 8'hdc == io_state_in_1 ? 8'h7f : _GEN_475; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_477 = 8'hdd == io_state_in_1 ? 8'h7c : _GEN_476; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_478 = 8'hde == io_state_in_1 ? 8'h79 : _GEN_477; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_479 = 8'hdf == io_state_in_1 ? 8'h7a : _GEN_478; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_480 = 8'he0 == io_state_in_1 ? 8'h3b : _GEN_479; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_481 = 8'he1 == io_state_in_1 ? 8'h38 : _GEN_480; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_482 = 8'he2 == io_state_in_1 ? 8'h3d : _GEN_481; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_483 = 8'he3 == io_state_in_1 ? 8'h3e : _GEN_482; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_484 = 8'he4 == io_state_in_1 ? 8'h37 : _GEN_483; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_485 = 8'he5 == io_state_in_1 ? 8'h34 : _GEN_484; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_486 = 8'he6 == io_state_in_1 ? 8'h31 : _GEN_485; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_487 = 8'he7 == io_state_in_1 ? 8'h32 : _GEN_486; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_488 = 8'he8 == io_state_in_1 ? 8'h23 : _GEN_487; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_489 = 8'he9 == io_state_in_1 ? 8'h20 : _GEN_488; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_490 = 8'hea == io_state_in_1 ? 8'h25 : _GEN_489; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_491 = 8'heb == io_state_in_1 ? 8'h26 : _GEN_490; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_492 = 8'hec == io_state_in_1 ? 8'h2f : _GEN_491; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_493 = 8'hed == io_state_in_1 ? 8'h2c : _GEN_492; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_494 = 8'hee == io_state_in_1 ? 8'h29 : _GEN_493; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_495 = 8'hef == io_state_in_1 ? 8'h2a : _GEN_494; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_496 = 8'hf0 == io_state_in_1 ? 8'hb : _GEN_495; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_497 = 8'hf1 == io_state_in_1 ? 8'h8 : _GEN_496; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_498 = 8'hf2 == io_state_in_1 ? 8'hd : _GEN_497; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_499 = 8'hf3 == io_state_in_1 ? 8'he : _GEN_498; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_500 = 8'hf4 == io_state_in_1 ? 8'h7 : _GEN_499; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_501 = 8'hf5 == io_state_in_1 ? 8'h4 : _GEN_500; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_502 = 8'hf6 == io_state_in_1 ? 8'h1 : _GEN_501; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_503 = 8'hf7 == io_state_in_1 ? 8'h2 : _GEN_502; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_504 = 8'hf8 == io_state_in_1 ? 8'h13 : _GEN_503; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_505 = 8'hf9 == io_state_in_1 ? 8'h10 : _GEN_504; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_506 = 8'hfa == io_state_in_1 ? 8'h15 : _GEN_505; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_507 = 8'hfb == io_state_in_1 ? 8'h16 : _GEN_506; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_508 = 8'hfc == io_state_in_1 ? 8'h1f : _GEN_507; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_509 = 8'hfd == io_state_in_1 ? 8'h1c : _GEN_508; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_510 = 8'hfe == io_state_in_1 ? 8'h19 : _GEN_509; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _GEN_511 = 8'hff == io_state_in_1 ? 8'h1a : _GEN_510; // @[MixColumns.scala 125:{41,41}]
  wire [7:0] _tmp_state_0_T = _GEN_255 ^ _GEN_511; // @[MixColumns.scala 125:41]
  wire [7:0] _tmp_state_0_T_1 = _tmp_state_0_T ^ io_state_in_2; // @[MixColumns.scala 125:65]
  wire [7:0] _GEN_513 = 8'h1 == io_state_in_1 ? 8'h2 : 8'h0; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_514 = 8'h2 == io_state_in_1 ? 8'h4 : _GEN_513; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_515 = 8'h3 == io_state_in_1 ? 8'h6 : _GEN_514; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_516 = 8'h4 == io_state_in_1 ? 8'h8 : _GEN_515; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_517 = 8'h5 == io_state_in_1 ? 8'ha : _GEN_516; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_518 = 8'h6 == io_state_in_1 ? 8'hc : _GEN_517; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_519 = 8'h7 == io_state_in_1 ? 8'he : _GEN_518; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_520 = 8'h8 == io_state_in_1 ? 8'h10 : _GEN_519; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_521 = 8'h9 == io_state_in_1 ? 8'h12 : _GEN_520; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_522 = 8'ha == io_state_in_1 ? 8'h14 : _GEN_521; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_523 = 8'hb == io_state_in_1 ? 8'h16 : _GEN_522; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_524 = 8'hc == io_state_in_1 ? 8'h18 : _GEN_523; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_525 = 8'hd == io_state_in_1 ? 8'h1a : _GEN_524; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_526 = 8'he == io_state_in_1 ? 8'h1c : _GEN_525; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_527 = 8'hf == io_state_in_1 ? 8'h1e : _GEN_526; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_528 = 8'h10 == io_state_in_1 ? 8'h20 : _GEN_527; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_529 = 8'h11 == io_state_in_1 ? 8'h22 : _GEN_528; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_530 = 8'h12 == io_state_in_1 ? 8'h24 : _GEN_529; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_531 = 8'h13 == io_state_in_1 ? 8'h26 : _GEN_530; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_532 = 8'h14 == io_state_in_1 ? 8'h28 : _GEN_531; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_533 = 8'h15 == io_state_in_1 ? 8'h2a : _GEN_532; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_534 = 8'h16 == io_state_in_1 ? 8'h2c : _GEN_533; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_535 = 8'h17 == io_state_in_1 ? 8'h2e : _GEN_534; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_536 = 8'h18 == io_state_in_1 ? 8'h30 : _GEN_535; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_537 = 8'h19 == io_state_in_1 ? 8'h32 : _GEN_536; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_538 = 8'h1a == io_state_in_1 ? 8'h34 : _GEN_537; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_539 = 8'h1b == io_state_in_1 ? 8'h36 : _GEN_538; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_540 = 8'h1c == io_state_in_1 ? 8'h38 : _GEN_539; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_541 = 8'h1d == io_state_in_1 ? 8'h3a : _GEN_540; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_542 = 8'h1e == io_state_in_1 ? 8'h3c : _GEN_541; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_543 = 8'h1f == io_state_in_1 ? 8'h3e : _GEN_542; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_544 = 8'h20 == io_state_in_1 ? 8'h40 : _GEN_543; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_545 = 8'h21 == io_state_in_1 ? 8'h42 : _GEN_544; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_546 = 8'h22 == io_state_in_1 ? 8'h44 : _GEN_545; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_547 = 8'h23 == io_state_in_1 ? 8'h46 : _GEN_546; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_548 = 8'h24 == io_state_in_1 ? 8'h48 : _GEN_547; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_549 = 8'h25 == io_state_in_1 ? 8'h4a : _GEN_548; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_550 = 8'h26 == io_state_in_1 ? 8'h4c : _GEN_549; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_551 = 8'h27 == io_state_in_1 ? 8'h4e : _GEN_550; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_552 = 8'h28 == io_state_in_1 ? 8'h50 : _GEN_551; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_553 = 8'h29 == io_state_in_1 ? 8'h52 : _GEN_552; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_554 = 8'h2a == io_state_in_1 ? 8'h54 : _GEN_553; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_555 = 8'h2b == io_state_in_1 ? 8'h56 : _GEN_554; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_556 = 8'h2c == io_state_in_1 ? 8'h58 : _GEN_555; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_557 = 8'h2d == io_state_in_1 ? 8'h5a : _GEN_556; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_558 = 8'h2e == io_state_in_1 ? 8'h5c : _GEN_557; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_559 = 8'h2f == io_state_in_1 ? 8'h5e : _GEN_558; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_560 = 8'h30 == io_state_in_1 ? 8'h60 : _GEN_559; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_561 = 8'h31 == io_state_in_1 ? 8'h62 : _GEN_560; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_562 = 8'h32 == io_state_in_1 ? 8'h64 : _GEN_561; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_563 = 8'h33 == io_state_in_1 ? 8'h66 : _GEN_562; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_564 = 8'h34 == io_state_in_1 ? 8'h68 : _GEN_563; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_565 = 8'h35 == io_state_in_1 ? 8'h6a : _GEN_564; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_566 = 8'h36 == io_state_in_1 ? 8'h6c : _GEN_565; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_567 = 8'h37 == io_state_in_1 ? 8'h6e : _GEN_566; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_568 = 8'h38 == io_state_in_1 ? 8'h70 : _GEN_567; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_569 = 8'h39 == io_state_in_1 ? 8'h72 : _GEN_568; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_570 = 8'h3a == io_state_in_1 ? 8'h74 : _GEN_569; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_571 = 8'h3b == io_state_in_1 ? 8'h76 : _GEN_570; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_572 = 8'h3c == io_state_in_1 ? 8'h78 : _GEN_571; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_573 = 8'h3d == io_state_in_1 ? 8'h7a : _GEN_572; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_574 = 8'h3e == io_state_in_1 ? 8'h7c : _GEN_573; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_575 = 8'h3f == io_state_in_1 ? 8'h7e : _GEN_574; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_576 = 8'h40 == io_state_in_1 ? 8'h80 : _GEN_575; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_577 = 8'h41 == io_state_in_1 ? 8'h82 : _GEN_576; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_578 = 8'h42 == io_state_in_1 ? 8'h84 : _GEN_577; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_579 = 8'h43 == io_state_in_1 ? 8'h86 : _GEN_578; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_580 = 8'h44 == io_state_in_1 ? 8'h88 : _GEN_579; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_581 = 8'h45 == io_state_in_1 ? 8'h8a : _GEN_580; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_582 = 8'h46 == io_state_in_1 ? 8'h8c : _GEN_581; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_583 = 8'h47 == io_state_in_1 ? 8'h8e : _GEN_582; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_584 = 8'h48 == io_state_in_1 ? 8'h90 : _GEN_583; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_585 = 8'h49 == io_state_in_1 ? 8'h92 : _GEN_584; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_586 = 8'h4a == io_state_in_1 ? 8'h94 : _GEN_585; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_587 = 8'h4b == io_state_in_1 ? 8'h96 : _GEN_586; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_588 = 8'h4c == io_state_in_1 ? 8'h98 : _GEN_587; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_589 = 8'h4d == io_state_in_1 ? 8'h9a : _GEN_588; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_590 = 8'h4e == io_state_in_1 ? 8'h9c : _GEN_589; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_591 = 8'h4f == io_state_in_1 ? 8'h9e : _GEN_590; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_592 = 8'h50 == io_state_in_1 ? 8'ha0 : _GEN_591; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_593 = 8'h51 == io_state_in_1 ? 8'ha2 : _GEN_592; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_594 = 8'h52 == io_state_in_1 ? 8'ha4 : _GEN_593; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_595 = 8'h53 == io_state_in_1 ? 8'ha6 : _GEN_594; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_596 = 8'h54 == io_state_in_1 ? 8'ha8 : _GEN_595; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_597 = 8'h55 == io_state_in_1 ? 8'haa : _GEN_596; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_598 = 8'h56 == io_state_in_1 ? 8'hac : _GEN_597; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_599 = 8'h57 == io_state_in_1 ? 8'hae : _GEN_598; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_600 = 8'h58 == io_state_in_1 ? 8'hb0 : _GEN_599; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_601 = 8'h59 == io_state_in_1 ? 8'hb2 : _GEN_600; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_602 = 8'h5a == io_state_in_1 ? 8'hb4 : _GEN_601; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_603 = 8'h5b == io_state_in_1 ? 8'hb6 : _GEN_602; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_604 = 8'h5c == io_state_in_1 ? 8'hb8 : _GEN_603; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_605 = 8'h5d == io_state_in_1 ? 8'hba : _GEN_604; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_606 = 8'h5e == io_state_in_1 ? 8'hbc : _GEN_605; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_607 = 8'h5f == io_state_in_1 ? 8'hbe : _GEN_606; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_608 = 8'h60 == io_state_in_1 ? 8'hc0 : _GEN_607; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_609 = 8'h61 == io_state_in_1 ? 8'hc2 : _GEN_608; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_610 = 8'h62 == io_state_in_1 ? 8'hc4 : _GEN_609; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_611 = 8'h63 == io_state_in_1 ? 8'hc6 : _GEN_610; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_612 = 8'h64 == io_state_in_1 ? 8'hc8 : _GEN_611; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_613 = 8'h65 == io_state_in_1 ? 8'hca : _GEN_612; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_614 = 8'h66 == io_state_in_1 ? 8'hcc : _GEN_613; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_615 = 8'h67 == io_state_in_1 ? 8'hce : _GEN_614; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_616 = 8'h68 == io_state_in_1 ? 8'hd0 : _GEN_615; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_617 = 8'h69 == io_state_in_1 ? 8'hd2 : _GEN_616; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_618 = 8'h6a == io_state_in_1 ? 8'hd4 : _GEN_617; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_619 = 8'h6b == io_state_in_1 ? 8'hd6 : _GEN_618; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_620 = 8'h6c == io_state_in_1 ? 8'hd8 : _GEN_619; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_621 = 8'h6d == io_state_in_1 ? 8'hda : _GEN_620; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_622 = 8'h6e == io_state_in_1 ? 8'hdc : _GEN_621; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_623 = 8'h6f == io_state_in_1 ? 8'hde : _GEN_622; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_624 = 8'h70 == io_state_in_1 ? 8'he0 : _GEN_623; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_625 = 8'h71 == io_state_in_1 ? 8'he2 : _GEN_624; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_626 = 8'h72 == io_state_in_1 ? 8'he4 : _GEN_625; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_627 = 8'h73 == io_state_in_1 ? 8'he6 : _GEN_626; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_628 = 8'h74 == io_state_in_1 ? 8'he8 : _GEN_627; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_629 = 8'h75 == io_state_in_1 ? 8'hea : _GEN_628; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_630 = 8'h76 == io_state_in_1 ? 8'hec : _GEN_629; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_631 = 8'h77 == io_state_in_1 ? 8'hee : _GEN_630; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_632 = 8'h78 == io_state_in_1 ? 8'hf0 : _GEN_631; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_633 = 8'h79 == io_state_in_1 ? 8'hf2 : _GEN_632; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_634 = 8'h7a == io_state_in_1 ? 8'hf4 : _GEN_633; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_635 = 8'h7b == io_state_in_1 ? 8'hf6 : _GEN_634; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_636 = 8'h7c == io_state_in_1 ? 8'hf8 : _GEN_635; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_637 = 8'h7d == io_state_in_1 ? 8'hfa : _GEN_636; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_638 = 8'h7e == io_state_in_1 ? 8'hfc : _GEN_637; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_639 = 8'h7f == io_state_in_1 ? 8'hfe : _GEN_638; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_640 = 8'h80 == io_state_in_1 ? 8'h1b : _GEN_639; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_641 = 8'h81 == io_state_in_1 ? 8'h19 : _GEN_640; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_642 = 8'h82 == io_state_in_1 ? 8'h1f : _GEN_641; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_643 = 8'h83 == io_state_in_1 ? 8'h1d : _GEN_642; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_644 = 8'h84 == io_state_in_1 ? 8'h13 : _GEN_643; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_645 = 8'h85 == io_state_in_1 ? 8'h11 : _GEN_644; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_646 = 8'h86 == io_state_in_1 ? 8'h17 : _GEN_645; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_647 = 8'h87 == io_state_in_1 ? 8'h15 : _GEN_646; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_648 = 8'h88 == io_state_in_1 ? 8'hb : _GEN_647; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_649 = 8'h89 == io_state_in_1 ? 8'h9 : _GEN_648; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_650 = 8'h8a == io_state_in_1 ? 8'hf : _GEN_649; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_651 = 8'h8b == io_state_in_1 ? 8'hd : _GEN_650; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_652 = 8'h8c == io_state_in_1 ? 8'h3 : _GEN_651; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_653 = 8'h8d == io_state_in_1 ? 8'h1 : _GEN_652; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_654 = 8'h8e == io_state_in_1 ? 8'h7 : _GEN_653; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_655 = 8'h8f == io_state_in_1 ? 8'h5 : _GEN_654; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_656 = 8'h90 == io_state_in_1 ? 8'h3b : _GEN_655; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_657 = 8'h91 == io_state_in_1 ? 8'h39 : _GEN_656; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_658 = 8'h92 == io_state_in_1 ? 8'h3f : _GEN_657; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_659 = 8'h93 == io_state_in_1 ? 8'h3d : _GEN_658; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_660 = 8'h94 == io_state_in_1 ? 8'h33 : _GEN_659; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_661 = 8'h95 == io_state_in_1 ? 8'h31 : _GEN_660; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_662 = 8'h96 == io_state_in_1 ? 8'h37 : _GEN_661; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_663 = 8'h97 == io_state_in_1 ? 8'h35 : _GEN_662; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_664 = 8'h98 == io_state_in_1 ? 8'h2b : _GEN_663; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_665 = 8'h99 == io_state_in_1 ? 8'h29 : _GEN_664; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_666 = 8'h9a == io_state_in_1 ? 8'h2f : _GEN_665; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_667 = 8'h9b == io_state_in_1 ? 8'h2d : _GEN_666; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_668 = 8'h9c == io_state_in_1 ? 8'h23 : _GEN_667; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_669 = 8'h9d == io_state_in_1 ? 8'h21 : _GEN_668; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_670 = 8'h9e == io_state_in_1 ? 8'h27 : _GEN_669; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_671 = 8'h9f == io_state_in_1 ? 8'h25 : _GEN_670; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_672 = 8'ha0 == io_state_in_1 ? 8'h5b : _GEN_671; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_673 = 8'ha1 == io_state_in_1 ? 8'h59 : _GEN_672; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_674 = 8'ha2 == io_state_in_1 ? 8'h5f : _GEN_673; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_675 = 8'ha3 == io_state_in_1 ? 8'h5d : _GEN_674; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_676 = 8'ha4 == io_state_in_1 ? 8'h53 : _GEN_675; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_677 = 8'ha5 == io_state_in_1 ? 8'h51 : _GEN_676; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_678 = 8'ha6 == io_state_in_1 ? 8'h57 : _GEN_677; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_679 = 8'ha7 == io_state_in_1 ? 8'h55 : _GEN_678; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_680 = 8'ha8 == io_state_in_1 ? 8'h4b : _GEN_679; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_681 = 8'ha9 == io_state_in_1 ? 8'h49 : _GEN_680; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_682 = 8'haa == io_state_in_1 ? 8'h4f : _GEN_681; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_683 = 8'hab == io_state_in_1 ? 8'h4d : _GEN_682; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_684 = 8'hac == io_state_in_1 ? 8'h43 : _GEN_683; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_685 = 8'had == io_state_in_1 ? 8'h41 : _GEN_684; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_686 = 8'hae == io_state_in_1 ? 8'h47 : _GEN_685; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_687 = 8'haf == io_state_in_1 ? 8'h45 : _GEN_686; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_688 = 8'hb0 == io_state_in_1 ? 8'h7b : _GEN_687; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_689 = 8'hb1 == io_state_in_1 ? 8'h79 : _GEN_688; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_690 = 8'hb2 == io_state_in_1 ? 8'h7f : _GEN_689; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_691 = 8'hb3 == io_state_in_1 ? 8'h7d : _GEN_690; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_692 = 8'hb4 == io_state_in_1 ? 8'h73 : _GEN_691; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_693 = 8'hb5 == io_state_in_1 ? 8'h71 : _GEN_692; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_694 = 8'hb6 == io_state_in_1 ? 8'h77 : _GEN_693; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_695 = 8'hb7 == io_state_in_1 ? 8'h75 : _GEN_694; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_696 = 8'hb8 == io_state_in_1 ? 8'h6b : _GEN_695; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_697 = 8'hb9 == io_state_in_1 ? 8'h69 : _GEN_696; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_698 = 8'hba == io_state_in_1 ? 8'h6f : _GEN_697; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_699 = 8'hbb == io_state_in_1 ? 8'h6d : _GEN_698; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_700 = 8'hbc == io_state_in_1 ? 8'h63 : _GEN_699; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_701 = 8'hbd == io_state_in_1 ? 8'h61 : _GEN_700; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_702 = 8'hbe == io_state_in_1 ? 8'h67 : _GEN_701; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_703 = 8'hbf == io_state_in_1 ? 8'h65 : _GEN_702; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_704 = 8'hc0 == io_state_in_1 ? 8'h9b : _GEN_703; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_705 = 8'hc1 == io_state_in_1 ? 8'h99 : _GEN_704; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_706 = 8'hc2 == io_state_in_1 ? 8'h9f : _GEN_705; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_707 = 8'hc3 == io_state_in_1 ? 8'h9d : _GEN_706; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_708 = 8'hc4 == io_state_in_1 ? 8'h93 : _GEN_707; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_709 = 8'hc5 == io_state_in_1 ? 8'h91 : _GEN_708; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_710 = 8'hc6 == io_state_in_1 ? 8'h97 : _GEN_709; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_711 = 8'hc7 == io_state_in_1 ? 8'h95 : _GEN_710; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_712 = 8'hc8 == io_state_in_1 ? 8'h8b : _GEN_711; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_713 = 8'hc9 == io_state_in_1 ? 8'h89 : _GEN_712; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_714 = 8'hca == io_state_in_1 ? 8'h8f : _GEN_713; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_715 = 8'hcb == io_state_in_1 ? 8'h8d : _GEN_714; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_716 = 8'hcc == io_state_in_1 ? 8'h83 : _GEN_715; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_717 = 8'hcd == io_state_in_1 ? 8'h81 : _GEN_716; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_718 = 8'hce == io_state_in_1 ? 8'h87 : _GEN_717; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_719 = 8'hcf == io_state_in_1 ? 8'h85 : _GEN_718; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_720 = 8'hd0 == io_state_in_1 ? 8'hbb : _GEN_719; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_721 = 8'hd1 == io_state_in_1 ? 8'hb9 : _GEN_720; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_722 = 8'hd2 == io_state_in_1 ? 8'hbf : _GEN_721; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_723 = 8'hd3 == io_state_in_1 ? 8'hbd : _GEN_722; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_724 = 8'hd4 == io_state_in_1 ? 8'hb3 : _GEN_723; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_725 = 8'hd5 == io_state_in_1 ? 8'hb1 : _GEN_724; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_726 = 8'hd6 == io_state_in_1 ? 8'hb7 : _GEN_725; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_727 = 8'hd7 == io_state_in_1 ? 8'hb5 : _GEN_726; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_728 = 8'hd8 == io_state_in_1 ? 8'hab : _GEN_727; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_729 = 8'hd9 == io_state_in_1 ? 8'ha9 : _GEN_728; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_730 = 8'hda == io_state_in_1 ? 8'haf : _GEN_729; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_731 = 8'hdb == io_state_in_1 ? 8'had : _GEN_730; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_732 = 8'hdc == io_state_in_1 ? 8'ha3 : _GEN_731; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_733 = 8'hdd == io_state_in_1 ? 8'ha1 : _GEN_732; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_734 = 8'hde == io_state_in_1 ? 8'ha7 : _GEN_733; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_735 = 8'hdf == io_state_in_1 ? 8'ha5 : _GEN_734; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_736 = 8'he0 == io_state_in_1 ? 8'hdb : _GEN_735; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_737 = 8'he1 == io_state_in_1 ? 8'hd9 : _GEN_736; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_738 = 8'he2 == io_state_in_1 ? 8'hdf : _GEN_737; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_739 = 8'he3 == io_state_in_1 ? 8'hdd : _GEN_738; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_740 = 8'he4 == io_state_in_1 ? 8'hd3 : _GEN_739; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_741 = 8'he5 == io_state_in_1 ? 8'hd1 : _GEN_740; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_742 = 8'he6 == io_state_in_1 ? 8'hd7 : _GEN_741; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_743 = 8'he7 == io_state_in_1 ? 8'hd5 : _GEN_742; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_744 = 8'he8 == io_state_in_1 ? 8'hcb : _GEN_743; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_745 = 8'he9 == io_state_in_1 ? 8'hc9 : _GEN_744; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_746 = 8'hea == io_state_in_1 ? 8'hcf : _GEN_745; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_747 = 8'heb == io_state_in_1 ? 8'hcd : _GEN_746; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_748 = 8'hec == io_state_in_1 ? 8'hc3 : _GEN_747; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_749 = 8'hed == io_state_in_1 ? 8'hc1 : _GEN_748; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_750 = 8'hee == io_state_in_1 ? 8'hc7 : _GEN_749; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_751 = 8'hef == io_state_in_1 ? 8'hc5 : _GEN_750; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_752 = 8'hf0 == io_state_in_1 ? 8'hfb : _GEN_751; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_753 = 8'hf1 == io_state_in_1 ? 8'hf9 : _GEN_752; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_754 = 8'hf2 == io_state_in_1 ? 8'hff : _GEN_753; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_755 = 8'hf3 == io_state_in_1 ? 8'hfd : _GEN_754; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_756 = 8'hf4 == io_state_in_1 ? 8'hf3 : _GEN_755; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_757 = 8'hf5 == io_state_in_1 ? 8'hf1 : _GEN_756; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_758 = 8'hf6 == io_state_in_1 ? 8'hf7 : _GEN_757; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_759 = 8'hf7 == io_state_in_1 ? 8'hf5 : _GEN_758; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_760 = 8'hf8 == io_state_in_1 ? 8'heb : _GEN_759; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_761 = 8'hf9 == io_state_in_1 ? 8'he9 : _GEN_760; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_762 = 8'hfa == io_state_in_1 ? 8'hef : _GEN_761; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_763 = 8'hfb == io_state_in_1 ? 8'hed : _GEN_762; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_764 = 8'hfc == io_state_in_1 ? 8'he3 : _GEN_763; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_765 = 8'hfd == io_state_in_1 ? 8'he1 : _GEN_764; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_766 = 8'hfe == io_state_in_1 ? 8'he7 : _GEN_765; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _GEN_767 = 8'hff == io_state_in_1 ? 8'he5 : _GEN_766; // @[MixColumns.scala 126:{34,34}]
  wire [7:0] _tmp_state_1_T = io_state_in_0 ^ _GEN_767; // @[MixColumns.scala 126:34]
  wire [7:0] _GEN_769 = 8'h1 == io_state_in_2 ? 8'h3 : 8'h0; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_770 = 8'h2 == io_state_in_2 ? 8'h6 : _GEN_769; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_771 = 8'h3 == io_state_in_2 ? 8'h5 : _GEN_770; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_772 = 8'h4 == io_state_in_2 ? 8'hc : _GEN_771; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_773 = 8'h5 == io_state_in_2 ? 8'hf : _GEN_772; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_774 = 8'h6 == io_state_in_2 ? 8'ha : _GEN_773; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_775 = 8'h7 == io_state_in_2 ? 8'h9 : _GEN_774; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_776 = 8'h8 == io_state_in_2 ? 8'h18 : _GEN_775; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_777 = 8'h9 == io_state_in_2 ? 8'h1b : _GEN_776; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_778 = 8'ha == io_state_in_2 ? 8'h1e : _GEN_777; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_779 = 8'hb == io_state_in_2 ? 8'h1d : _GEN_778; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_780 = 8'hc == io_state_in_2 ? 8'h14 : _GEN_779; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_781 = 8'hd == io_state_in_2 ? 8'h17 : _GEN_780; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_782 = 8'he == io_state_in_2 ? 8'h12 : _GEN_781; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_783 = 8'hf == io_state_in_2 ? 8'h11 : _GEN_782; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_784 = 8'h10 == io_state_in_2 ? 8'h30 : _GEN_783; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_785 = 8'h11 == io_state_in_2 ? 8'h33 : _GEN_784; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_786 = 8'h12 == io_state_in_2 ? 8'h36 : _GEN_785; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_787 = 8'h13 == io_state_in_2 ? 8'h35 : _GEN_786; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_788 = 8'h14 == io_state_in_2 ? 8'h3c : _GEN_787; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_789 = 8'h15 == io_state_in_2 ? 8'h3f : _GEN_788; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_790 = 8'h16 == io_state_in_2 ? 8'h3a : _GEN_789; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_791 = 8'h17 == io_state_in_2 ? 8'h39 : _GEN_790; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_792 = 8'h18 == io_state_in_2 ? 8'h28 : _GEN_791; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_793 = 8'h19 == io_state_in_2 ? 8'h2b : _GEN_792; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_794 = 8'h1a == io_state_in_2 ? 8'h2e : _GEN_793; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_795 = 8'h1b == io_state_in_2 ? 8'h2d : _GEN_794; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_796 = 8'h1c == io_state_in_2 ? 8'h24 : _GEN_795; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_797 = 8'h1d == io_state_in_2 ? 8'h27 : _GEN_796; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_798 = 8'h1e == io_state_in_2 ? 8'h22 : _GEN_797; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_799 = 8'h1f == io_state_in_2 ? 8'h21 : _GEN_798; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_800 = 8'h20 == io_state_in_2 ? 8'h60 : _GEN_799; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_801 = 8'h21 == io_state_in_2 ? 8'h63 : _GEN_800; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_802 = 8'h22 == io_state_in_2 ? 8'h66 : _GEN_801; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_803 = 8'h23 == io_state_in_2 ? 8'h65 : _GEN_802; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_804 = 8'h24 == io_state_in_2 ? 8'h6c : _GEN_803; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_805 = 8'h25 == io_state_in_2 ? 8'h6f : _GEN_804; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_806 = 8'h26 == io_state_in_2 ? 8'h6a : _GEN_805; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_807 = 8'h27 == io_state_in_2 ? 8'h69 : _GEN_806; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_808 = 8'h28 == io_state_in_2 ? 8'h78 : _GEN_807; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_809 = 8'h29 == io_state_in_2 ? 8'h7b : _GEN_808; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_810 = 8'h2a == io_state_in_2 ? 8'h7e : _GEN_809; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_811 = 8'h2b == io_state_in_2 ? 8'h7d : _GEN_810; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_812 = 8'h2c == io_state_in_2 ? 8'h74 : _GEN_811; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_813 = 8'h2d == io_state_in_2 ? 8'h77 : _GEN_812; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_814 = 8'h2e == io_state_in_2 ? 8'h72 : _GEN_813; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_815 = 8'h2f == io_state_in_2 ? 8'h71 : _GEN_814; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_816 = 8'h30 == io_state_in_2 ? 8'h50 : _GEN_815; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_817 = 8'h31 == io_state_in_2 ? 8'h53 : _GEN_816; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_818 = 8'h32 == io_state_in_2 ? 8'h56 : _GEN_817; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_819 = 8'h33 == io_state_in_2 ? 8'h55 : _GEN_818; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_820 = 8'h34 == io_state_in_2 ? 8'h5c : _GEN_819; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_821 = 8'h35 == io_state_in_2 ? 8'h5f : _GEN_820; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_822 = 8'h36 == io_state_in_2 ? 8'h5a : _GEN_821; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_823 = 8'h37 == io_state_in_2 ? 8'h59 : _GEN_822; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_824 = 8'h38 == io_state_in_2 ? 8'h48 : _GEN_823; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_825 = 8'h39 == io_state_in_2 ? 8'h4b : _GEN_824; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_826 = 8'h3a == io_state_in_2 ? 8'h4e : _GEN_825; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_827 = 8'h3b == io_state_in_2 ? 8'h4d : _GEN_826; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_828 = 8'h3c == io_state_in_2 ? 8'h44 : _GEN_827; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_829 = 8'h3d == io_state_in_2 ? 8'h47 : _GEN_828; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_830 = 8'h3e == io_state_in_2 ? 8'h42 : _GEN_829; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_831 = 8'h3f == io_state_in_2 ? 8'h41 : _GEN_830; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_832 = 8'h40 == io_state_in_2 ? 8'hc0 : _GEN_831; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_833 = 8'h41 == io_state_in_2 ? 8'hc3 : _GEN_832; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_834 = 8'h42 == io_state_in_2 ? 8'hc6 : _GEN_833; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_835 = 8'h43 == io_state_in_2 ? 8'hc5 : _GEN_834; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_836 = 8'h44 == io_state_in_2 ? 8'hcc : _GEN_835; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_837 = 8'h45 == io_state_in_2 ? 8'hcf : _GEN_836; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_838 = 8'h46 == io_state_in_2 ? 8'hca : _GEN_837; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_839 = 8'h47 == io_state_in_2 ? 8'hc9 : _GEN_838; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_840 = 8'h48 == io_state_in_2 ? 8'hd8 : _GEN_839; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_841 = 8'h49 == io_state_in_2 ? 8'hdb : _GEN_840; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_842 = 8'h4a == io_state_in_2 ? 8'hde : _GEN_841; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_843 = 8'h4b == io_state_in_2 ? 8'hdd : _GEN_842; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_844 = 8'h4c == io_state_in_2 ? 8'hd4 : _GEN_843; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_845 = 8'h4d == io_state_in_2 ? 8'hd7 : _GEN_844; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_846 = 8'h4e == io_state_in_2 ? 8'hd2 : _GEN_845; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_847 = 8'h4f == io_state_in_2 ? 8'hd1 : _GEN_846; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_848 = 8'h50 == io_state_in_2 ? 8'hf0 : _GEN_847; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_849 = 8'h51 == io_state_in_2 ? 8'hf3 : _GEN_848; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_850 = 8'h52 == io_state_in_2 ? 8'hf6 : _GEN_849; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_851 = 8'h53 == io_state_in_2 ? 8'hf5 : _GEN_850; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_852 = 8'h54 == io_state_in_2 ? 8'hfc : _GEN_851; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_853 = 8'h55 == io_state_in_2 ? 8'hff : _GEN_852; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_854 = 8'h56 == io_state_in_2 ? 8'hfa : _GEN_853; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_855 = 8'h57 == io_state_in_2 ? 8'hf9 : _GEN_854; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_856 = 8'h58 == io_state_in_2 ? 8'he8 : _GEN_855; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_857 = 8'h59 == io_state_in_2 ? 8'heb : _GEN_856; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_858 = 8'h5a == io_state_in_2 ? 8'hee : _GEN_857; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_859 = 8'h5b == io_state_in_2 ? 8'hed : _GEN_858; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_860 = 8'h5c == io_state_in_2 ? 8'he4 : _GEN_859; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_861 = 8'h5d == io_state_in_2 ? 8'he7 : _GEN_860; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_862 = 8'h5e == io_state_in_2 ? 8'he2 : _GEN_861; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_863 = 8'h5f == io_state_in_2 ? 8'he1 : _GEN_862; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_864 = 8'h60 == io_state_in_2 ? 8'ha0 : _GEN_863; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_865 = 8'h61 == io_state_in_2 ? 8'ha3 : _GEN_864; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_866 = 8'h62 == io_state_in_2 ? 8'ha6 : _GEN_865; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_867 = 8'h63 == io_state_in_2 ? 8'ha5 : _GEN_866; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_868 = 8'h64 == io_state_in_2 ? 8'hac : _GEN_867; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_869 = 8'h65 == io_state_in_2 ? 8'haf : _GEN_868; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_870 = 8'h66 == io_state_in_2 ? 8'haa : _GEN_869; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_871 = 8'h67 == io_state_in_2 ? 8'ha9 : _GEN_870; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_872 = 8'h68 == io_state_in_2 ? 8'hb8 : _GEN_871; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_873 = 8'h69 == io_state_in_2 ? 8'hbb : _GEN_872; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_874 = 8'h6a == io_state_in_2 ? 8'hbe : _GEN_873; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_875 = 8'h6b == io_state_in_2 ? 8'hbd : _GEN_874; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_876 = 8'h6c == io_state_in_2 ? 8'hb4 : _GEN_875; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_877 = 8'h6d == io_state_in_2 ? 8'hb7 : _GEN_876; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_878 = 8'h6e == io_state_in_2 ? 8'hb2 : _GEN_877; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_879 = 8'h6f == io_state_in_2 ? 8'hb1 : _GEN_878; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_880 = 8'h70 == io_state_in_2 ? 8'h90 : _GEN_879; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_881 = 8'h71 == io_state_in_2 ? 8'h93 : _GEN_880; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_882 = 8'h72 == io_state_in_2 ? 8'h96 : _GEN_881; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_883 = 8'h73 == io_state_in_2 ? 8'h95 : _GEN_882; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_884 = 8'h74 == io_state_in_2 ? 8'h9c : _GEN_883; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_885 = 8'h75 == io_state_in_2 ? 8'h9f : _GEN_884; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_886 = 8'h76 == io_state_in_2 ? 8'h9a : _GEN_885; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_887 = 8'h77 == io_state_in_2 ? 8'h99 : _GEN_886; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_888 = 8'h78 == io_state_in_2 ? 8'h88 : _GEN_887; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_889 = 8'h79 == io_state_in_2 ? 8'h8b : _GEN_888; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_890 = 8'h7a == io_state_in_2 ? 8'h8e : _GEN_889; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_891 = 8'h7b == io_state_in_2 ? 8'h8d : _GEN_890; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_892 = 8'h7c == io_state_in_2 ? 8'h84 : _GEN_891; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_893 = 8'h7d == io_state_in_2 ? 8'h87 : _GEN_892; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_894 = 8'h7e == io_state_in_2 ? 8'h82 : _GEN_893; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_895 = 8'h7f == io_state_in_2 ? 8'h81 : _GEN_894; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_896 = 8'h80 == io_state_in_2 ? 8'h9b : _GEN_895; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_897 = 8'h81 == io_state_in_2 ? 8'h98 : _GEN_896; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_898 = 8'h82 == io_state_in_2 ? 8'h9d : _GEN_897; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_899 = 8'h83 == io_state_in_2 ? 8'h9e : _GEN_898; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_900 = 8'h84 == io_state_in_2 ? 8'h97 : _GEN_899; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_901 = 8'h85 == io_state_in_2 ? 8'h94 : _GEN_900; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_902 = 8'h86 == io_state_in_2 ? 8'h91 : _GEN_901; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_903 = 8'h87 == io_state_in_2 ? 8'h92 : _GEN_902; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_904 = 8'h88 == io_state_in_2 ? 8'h83 : _GEN_903; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_905 = 8'h89 == io_state_in_2 ? 8'h80 : _GEN_904; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_906 = 8'h8a == io_state_in_2 ? 8'h85 : _GEN_905; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_907 = 8'h8b == io_state_in_2 ? 8'h86 : _GEN_906; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_908 = 8'h8c == io_state_in_2 ? 8'h8f : _GEN_907; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_909 = 8'h8d == io_state_in_2 ? 8'h8c : _GEN_908; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_910 = 8'h8e == io_state_in_2 ? 8'h89 : _GEN_909; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_911 = 8'h8f == io_state_in_2 ? 8'h8a : _GEN_910; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_912 = 8'h90 == io_state_in_2 ? 8'hab : _GEN_911; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_913 = 8'h91 == io_state_in_2 ? 8'ha8 : _GEN_912; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_914 = 8'h92 == io_state_in_2 ? 8'had : _GEN_913; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_915 = 8'h93 == io_state_in_2 ? 8'hae : _GEN_914; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_916 = 8'h94 == io_state_in_2 ? 8'ha7 : _GEN_915; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_917 = 8'h95 == io_state_in_2 ? 8'ha4 : _GEN_916; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_918 = 8'h96 == io_state_in_2 ? 8'ha1 : _GEN_917; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_919 = 8'h97 == io_state_in_2 ? 8'ha2 : _GEN_918; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_920 = 8'h98 == io_state_in_2 ? 8'hb3 : _GEN_919; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_921 = 8'h99 == io_state_in_2 ? 8'hb0 : _GEN_920; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_922 = 8'h9a == io_state_in_2 ? 8'hb5 : _GEN_921; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_923 = 8'h9b == io_state_in_2 ? 8'hb6 : _GEN_922; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_924 = 8'h9c == io_state_in_2 ? 8'hbf : _GEN_923; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_925 = 8'h9d == io_state_in_2 ? 8'hbc : _GEN_924; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_926 = 8'h9e == io_state_in_2 ? 8'hb9 : _GEN_925; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_927 = 8'h9f == io_state_in_2 ? 8'hba : _GEN_926; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_928 = 8'ha0 == io_state_in_2 ? 8'hfb : _GEN_927; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_929 = 8'ha1 == io_state_in_2 ? 8'hf8 : _GEN_928; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_930 = 8'ha2 == io_state_in_2 ? 8'hfd : _GEN_929; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_931 = 8'ha3 == io_state_in_2 ? 8'hfe : _GEN_930; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_932 = 8'ha4 == io_state_in_2 ? 8'hf7 : _GEN_931; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_933 = 8'ha5 == io_state_in_2 ? 8'hf4 : _GEN_932; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_934 = 8'ha6 == io_state_in_2 ? 8'hf1 : _GEN_933; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_935 = 8'ha7 == io_state_in_2 ? 8'hf2 : _GEN_934; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_936 = 8'ha8 == io_state_in_2 ? 8'he3 : _GEN_935; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_937 = 8'ha9 == io_state_in_2 ? 8'he0 : _GEN_936; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_938 = 8'haa == io_state_in_2 ? 8'he5 : _GEN_937; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_939 = 8'hab == io_state_in_2 ? 8'he6 : _GEN_938; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_940 = 8'hac == io_state_in_2 ? 8'hef : _GEN_939; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_941 = 8'had == io_state_in_2 ? 8'hec : _GEN_940; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_942 = 8'hae == io_state_in_2 ? 8'he9 : _GEN_941; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_943 = 8'haf == io_state_in_2 ? 8'hea : _GEN_942; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_944 = 8'hb0 == io_state_in_2 ? 8'hcb : _GEN_943; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_945 = 8'hb1 == io_state_in_2 ? 8'hc8 : _GEN_944; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_946 = 8'hb2 == io_state_in_2 ? 8'hcd : _GEN_945; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_947 = 8'hb3 == io_state_in_2 ? 8'hce : _GEN_946; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_948 = 8'hb4 == io_state_in_2 ? 8'hc7 : _GEN_947; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_949 = 8'hb5 == io_state_in_2 ? 8'hc4 : _GEN_948; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_950 = 8'hb6 == io_state_in_2 ? 8'hc1 : _GEN_949; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_951 = 8'hb7 == io_state_in_2 ? 8'hc2 : _GEN_950; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_952 = 8'hb8 == io_state_in_2 ? 8'hd3 : _GEN_951; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_953 = 8'hb9 == io_state_in_2 ? 8'hd0 : _GEN_952; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_954 = 8'hba == io_state_in_2 ? 8'hd5 : _GEN_953; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_955 = 8'hbb == io_state_in_2 ? 8'hd6 : _GEN_954; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_956 = 8'hbc == io_state_in_2 ? 8'hdf : _GEN_955; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_957 = 8'hbd == io_state_in_2 ? 8'hdc : _GEN_956; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_958 = 8'hbe == io_state_in_2 ? 8'hd9 : _GEN_957; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_959 = 8'hbf == io_state_in_2 ? 8'hda : _GEN_958; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_960 = 8'hc0 == io_state_in_2 ? 8'h5b : _GEN_959; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_961 = 8'hc1 == io_state_in_2 ? 8'h58 : _GEN_960; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_962 = 8'hc2 == io_state_in_2 ? 8'h5d : _GEN_961; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_963 = 8'hc3 == io_state_in_2 ? 8'h5e : _GEN_962; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_964 = 8'hc4 == io_state_in_2 ? 8'h57 : _GEN_963; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_965 = 8'hc5 == io_state_in_2 ? 8'h54 : _GEN_964; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_966 = 8'hc6 == io_state_in_2 ? 8'h51 : _GEN_965; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_967 = 8'hc7 == io_state_in_2 ? 8'h52 : _GEN_966; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_968 = 8'hc8 == io_state_in_2 ? 8'h43 : _GEN_967; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_969 = 8'hc9 == io_state_in_2 ? 8'h40 : _GEN_968; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_970 = 8'hca == io_state_in_2 ? 8'h45 : _GEN_969; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_971 = 8'hcb == io_state_in_2 ? 8'h46 : _GEN_970; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_972 = 8'hcc == io_state_in_2 ? 8'h4f : _GEN_971; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_973 = 8'hcd == io_state_in_2 ? 8'h4c : _GEN_972; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_974 = 8'hce == io_state_in_2 ? 8'h49 : _GEN_973; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_975 = 8'hcf == io_state_in_2 ? 8'h4a : _GEN_974; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_976 = 8'hd0 == io_state_in_2 ? 8'h6b : _GEN_975; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_977 = 8'hd1 == io_state_in_2 ? 8'h68 : _GEN_976; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_978 = 8'hd2 == io_state_in_2 ? 8'h6d : _GEN_977; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_979 = 8'hd3 == io_state_in_2 ? 8'h6e : _GEN_978; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_980 = 8'hd4 == io_state_in_2 ? 8'h67 : _GEN_979; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_981 = 8'hd5 == io_state_in_2 ? 8'h64 : _GEN_980; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_982 = 8'hd6 == io_state_in_2 ? 8'h61 : _GEN_981; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_983 = 8'hd7 == io_state_in_2 ? 8'h62 : _GEN_982; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_984 = 8'hd8 == io_state_in_2 ? 8'h73 : _GEN_983; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_985 = 8'hd9 == io_state_in_2 ? 8'h70 : _GEN_984; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_986 = 8'hda == io_state_in_2 ? 8'h75 : _GEN_985; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_987 = 8'hdb == io_state_in_2 ? 8'h76 : _GEN_986; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_988 = 8'hdc == io_state_in_2 ? 8'h7f : _GEN_987; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_989 = 8'hdd == io_state_in_2 ? 8'h7c : _GEN_988; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_990 = 8'hde == io_state_in_2 ? 8'h79 : _GEN_989; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_991 = 8'hdf == io_state_in_2 ? 8'h7a : _GEN_990; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_992 = 8'he0 == io_state_in_2 ? 8'h3b : _GEN_991; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_993 = 8'he1 == io_state_in_2 ? 8'h38 : _GEN_992; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_994 = 8'he2 == io_state_in_2 ? 8'h3d : _GEN_993; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_995 = 8'he3 == io_state_in_2 ? 8'h3e : _GEN_994; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_996 = 8'he4 == io_state_in_2 ? 8'h37 : _GEN_995; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_997 = 8'he5 == io_state_in_2 ? 8'h34 : _GEN_996; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_998 = 8'he6 == io_state_in_2 ? 8'h31 : _GEN_997; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_999 = 8'he7 == io_state_in_2 ? 8'h32 : _GEN_998; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1000 = 8'he8 == io_state_in_2 ? 8'h23 : _GEN_999; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1001 = 8'he9 == io_state_in_2 ? 8'h20 : _GEN_1000; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1002 = 8'hea == io_state_in_2 ? 8'h25 : _GEN_1001; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1003 = 8'heb == io_state_in_2 ? 8'h26 : _GEN_1002; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1004 = 8'hec == io_state_in_2 ? 8'h2f : _GEN_1003; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1005 = 8'hed == io_state_in_2 ? 8'h2c : _GEN_1004; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1006 = 8'hee == io_state_in_2 ? 8'h29 : _GEN_1005; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1007 = 8'hef == io_state_in_2 ? 8'h2a : _GEN_1006; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1008 = 8'hf0 == io_state_in_2 ? 8'hb : _GEN_1007; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1009 = 8'hf1 == io_state_in_2 ? 8'h8 : _GEN_1008; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1010 = 8'hf2 == io_state_in_2 ? 8'hd : _GEN_1009; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1011 = 8'hf3 == io_state_in_2 ? 8'he : _GEN_1010; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1012 = 8'hf4 == io_state_in_2 ? 8'h7 : _GEN_1011; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1013 = 8'hf5 == io_state_in_2 ? 8'h4 : _GEN_1012; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1014 = 8'hf6 == io_state_in_2 ? 8'h1 : _GEN_1013; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1015 = 8'hf7 == io_state_in_2 ? 8'h2 : _GEN_1014; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1016 = 8'hf8 == io_state_in_2 ? 8'h13 : _GEN_1015; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1017 = 8'hf9 == io_state_in_2 ? 8'h10 : _GEN_1016; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1018 = 8'hfa == io_state_in_2 ? 8'h15 : _GEN_1017; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1019 = 8'hfb == io_state_in_2 ? 8'h16 : _GEN_1018; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1020 = 8'hfc == io_state_in_2 ? 8'h1f : _GEN_1019; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1021 = 8'hfd == io_state_in_2 ? 8'h1c : _GEN_1020; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1022 = 8'hfe == io_state_in_2 ? 8'h19 : _GEN_1021; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _GEN_1023 = 8'hff == io_state_in_2 ? 8'h1a : _GEN_1022; // @[MixColumns.scala 126:{58,58}]
  wire [7:0] _tmp_state_1_T_1 = _tmp_state_1_T ^ _GEN_1023; // @[MixColumns.scala 126:58]
  wire [7:0] _tmp_state_2_T = io_state_in_0 ^ io_state_in_1; // @[MixColumns.scala 127:34]
  wire [7:0] _GEN_1025 = 8'h1 == io_state_in_2 ? 8'h2 : 8'h0; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1026 = 8'h2 == io_state_in_2 ? 8'h4 : _GEN_1025; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1027 = 8'h3 == io_state_in_2 ? 8'h6 : _GEN_1026; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1028 = 8'h4 == io_state_in_2 ? 8'h8 : _GEN_1027; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1029 = 8'h5 == io_state_in_2 ? 8'ha : _GEN_1028; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1030 = 8'h6 == io_state_in_2 ? 8'hc : _GEN_1029; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1031 = 8'h7 == io_state_in_2 ? 8'he : _GEN_1030; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1032 = 8'h8 == io_state_in_2 ? 8'h10 : _GEN_1031; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1033 = 8'h9 == io_state_in_2 ? 8'h12 : _GEN_1032; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1034 = 8'ha == io_state_in_2 ? 8'h14 : _GEN_1033; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1035 = 8'hb == io_state_in_2 ? 8'h16 : _GEN_1034; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1036 = 8'hc == io_state_in_2 ? 8'h18 : _GEN_1035; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1037 = 8'hd == io_state_in_2 ? 8'h1a : _GEN_1036; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1038 = 8'he == io_state_in_2 ? 8'h1c : _GEN_1037; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1039 = 8'hf == io_state_in_2 ? 8'h1e : _GEN_1038; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1040 = 8'h10 == io_state_in_2 ? 8'h20 : _GEN_1039; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1041 = 8'h11 == io_state_in_2 ? 8'h22 : _GEN_1040; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1042 = 8'h12 == io_state_in_2 ? 8'h24 : _GEN_1041; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1043 = 8'h13 == io_state_in_2 ? 8'h26 : _GEN_1042; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1044 = 8'h14 == io_state_in_2 ? 8'h28 : _GEN_1043; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1045 = 8'h15 == io_state_in_2 ? 8'h2a : _GEN_1044; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1046 = 8'h16 == io_state_in_2 ? 8'h2c : _GEN_1045; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1047 = 8'h17 == io_state_in_2 ? 8'h2e : _GEN_1046; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1048 = 8'h18 == io_state_in_2 ? 8'h30 : _GEN_1047; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1049 = 8'h19 == io_state_in_2 ? 8'h32 : _GEN_1048; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1050 = 8'h1a == io_state_in_2 ? 8'h34 : _GEN_1049; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1051 = 8'h1b == io_state_in_2 ? 8'h36 : _GEN_1050; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1052 = 8'h1c == io_state_in_2 ? 8'h38 : _GEN_1051; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1053 = 8'h1d == io_state_in_2 ? 8'h3a : _GEN_1052; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1054 = 8'h1e == io_state_in_2 ? 8'h3c : _GEN_1053; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1055 = 8'h1f == io_state_in_2 ? 8'h3e : _GEN_1054; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1056 = 8'h20 == io_state_in_2 ? 8'h40 : _GEN_1055; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1057 = 8'h21 == io_state_in_2 ? 8'h42 : _GEN_1056; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1058 = 8'h22 == io_state_in_2 ? 8'h44 : _GEN_1057; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1059 = 8'h23 == io_state_in_2 ? 8'h46 : _GEN_1058; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1060 = 8'h24 == io_state_in_2 ? 8'h48 : _GEN_1059; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1061 = 8'h25 == io_state_in_2 ? 8'h4a : _GEN_1060; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1062 = 8'h26 == io_state_in_2 ? 8'h4c : _GEN_1061; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1063 = 8'h27 == io_state_in_2 ? 8'h4e : _GEN_1062; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1064 = 8'h28 == io_state_in_2 ? 8'h50 : _GEN_1063; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1065 = 8'h29 == io_state_in_2 ? 8'h52 : _GEN_1064; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1066 = 8'h2a == io_state_in_2 ? 8'h54 : _GEN_1065; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1067 = 8'h2b == io_state_in_2 ? 8'h56 : _GEN_1066; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1068 = 8'h2c == io_state_in_2 ? 8'h58 : _GEN_1067; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1069 = 8'h2d == io_state_in_2 ? 8'h5a : _GEN_1068; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1070 = 8'h2e == io_state_in_2 ? 8'h5c : _GEN_1069; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1071 = 8'h2f == io_state_in_2 ? 8'h5e : _GEN_1070; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1072 = 8'h30 == io_state_in_2 ? 8'h60 : _GEN_1071; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1073 = 8'h31 == io_state_in_2 ? 8'h62 : _GEN_1072; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1074 = 8'h32 == io_state_in_2 ? 8'h64 : _GEN_1073; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1075 = 8'h33 == io_state_in_2 ? 8'h66 : _GEN_1074; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1076 = 8'h34 == io_state_in_2 ? 8'h68 : _GEN_1075; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1077 = 8'h35 == io_state_in_2 ? 8'h6a : _GEN_1076; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1078 = 8'h36 == io_state_in_2 ? 8'h6c : _GEN_1077; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1079 = 8'h37 == io_state_in_2 ? 8'h6e : _GEN_1078; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1080 = 8'h38 == io_state_in_2 ? 8'h70 : _GEN_1079; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1081 = 8'h39 == io_state_in_2 ? 8'h72 : _GEN_1080; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1082 = 8'h3a == io_state_in_2 ? 8'h74 : _GEN_1081; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1083 = 8'h3b == io_state_in_2 ? 8'h76 : _GEN_1082; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1084 = 8'h3c == io_state_in_2 ? 8'h78 : _GEN_1083; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1085 = 8'h3d == io_state_in_2 ? 8'h7a : _GEN_1084; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1086 = 8'h3e == io_state_in_2 ? 8'h7c : _GEN_1085; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1087 = 8'h3f == io_state_in_2 ? 8'h7e : _GEN_1086; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1088 = 8'h40 == io_state_in_2 ? 8'h80 : _GEN_1087; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1089 = 8'h41 == io_state_in_2 ? 8'h82 : _GEN_1088; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1090 = 8'h42 == io_state_in_2 ? 8'h84 : _GEN_1089; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1091 = 8'h43 == io_state_in_2 ? 8'h86 : _GEN_1090; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1092 = 8'h44 == io_state_in_2 ? 8'h88 : _GEN_1091; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1093 = 8'h45 == io_state_in_2 ? 8'h8a : _GEN_1092; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1094 = 8'h46 == io_state_in_2 ? 8'h8c : _GEN_1093; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1095 = 8'h47 == io_state_in_2 ? 8'h8e : _GEN_1094; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1096 = 8'h48 == io_state_in_2 ? 8'h90 : _GEN_1095; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1097 = 8'h49 == io_state_in_2 ? 8'h92 : _GEN_1096; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1098 = 8'h4a == io_state_in_2 ? 8'h94 : _GEN_1097; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1099 = 8'h4b == io_state_in_2 ? 8'h96 : _GEN_1098; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1100 = 8'h4c == io_state_in_2 ? 8'h98 : _GEN_1099; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1101 = 8'h4d == io_state_in_2 ? 8'h9a : _GEN_1100; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1102 = 8'h4e == io_state_in_2 ? 8'h9c : _GEN_1101; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1103 = 8'h4f == io_state_in_2 ? 8'h9e : _GEN_1102; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1104 = 8'h50 == io_state_in_2 ? 8'ha0 : _GEN_1103; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1105 = 8'h51 == io_state_in_2 ? 8'ha2 : _GEN_1104; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1106 = 8'h52 == io_state_in_2 ? 8'ha4 : _GEN_1105; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1107 = 8'h53 == io_state_in_2 ? 8'ha6 : _GEN_1106; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1108 = 8'h54 == io_state_in_2 ? 8'ha8 : _GEN_1107; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1109 = 8'h55 == io_state_in_2 ? 8'haa : _GEN_1108; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1110 = 8'h56 == io_state_in_2 ? 8'hac : _GEN_1109; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1111 = 8'h57 == io_state_in_2 ? 8'hae : _GEN_1110; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1112 = 8'h58 == io_state_in_2 ? 8'hb0 : _GEN_1111; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1113 = 8'h59 == io_state_in_2 ? 8'hb2 : _GEN_1112; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1114 = 8'h5a == io_state_in_2 ? 8'hb4 : _GEN_1113; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1115 = 8'h5b == io_state_in_2 ? 8'hb6 : _GEN_1114; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1116 = 8'h5c == io_state_in_2 ? 8'hb8 : _GEN_1115; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1117 = 8'h5d == io_state_in_2 ? 8'hba : _GEN_1116; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1118 = 8'h5e == io_state_in_2 ? 8'hbc : _GEN_1117; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1119 = 8'h5f == io_state_in_2 ? 8'hbe : _GEN_1118; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1120 = 8'h60 == io_state_in_2 ? 8'hc0 : _GEN_1119; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1121 = 8'h61 == io_state_in_2 ? 8'hc2 : _GEN_1120; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1122 = 8'h62 == io_state_in_2 ? 8'hc4 : _GEN_1121; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1123 = 8'h63 == io_state_in_2 ? 8'hc6 : _GEN_1122; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1124 = 8'h64 == io_state_in_2 ? 8'hc8 : _GEN_1123; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1125 = 8'h65 == io_state_in_2 ? 8'hca : _GEN_1124; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1126 = 8'h66 == io_state_in_2 ? 8'hcc : _GEN_1125; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1127 = 8'h67 == io_state_in_2 ? 8'hce : _GEN_1126; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1128 = 8'h68 == io_state_in_2 ? 8'hd0 : _GEN_1127; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1129 = 8'h69 == io_state_in_2 ? 8'hd2 : _GEN_1128; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1130 = 8'h6a == io_state_in_2 ? 8'hd4 : _GEN_1129; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1131 = 8'h6b == io_state_in_2 ? 8'hd6 : _GEN_1130; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1132 = 8'h6c == io_state_in_2 ? 8'hd8 : _GEN_1131; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1133 = 8'h6d == io_state_in_2 ? 8'hda : _GEN_1132; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1134 = 8'h6e == io_state_in_2 ? 8'hdc : _GEN_1133; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1135 = 8'h6f == io_state_in_2 ? 8'hde : _GEN_1134; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1136 = 8'h70 == io_state_in_2 ? 8'he0 : _GEN_1135; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1137 = 8'h71 == io_state_in_2 ? 8'he2 : _GEN_1136; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1138 = 8'h72 == io_state_in_2 ? 8'he4 : _GEN_1137; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1139 = 8'h73 == io_state_in_2 ? 8'he6 : _GEN_1138; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1140 = 8'h74 == io_state_in_2 ? 8'he8 : _GEN_1139; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1141 = 8'h75 == io_state_in_2 ? 8'hea : _GEN_1140; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1142 = 8'h76 == io_state_in_2 ? 8'hec : _GEN_1141; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1143 = 8'h77 == io_state_in_2 ? 8'hee : _GEN_1142; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1144 = 8'h78 == io_state_in_2 ? 8'hf0 : _GEN_1143; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1145 = 8'h79 == io_state_in_2 ? 8'hf2 : _GEN_1144; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1146 = 8'h7a == io_state_in_2 ? 8'hf4 : _GEN_1145; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1147 = 8'h7b == io_state_in_2 ? 8'hf6 : _GEN_1146; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1148 = 8'h7c == io_state_in_2 ? 8'hf8 : _GEN_1147; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1149 = 8'h7d == io_state_in_2 ? 8'hfa : _GEN_1148; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1150 = 8'h7e == io_state_in_2 ? 8'hfc : _GEN_1149; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1151 = 8'h7f == io_state_in_2 ? 8'hfe : _GEN_1150; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1152 = 8'h80 == io_state_in_2 ? 8'h1b : _GEN_1151; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1153 = 8'h81 == io_state_in_2 ? 8'h19 : _GEN_1152; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1154 = 8'h82 == io_state_in_2 ? 8'h1f : _GEN_1153; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1155 = 8'h83 == io_state_in_2 ? 8'h1d : _GEN_1154; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1156 = 8'h84 == io_state_in_2 ? 8'h13 : _GEN_1155; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1157 = 8'h85 == io_state_in_2 ? 8'h11 : _GEN_1156; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1158 = 8'h86 == io_state_in_2 ? 8'h17 : _GEN_1157; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1159 = 8'h87 == io_state_in_2 ? 8'h15 : _GEN_1158; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1160 = 8'h88 == io_state_in_2 ? 8'hb : _GEN_1159; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1161 = 8'h89 == io_state_in_2 ? 8'h9 : _GEN_1160; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1162 = 8'h8a == io_state_in_2 ? 8'hf : _GEN_1161; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1163 = 8'h8b == io_state_in_2 ? 8'hd : _GEN_1162; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1164 = 8'h8c == io_state_in_2 ? 8'h3 : _GEN_1163; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1165 = 8'h8d == io_state_in_2 ? 8'h1 : _GEN_1164; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1166 = 8'h8e == io_state_in_2 ? 8'h7 : _GEN_1165; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1167 = 8'h8f == io_state_in_2 ? 8'h5 : _GEN_1166; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1168 = 8'h90 == io_state_in_2 ? 8'h3b : _GEN_1167; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1169 = 8'h91 == io_state_in_2 ? 8'h39 : _GEN_1168; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1170 = 8'h92 == io_state_in_2 ? 8'h3f : _GEN_1169; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1171 = 8'h93 == io_state_in_2 ? 8'h3d : _GEN_1170; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1172 = 8'h94 == io_state_in_2 ? 8'h33 : _GEN_1171; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1173 = 8'h95 == io_state_in_2 ? 8'h31 : _GEN_1172; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1174 = 8'h96 == io_state_in_2 ? 8'h37 : _GEN_1173; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1175 = 8'h97 == io_state_in_2 ? 8'h35 : _GEN_1174; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1176 = 8'h98 == io_state_in_2 ? 8'h2b : _GEN_1175; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1177 = 8'h99 == io_state_in_2 ? 8'h29 : _GEN_1176; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1178 = 8'h9a == io_state_in_2 ? 8'h2f : _GEN_1177; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1179 = 8'h9b == io_state_in_2 ? 8'h2d : _GEN_1178; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1180 = 8'h9c == io_state_in_2 ? 8'h23 : _GEN_1179; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1181 = 8'h9d == io_state_in_2 ? 8'h21 : _GEN_1180; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1182 = 8'h9e == io_state_in_2 ? 8'h27 : _GEN_1181; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1183 = 8'h9f == io_state_in_2 ? 8'h25 : _GEN_1182; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1184 = 8'ha0 == io_state_in_2 ? 8'h5b : _GEN_1183; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1185 = 8'ha1 == io_state_in_2 ? 8'h59 : _GEN_1184; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1186 = 8'ha2 == io_state_in_2 ? 8'h5f : _GEN_1185; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1187 = 8'ha3 == io_state_in_2 ? 8'h5d : _GEN_1186; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1188 = 8'ha4 == io_state_in_2 ? 8'h53 : _GEN_1187; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1189 = 8'ha5 == io_state_in_2 ? 8'h51 : _GEN_1188; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1190 = 8'ha6 == io_state_in_2 ? 8'h57 : _GEN_1189; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1191 = 8'ha7 == io_state_in_2 ? 8'h55 : _GEN_1190; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1192 = 8'ha8 == io_state_in_2 ? 8'h4b : _GEN_1191; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1193 = 8'ha9 == io_state_in_2 ? 8'h49 : _GEN_1192; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1194 = 8'haa == io_state_in_2 ? 8'h4f : _GEN_1193; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1195 = 8'hab == io_state_in_2 ? 8'h4d : _GEN_1194; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1196 = 8'hac == io_state_in_2 ? 8'h43 : _GEN_1195; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1197 = 8'had == io_state_in_2 ? 8'h41 : _GEN_1196; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1198 = 8'hae == io_state_in_2 ? 8'h47 : _GEN_1197; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1199 = 8'haf == io_state_in_2 ? 8'h45 : _GEN_1198; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1200 = 8'hb0 == io_state_in_2 ? 8'h7b : _GEN_1199; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1201 = 8'hb1 == io_state_in_2 ? 8'h79 : _GEN_1200; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1202 = 8'hb2 == io_state_in_2 ? 8'h7f : _GEN_1201; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1203 = 8'hb3 == io_state_in_2 ? 8'h7d : _GEN_1202; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1204 = 8'hb4 == io_state_in_2 ? 8'h73 : _GEN_1203; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1205 = 8'hb5 == io_state_in_2 ? 8'h71 : _GEN_1204; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1206 = 8'hb6 == io_state_in_2 ? 8'h77 : _GEN_1205; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1207 = 8'hb7 == io_state_in_2 ? 8'h75 : _GEN_1206; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1208 = 8'hb8 == io_state_in_2 ? 8'h6b : _GEN_1207; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1209 = 8'hb9 == io_state_in_2 ? 8'h69 : _GEN_1208; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1210 = 8'hba == io_state_in_2 ? 8'h6f : _GEN_1209; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1211 = 8'hbb == io_state_in_2 ? 8'h6d : _GEN_1210; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1212 = 8'hbc == io_state_in_2 ? 8'h63 : _GEN_1211; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1213 = 8'hbd == io_state_in_2 ? 8'h61 : _GEN_1212; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1214 = 8'hbe == io_state_in_2 ? 8'h67 : _GEN_1213; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1215 = 8'hbf == io_state_in_2 ? 8'h65 : _GEN_1214; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1216 = 8'hc0 == io_state_in_2 ? 8'h9b : _GEN_1215; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1217 = 8'hc1 == io_state_in_2 ? 8'h99 : _GEN_1216; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1218 = 8'hc2 == io_state_in_2 ? 8'h9f : _GEN_1217; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1219 = 8'hc3 == io_state_in_2 ? 8'h9d : _GEN_1218; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1220 = 8'hc4 == io_state_in_2 ? 8'h93 : _GEN_1219; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1221 = 8'hc5 == io_state_in_2 ? 8'h91 : _GEN_1220; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1222 = 8'hc6 == io_state_in_2 ? 8'h97 : _GEN_1221; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1223 = 8'hc7 == io_state_in_2 ? 8'h95 : _GEN_1222; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1224 = 8'hc8 == io_state_in_2 ? 8'h8b : _GEN_1223; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1225 = 8'hc9 == io_state_in_2 ? 8'h89 : _GEN_1224; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1226 = 8'hca == io_state_in_2 ? 8'h8f : _GEN_1225; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1227 = 8'hcb == io_state_in_2 ? 8'h8d : _GEN_1226; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1228 = 8'hcc == io_state_in_2 ? 8'h83 : _GEN_1227; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1229 = 8'hcd == io_state_in_2 ? 8'h81 : _GEN_1228; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1230 = 8'hce == io_state_in_2 ? 8'h87 : _GEN_1229; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1231 = 8'hcf == io_state_in_2 ? 8'h85 : _GEN_1230; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1232 = 8'hd0 == io_state_in_2 ? 8'hbb : _GEN_1231; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1233 = 8'hd1 == io_state_in_2 ? 8'hb9 : _GEN_1232; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1234 = 8'hd2 == io_state_in_2 ? 8'hbf : _GEN_1233; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1235 = 8'hd3 == io_state_in_2 ? 8'hbd : _GEN_1234; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1236 = 8'hd4 == io_state_in_2 ? 8'hb3 : _GEN_1235; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1237 = 8'hd5 == io_state_in_2 ? 8'hb1 : _GEN_1236; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1238 = 8'hd6 == io_state_in_2 ? 8'hb7 : _GEN_1237; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1239 = 8'hd7 == io_state_in_2 ? 8'hb5 : _GEN_1238; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1240 = 8'hd8 == io_state_in_2 ? 8'hab : _GEN_1239; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1241 = 8'hd9 == io_state_in_2 ? 8'ha9 : _GEN_1240; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1242 = 8'hda == io_state_in_2 ? 8'haf : _GEN_1241; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1243 = 8'hdb == io_state_in_2 ? 8'had : _GEN_1242; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1244 = 8'hdc == io_state_in_2 ? 8'ha3 : _GEN_1243; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1245 = 8'hdd == io_state_in_2 ? 8'ha1 : _GEN_1244; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1246 = 8'hde == io_state_in_2 ? 8'ha7 : _GEN_1245; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1247 = 8'hdf == io_state_in_2 ? 8'ha5 : _GEN_1246; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1248 = 8'he0 == io_state_in_2 ? 8'hdb : _GEN_1247; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1249 = 8'he1 == io_state_in_2 ? 8'hd9 : _GEN_1248; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1250 = 8'he2 == io_state_in_2 ? 8'hdf : _GEN_1249; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1251 = 8'he3 == io_state_in_2 ? 8'hdd : _GEN_1250; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1252 = 8'he4 == io_state_in_2 ? 8'hd3 : _GEN_1251; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1253 = 8'he5 == io_state_in_2 ? 8'hd1 : _GEN_1252; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1254 = 8'he6 == io_state_in_2 ? 8'hd7 : _GEN_1253; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1255 = 8'he7 == io_state_in_2 ? 8'hd5 : _GEN_1254; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1256 = 8'he8 == io_state_in_2 ? 8'hcb : _GEN_1255; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1257 = 8'he9 == io_state_in_2 ? 8'hc9 : _GEN_1256; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1258 = 8'hea == io_state_in_2 ? 8'hcf : _GEN_1257; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1259 = 8'heb == io_state_in_2 ? 8'hcd : _GEN_1258; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1260 = 8'hec == io_state_in_2 ? 8'hc3 : _GEN_1259; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1261 = 8'hed == io_state_in_2 ? 8'hc1 : _GEN_1260; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1262 = 8'hee == io_state_in_2 ? 8'hc7 : _GEN_1261; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1263 = 8'hef == io_state_in_2 ? 8'hc5 : _GEN_1262; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1264 = 8'hf0 == io_state_in_2 ? 8'hfb : _GEN_1263; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1265 = 8'hf1 == io_state_in_2 ? 8'hf9 : _GEN_1264; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1266 = 8'hf2 == io_state_in_2 ? 8'hff : _GEN_1265; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1267 = 8'hf3 == io_state_in_2 ? 8'hfd : _GEN_1266; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1268 = 8'hf4 == io_state_in_2 ? 8'hf3 : _GEN_1267; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1269 = 8'hf5 == io_state_in_2 ? 8'hf1 : _GEN_1268; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1270 = 8'hf6 == io_state_in_2 ? 8'hf7 : _GEN_1269; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1271 = 8'hf7 == io_state_in_2 ? 8'hf5 : _GEN_1270; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1272 = 8'hf8 == io_state_in_2 ? 8'heb : _GEN_1271; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1273 = 8'hf9 == io_state_in_2 ? 8'he9 : _GEN_1272; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1274 = 8'hfa == io_state_in_2 ? 8'hef : _GEN_1273; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1275 = 8'hfb == io_state_in_2 ? 8'hed : _GEN_1274; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1276 = 8'hfc == io_state_in_2 ? 8'he3 : _GEN_1275; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1277 = 8'hfd == io_state_in_2 ? 8'he1 : _GEN_1276; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1278 = 8'hfe == io_state_in_2 ? 8'he7 : _GEN_1277; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _GEN_1279 = 8'hff == io_state_in_2 ? 8'he5 : _GEN_1278; // @[MixColumns.scala 127:{51,51}]
  wire [7:0] _tmp_state_2_T_1 = _tmp_state_2_T ^ _GEN_1279; // @[MixColumns.scala 127:51]
  wire [7:0] _GEN_1281 = 8'h1 == io_state_in_3 ? 8'h3 : 8'h0; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1282 = 8'h2 == io_state_in_3 ? 8'h6 : _GEN_1281; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1283 = 8'h3 == io_state_in_3 ? 8'h5 : _GEN_1282; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1284 = 8'h4 == io_state_in_3 ? 8'hc : _GEN_1283; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1285 = 8'h5 == io_state_in_3 ? 8'hf : _GEN_1284; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1286 = 8'h6 == io_state_in_3 ? 8'ha : _GEN_1285; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1287 = 8'h7 == io_state_in_3 ? 8'h9 : _GEN_1286; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1288 = 8'h8 == io_state_in_3 ? 8'h18 : _GEN_1287; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1289 = 8'h9 == io_state_in_3 ? 8'h1b : _GEN_1288; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1290 = 8'ha == io_state_in_3 ? 8'h1e : _GEN_1289; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1291 = 8'hb == io_state_in_3 ? 8'h1d : _GEN_1290; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1292 = 8'hc == io_state_in_3 ? 8'h14 : _GEN_1291; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1293 = 8'hd == io_state_in_3 ? 8'h17 : _GEN_1292; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1294 = 8'he == io_state_in_3 ? 8'h12 : _GEN_1293; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1295 = 8'hf == io_state_in_3 ? 8'h11 : _GEN_1294; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1296 = 8'h10 == io_state_in_3 ? 8'h30 : _GEN_1295; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1297 = 8'h11 == io_state_in_3 ? 8'h33 : _GEN_1296; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1298 = 8'h12 == io_state_in_3 ? 8'h36 : _GEN_1297; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1299 = 8'h13 == io_state_in_3 ? 8'h35 : _GEN_1298; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1300 = 8'h14 == io_state_in_3 ? 8'h3c : _GEN_1299; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1301 = 8'h15 == io_state_in_3 ? 8'h3f : _GEN_1300; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1302 = 8'h16 == io_state_in_3 ? 8'h3a : _GEN_1301; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1303 = 8'h17 == io_state_in_3 ? 8'h39 : _GEN_1302; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1304 = 8'h18 == io_state_in_3 ? 8'h28 : _GEN_1303; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1305 = 8'h19 == io_state_in_3 ? 8'h2b : _GEN_1304; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1306 = 8'h1a == io_state_in_3 ? 8'h2e : _GEN_1305; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1307 = 8'h1b == io_state_in_3 ? 8'h2d : _GEN_1306; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1308 = 8'h1c == io_state_in_3 ? 8'h24 : _GEN_1307; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1309 = 8'h1d == io_state_in_3 ? 8'h27 : _GEN_1308; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1310 = 8'h1e == io_state_in_3 ? 8'h22 : _GEN_1309; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1311 = 8'h1f == io_state_in_3 ? 8'h21 : _GEN_1310; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1312 = 8'h20 == io_state_in_3 ? 8'h60 : _GEN_1311; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1313 = 8'h21 == io_state_in_3 ? 8'h63 : _GEN_1312; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1314 = 8'h22 == io_state_in_3 ? 8'h66 : _GEN_1313; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1315 = 8'h23 == io_state_in_3 ? 8'h65 : _GEN_1314; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1316 = 8'h24 == io_state_in_3 ? 8'h6c : _GEN_1315; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1317 = 8'h25 == io_state_in_3 ? 8'h6f : _GEN_1316; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1318 = 8'h26 == io_state_in_3 ? 8'h6a : _GEN_1317; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1319 = 8'h27 == io_state_in_3 ? 8'h69 : _GEN_1318; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1320 = 8'h28 == io_state_in_3 ? 8'h78 : _GEN_1319; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1321 = 8'h29 == io_state_in_3 ? 8'h7b : _GEN_1320; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1322 = 8'h2a == io_state_in_3 ? 8'h7e : _GEN_1321; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1323 = 8'h2b == io_state_in_3 ? 8'h7d : _GEN_1322; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1324 = 8'h2c == io_state_in_3 ? 8'h74 : _GEN_1323; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1325 = 8'h2d == io_state_in_3 ? 8'h77 : _GEN_1324; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1326 = 8'h2e == io_state_in_3 ? 8'h72 : _GEN_1325; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1327 = 8'h2f == io_state_in_3 ? 8'h71 : _GEN_1326; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1328 = 8'h30 == io_state_in_3 ? 8'h50 : _GEN_1327; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1329 = 8'h31 == io_state_in_3 ? 8'h53 : _GEN_1328; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1330 = 8'h32 == io_state_in_3 ? 8'h56 : _GEN_1329; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1331 = 8'h33 == io_state_in_3 ? 8'h55 : _GEN_1330; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1332 = 8'h34 == io_state_in_3 ? 8'h5c : _GEN_1331; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1333 = 8'h35 == io_state_in_3 ? 8'h5f : _GEN_1332; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1334 = 8'h36 == io_state_in_3 ? 8'h5a : _GEN_1333; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1335 = 8'h37 == io_state_in_3 ? 8'h59 : _GEN_1334; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1336 = 8'h38 == io_state_in_3 ? 8'h48 : _GEN_1335; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1337 = 8'h39 == io_state_in_3 ? 8'h4b : _GEN_1336; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1338 = 8'h3a == io_state_in_3 ? 8'h4e : _GEN_1337; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1339 = 8'h3b == io_state_in_3 ? 8'h4d : _GEN_1338; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1340 = 8'h3c == io_state_in_3 ? 8'h44 : _GEN_1339; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1341 = 8'h3d == io_state_in_3 ? 8'h47 : _GEN_1340; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1342 = 8'h3e == io_state_in_3 ? 8'h42 : _GEN_1341; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1343 = 8'h3f == io_state_in_3 ? 8'h41 : _GEN_1342; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1344 = 8'h40 == io_state_in_3 ? 8'hc0 : _GEN_1343; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1345 = 8'h41 == io_state_in_3 ? 8'hc3 : _GEN_1344; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1346 = 8'h42 == io_state_in_3 ? 8'hc6 : _GEN_1345; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1347 = 8'h43 == io_state_in_3 ? 8'hc5 : _GEN_1346; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1348 = 8'h44 == io_state_in_3 ? 8'hcc : _GEN_1347; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1349 = 8'h45 == io_state_in_3 ? 8'hcf : _GEN_1348; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1350 = 8'h46 == io_state_in_3 ? 8'hca : _GEN_1349; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1351 = 8'h47 == io_state_in_3 ? 8'hc9 : _GEN_1350; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1352 = 8'h48 == io_state_in_3 ? 8'hd8 : _GEN_1351; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1353 = 8'h49 == io_state_in_3 ? 8'hdb : _GEN_1352; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1354 = 8'h4a == io_state_in_3 ? 8'hde : _GEN_1353; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1355 = 8'h4b == io_state_in_3 ? 8'hdd : _GEN_1354; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1356 = 8'h4c == io_state_in_3 ? 8'hd4 : _GEN_1355; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1357 = 8'h4d == io_state_in_3 ? 8'hd7 : _GEN_1356; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1358 = 8'h4e == io_state_in_3 ? 8'hd2 : _GEN_1357; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1359 = 8'h4f == io_state_in_3 ? 8'hd1 : _GEN_1358; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1360 = 8'h50 == io_state_in_3 ? 8'hf0 : _GEN_1359; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1361 = 8'h51 == io_state_in_3 ? 8'hf3 : _GEN_1360; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1362 = 8'h52 == io_state_in_3 ? 8'hf6 : _GEN_1361; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1363 = 8'h53 == io_state_in_3 ? 8'hf5 : _GEN_1362; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1364 = 8'h54 == io_state_in_3 ? 8'hfc : _GEN_1363; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1365 = 8'h55 == io_state_in_3 ? 8'hff : _GEN_1364; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1366 = 8'h56 == io_state_in_3 ? 8'hfa : _GEN_1365; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1367 = 8'h57 == io_state_in_3 ? 8'hf9 : _GEN_1366; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1368 = 8'h58 == io_state_in_3 ? 8'he8 : _GEN_1367; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1369 = 8'h59 == io_state_in_3 ? 8'heb : _GEN_1368; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1370 = 8'h5a == io_state_in_3 ? 8'hee : _GEN_1369; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1371 = 8'h5b == io_state_in_3 ? 8'hed : _GEN_1370; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1372 = 8'h5c == io_state_in_3 ? 8'he4 : _GEN_1371; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1373 = 8'h5d == io_state_in_3 ? 8'he7 : _GEN_1372; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1374 = 8'h5e == io_state_in_3 ? 8'he2 : _GEN_1373; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1375 = 8'h5f == io_state_in_3 ? 8'he1 : _GEN_1374; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1376 = 8'h60 == io_state_in_3 ? 8'ha0 : _GEN_1375; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1377 = 8'h61 == io_state_in_3 ? 8'ha3 : _GEN_1376; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1378 = 8'h62 == io_state_in_3 ? 8'ha6 : _GEN_1377; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1379 = 8'h63 == io_state_in_3 ? 8'ha5 : _GEN_1378; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1380 = 8'h64 == io_state_in_3 ? 8'hac : _GEN_1379; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1381 = 8'h65 == io_state_in_3 ? 8'haf : _GEN_1380; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1382 = 8'h66 == io_state_in_3 ? 8'haa : _GEN_1381; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1383 = 8'h67 == io_state_in_3 ? 8'ha9 : _GEN_1382; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1384 = 8'h68 == io_state_in_3 ? 8'hb8 : _GEN_1383; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1385 = 8'h69 == io_state_in_3 ? 8'hbb : _GEN_1384; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1386 = 8'h6a == io_state_in_3 ? 8'hbe : _GEN_1385; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1387 = 8'h6b == io_state_in_3 ? 8'hbd : _GEN_1386; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1388 = 8'h6c == io_state_in_3 ? 8'hb4 : _GEN_1387; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1389 = 8'h6d == io_state_in_3 ? 8'hb7 : _GEN_1388; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1390 = 8'h6e == io_state_in_3 ? 8'hb2 : _GEN_1389; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1391 = 8'h6f == io_state_in_3 ? 8'hb1 : _GEN_1390; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1392 = 8'h70 == io_state_in_3 ? 8'h90 : _GEN_1391; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1393 = 8'h71 == io_state_in_3 ? 8'h93 : _GEN_1392; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1394 = 8'h72 == io_state_in_3 ? 8'h96 : _GEN_1393; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1395 = 8'h73 == io_state_in_3 ? 8'h95 : _GEN_1394; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1396 = 8'h74 == io_state_in_3 ? 8'h9c : _GEN_1395; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1397 = 8'h75 == io_state_in_3 ? 8'h9f : _GEN_1396; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1398 = 8'h76 == io_state_in_3 ? 8'h9a : _GEN_1397; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1399 = 8'h77 == io_state_in_3 ? 8'h99 : _GEN_1398; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1400 = 8'h78 == io_state_in_3 ? 8'h88 : _GEN_1399; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1401 = 8'h79 == io_state_in_3 ? 8'h8b : _GEN_1400; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1402 = 8'h7a == io_state_in_3 ? 8'h8e : _GEN_1401; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1403 = 8'h7b == io_state_in_3 ? 8'h8d : _GEN_1402; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1404 = 8'h7c == io_state_in_3 ? 8'h84 : _GEN_1403; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1405 = 8'h7d == io_state_in_3 ? 8'h87 : _GEN_1404; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1406 = 8'h7e == io_state_in_3 ? 8'h82 : _GEN_1405; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1407 = 8'h7f == io_state_in_3 ? 8'h81 : _GEN_1406; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1408 = 8'h80 == io_state_in_3 ? 8'h9b : _GEN_1407; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1409 = 8'h81 == io_state_in_3 ? 8'h98 : _GEN_1408; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1410 = 8'h82 == io_state_in_3 ? 8'h9d : _GEN_1409; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1411 = 8'h83 == io_state_in_3 ? 8'h9e : _GEN_1410; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1412 = 8'h84 == io_state_in_3 ? 8'h97 : _GEN_1411; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1413 = 8'h85 == io_state_in_3 ? 8'h94 : _GEN_1412; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1414 = 8'h86 == io_state_in_3 ? 8'h91 : _GEN_1413; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1415 = 8'h87 == io_state_in_3 ? 8'h92 : _GEN_1414; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1416 = 8'h88 == io_state_in_3 ? 8'h83 : _GEN_1415; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1417 = 8'h89 == io_state_in_3 ? 8'h80 : _GEN_1416; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1418 = 8'h8a == io_state_in_3 ? 8'h85 : _GEN_1417; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1419 = 8'h8b == io_state_in_3 ? 8'h86 : _GEN_1418; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1420 = 8'h8c == io_state_in_3 ? 8'h8f : _GEN_1419; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1421 = 8'h8d == io_state_in_3 ? 8'h8c : _GEN_1420; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1422 = 8'h8e == io_state_in_3 ? 8'h89 : _GEN_1421; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1423 = 8'h8f == io_state_in_3 ? 8'h8a : _GEN_1422; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1424 = 8'h90 == io_state_in_3 ? 8'hab : _GEN_1423; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1425 = 8'h91 == io_state_in_3 ? 8'ha8 : _GEN_1424; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1426 = 8'h92 == io_state_in_3 ? 8'had : _GEN_1425; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1427 = 8'h93 == io_state_in_3 ? 8'hae : _GEN_1426; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1428 = 8'h94 == io_state_in_3 ? 8'ha7 : _GEN_1427; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1429 = 8'h95 == io_state_in_3 ? 8'ha4 : _GEN_1428; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1430 = 8'h96 == io_state_in_3 ? 8'ha1 : _GEN_1429; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1431 = 8'h97 == io_state_in_3 ? 8'ha2 : _GEN_1430; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1432 = 8'h98 == io_state_in_3 ? 8'hb3 : _GEN_1431; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1433 = 8'h99 == io_state_in_3 ? 8'hb0 : _GEN_1432; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1434 = 8'h9a == io_state_in_3 ? 8'hb5 : _GEN_1433; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1435 = 8'h9b == io_state_in_3 ? 8'hb6 : _GEN_1434; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1436 = 8'h9c == io_state_in_3 ? 8'hbf : _GEN_1435; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1437 = 8'h9d == io_state_in_3 ? 8'hbc : _GEN_1436; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1438 = 8'h9e == io_state_in_3 ? 8'hb9 : _GEN_1437; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1439 = 8'h9f == io_state_in_3 ? 8'hba : _GEN_1438; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1440 = 8'ha0 == io_state_in_3 ? 8'hfb : _GEN_1439; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1441 = 8'ha1 == io_state_in_3 ? 8'hf8 : _GEN_1440; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1442 = 8'ha2 == io_state_in_3 ? 8'hfd : _GEN_1441; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1443 = 8'ha3 == io_state_in_3 ? 8'hfe : _GEN_1442; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1444 = 8'ha4 == io_state_in_3 ? 8'hf7 : _GEN_1443; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1445 = 8'ha5 == io_state_in_3 ? 8'hf4 : _GEN_1444; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1446 = 8'ha6 == io_state_in_3 ? 8'hf1 : _GEN_1445; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1447 = 8'ha7 == io_state_in_3 ? 8'hf2 : _GEN_1446; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1448 = 8'ha8 == io_state_in_3 ? 8'he3 : _GEN_1447; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1449 = 8'ha9 == io_state_in_3 ? 8'he0 : _GEN_1448; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1450 = 8'haa == io_state_in_3 ? 8'he5 : _GEN_1449; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1451 = 8'hab == io_state_in_3 ? 8'he6 : _GEN_1450; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1452 = 8'hac == io_state_in_3 ? 8'hef : _GEN_1451; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1453 = 8'had == io_state_in_3 ? 8'hec : _GEN_1452; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1454 = 8'hae == io_state_in_3 ? 8'he9 : _GEN_1453; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1455 = 8'haf == io_state_in_3 ? 8'hea : _GEN_1454; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1456 = 8'hb0 == io_state_in_3 ? 8'hcb : _GEN_1455; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1457 = 8'hb1 == io_state_in_3 ? 8'hc8 : _GEN_1456; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1458 = 8'hb2 == io_state_in_3 ? 8'hcd : _GEN_1457; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1459 = 8'hb3 == io_state_in_3 ? 8'hce : _GEN_1458; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1460 = 8'hb4 == io_state_in_3 ? 8'hc7 : _GEN_1459; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1461 = 8'hb5 == io_state_in_3 ? 8'hc4 : _GEN_1460; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1462 = 8'hb6 == io_state_in_3 ? 8'hc1 : _GEN_1461; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1463 = 8'hb7 == io_state_in_3 ? 8'hc2 : _GEN_1462; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1464 = 8'hb8 == io_state_in_3 ? 8'hd3 : _GEN_1463; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1465 = 8'hb9 == io_state_in_3 ? 8'hd0 : _GEN_1464; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1466 = 8'hba == io_state_in_3 ? 8'hd5 : _GEN_1465; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1467 = 8'hbb == io_state_in_3 ? 8'hd6 : _GEN_1466; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1468 = 8'hbc == io_state_in_3 ? 8'hdf : _GEN_1467; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1469 = 8'hbd == io_state_in_3 ? 8'hdc : _GEN_1468; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1470 = 8'hbe == io_state_in_3 ? 8'hd9 : _GEN_1469; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1471 = 8'hbf == io_state_in_3 ? 8'hda : _GEN_1470; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1472 = 8'hc0 == io_state_in_3 ? 8'h5b : _GEN_1471; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1473 = 8'hc1 == io_state_in_3 ? 8'h58 : _GEN_1472; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1474 = 8'hc2 == io_state_in_3 ? 8'h5d : _GEN_1473; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1475 = 8'hc3 == io_state_in_3 ? 8'h5e : _GEN_1474; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1476 = 8'hc4 == io_state_in_3 ? 8'h57 : _GEN_1475; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1477 = 8'hc5 == io_state_in_3 ? 8'h54 : _GEN_1476; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1478 = 8'hc6 == io_state_in_3 ? 8'h51 : _GEN_1477; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1479 = 8'hc7 == io_state_in_3 ? 8'h52 : _GEN_1478; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1480 = 8'hc8 == io_state_in_3 ? 8'h43 : _GEN_1479; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1481 = 8'hc9 == io_state_in_3 ? 8'h40 : _GEN_1480; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1482 = 8'hca == io_state_in_3 ? 8'h45 : _GEN_1481; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1483 = 8'hcb == io_state_in_3 ? 8'h46 : _GEN_1482; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1484 = 8'hcc == io_state_in_3 ? 8'h4f : _GEN_1483; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1485 = 8'hcd == io_state_in_3 ? 8'h4c : _GEN_1484; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1486 = 8'hce == io_state_in_3 ? 8'h49 : _GEN_1485; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1487 = 8'hcf == io_state_in_3 ? 8'h4a : _GEN_1486; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1488 = 8'hd0 == io_state_in_3 ? 8'h6b : _GEN_1487; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1489 = 8'hd1 == io_state_in_3 ? 8'h68 : _GEN_1488; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1490 = 8'hd2 == io_state_in_3 ? 8'h6d : _GEN_1489; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1491 = 8'hd3 == io_state_in_3 ? 8'h6e : _GEN_1490; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1492 = 8'hd4 == io_state_in_3 ? 8'h67 : _GEN_1491; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1493 = 8'hd5 == io_state_in_3 ? 8'h64 : _GEN_1492; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1494 = 8'hd6 == io_state_in_3 ? 8'h61 : _GEN_1493; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1495 = 8'hd7 == io_state_in_3 ? 8'h62 : _GEN_1494; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1496 = 8'hd8 == io_state_in_3 ? 8'h73 : _GEN_1495; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1497 = 8'hd9 == io_state_in_3 ? 8'h70 : _GEN_1496; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1498 = 8'hda == io_state_in_3 ? 8'h75 : _GEN_1497; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1499 = 8'hdb == io_state_in_3 ? 8'h76 : _GEN_1498; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1500 = 8'hdc == io_state_in_3 ? 8'h7f : _GEN_1499; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1501 = 8'hdd == io_state_in_3 ? 8'h7c : _GEN_1500; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1502 = 8'hde == io_state_in_3 ? 8'h79 : _GEN_1501; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1503 = 8'hdf == io_state_in_3 ? 8'h7a : _GEN_1502; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1504 = 8'he0 == io_state_in_3 ? 8'h3b : _GEN_1503; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1505 = 8'he1 == io_state_in_3 ? 8'h38 : _GEN_1504; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1506 = 8'he2 == io_state_in_3 ? 8'h3d : _GEN_1505; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1507 = 8'he3 == io_state_in_3 ? 8'h3e : _GEN_1506; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1508 = 8'he4 == io_state_in_3 ? 8'h37 : _GEN_1507; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1509 = 8'he5 == io_state_in_3 ? 8'h34 : _GEN_1508; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1510 = 8'he6 == io_state_in_3 ? 8'h31 : _GEN_1509; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1511 = 8'he7 == io_state_in_3 ? 8'h32 : _GEN_1510; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1512 = 8'he8 == io_state_in_3 ? 8'h23 : _GEN_1511; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1513 = 8'he9 == io_state_in_3 ? 8'h20 : _GEN_1512; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1514 = 8'hea == io_state_in_3 ? 8'h25 : _GEN_1513; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1515 = 8'heb == io_state_in_3 ? 8'h26 : _GEN_1514; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1516 = 8'hec == io_state_in_3 ? 8'h2f : _GEN_1515; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1517 = 8'hed == io_state_in_3 ? 8'h2c : _GEN_1516; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1518 = 8'hee == io_state_in_3 ? 8'h29 : _GEN_1517; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1519 = 8'hef == io_state_in_3 ? 8'h2a : _GEN_1518; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1520 = 8'hf0 == io_state_in_3 ? 8'hb : _GEN_1519; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1521 = 8'hf1 == io_state_in_3 ? 8'h8 : _GEN_1520; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1522 = 8'hf2 == io_state_in_3 ? 8'hd : _GEN_1521; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1523 = 8'hf3 == io_state_in_3 ? 8'he : _GEN_1522; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1524 = 8'hf4 == io_state_in_3 ? 8'h7 : _GEN_1523; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1525 = 8'hf5 == io_state_in_3 ? 8'h4 : _GEN_1524; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1526 = 8'hf6 == io_state_in_3 ? 8'h1 : _GEN_1525; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1527 = 8'hf7 == io_state_in_3 ? 8'h2 : _GEN_1526; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1528 = 8'hf8 == io_state_in_3 ? 8'h13 : _GEN_1527; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1529 = 8'hf9 == io_state_in_3 ? 8'h10 : _GEN_1528; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1530 = 8'hfa == io_state_in_3 ? 8'h15 : _GEN_1529; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1531 = 8'hfb == io_state_in_3 ? 8'h16 : _GEN_1530; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1532 = 8'hfc == io_state_in_3 ? 8'h1f : _GEN_1531; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1533 = 8'hfd == io_state_in_3 ? 8'h1c : _GEN_1532; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1534 = 8'hfe == io_state_in_3 ? 8'h19 : _GEN_1533; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1535 = 8'hff == io_state_in_3 ? 8'h1a : _GEN_1534; // @[MixColumns.scala 127:{75,75}]
  wire [7:0] _GEN_1537 = 8'h1 == io_state_in_0 ? 8'h3 : 8'h0; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1538 = 8'h2 == io_state_in_0 ? 8'h6 : _GEN_1537; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1539 = 8'h3 == io_state_in_0 ? 8'h5 : _GEN_1538; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1540 = 8'h4 == io_state_in_0 ? 8'hc : _GEN_1539; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1541 = 8'h5 == io_state_in_0 ? 8'hf : _GEN_1540; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1542 = 8'h6 == io_state_in_0 ? 8'ha : _GEN_1541; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1543 = 8'h7 == io_state_in_0 ? 8'h9 : _GEN_1542; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1544 = 8'h8 == io_state_in_0 ? 8'h18 : _GEN_1543; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1545 = 8'h9 == io_state_in_0 ? 8'h1b : _GEN_1544; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1546 = 8'ha == io_state_in_0 ? 8'h1e : _GEN_1545; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1547 = 8'hb == io_state_in_0 ? 8'h1d : _GEN_1546; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1548 = 8'hc == io_state_in_0 ? 8'h14 : _GEN_1547; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1549 = 8'hd == io_state_in_0 ? 8'h17 : _GEN_1548; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1550 = 8'he == io_state_in_0 ? 8'h12 : _GEN_1549; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1551 = 8'hf == io_state_in_0 ? 8'h11 : _GEN_1550; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1552 = 8'h10 == io_state_in_0 ? 8'h30 : _GEN_1551; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1553 = 8'h11 == io_state_in_0 ? 8'h33 : _GEN_1552; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1554 = 8'h12 == io_state_in_0 ? 8'h36 : _GEN_1553; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1555 = 8'h13 == io_state_in_0 ? 8'h35 : _GEN_1554; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1556 = 8'h14 == io_state_in_0 ? 8'h3c : _GEN_1555; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1557 = 8'h15 == io_state_in_0 ? 8'h3f : _GEN_1556; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1558 = 8'h16 == io_state_in_0 ? 8'h3a : _GEN_1557; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1559 = 8'h17 == io_state_in_0 ? 8'h39 : _GEN_1558; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1560 = 8'h18 == io_state_in_0 ? 8'h28 : _GEN_1559; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1561 = 8'h19 == io_state_in_0 ? 8'h2b : _GEN_1560; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1562 = 8'h1a == io_state_in_0 ? 8'h2e : _GEN_1561; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1563 = 8'h1b == io_state_in_0 ? 8'h2d : _GEN_1562; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1564 = 8'h1c == io_state_in_0 ? 8'h24 : _GEN_1563; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1565 = 8'h1d == io_state_in_0 ? 8'h27 : _GEN_1564; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1566 = 8'h1e == io_state_in_0 ? 8'h22 : _GEN_1565; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1567 = 8'h1f == io_state_in_0 ? 8'h21 : _GEN_1566; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1568 = 8'h20 == io_state_in_0 ? 8'h60 : _GEN_1567; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1569 = 8'h21 == io_state_in_0 ? 8'h63 : _GEN_1568; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1570 = 8'h22 == io_state_in_0 ? 8'h66 : _GEN_1569; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1571 = 8'h23 == io_state_in_0 ? 8'h65 : _GEN_1570; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1572 = 8'h24 == io_state_in_0 ? 8'h6c : _GEN_1571; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1573 = 8'h25 == io_state_in_0 ? 8'h6f : _GEN_1572; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1574 = 8'h26 == io_state_in_0 ? 8'h6a : _GEN_1573; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1575 = 8'h27 == io_state_in_0 ? 8'h69 : _GEN_1574; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1576 = 8'h28 == io_state_in_0 ? 8'h78 : _GEN_1575; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1577 = 8'h29 == io_state_in_0 ? 8'h7b : _GEN_1576; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1578 = 8'h2a == io_state_in_0 ? 8'h7e : _GEN_1577; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1579 = 8'h2b == io_state_in_0 ? 8'h7d : _GEN_1578; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1580 = 8'h2c == io_state_in_0 ? 8'h74 : _GEN_1579; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1581 = 8'h2d == io_state_in_0 ? 8'h77 : _GEN_1580; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1582 = 8'h2e == io_state_in_0 ? 8'h72 : _GEN_1581; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1583 = 8'h2f == io_state_in_0 ? 8'h71 : _GEN_1582; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1584 = 8'h30 == io_state_in_0 ? 8'h50 : _GEN_1583; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1585 = 8'h31 == io_state_in_0 ? 8'h53 : _GEN_1584; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1586 = 8'h32 == io_state_in_0 ? 8'h56 : _GEN_1585; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1587 = 8'h33 == io_state_in_0 ? 8'h55 : _GEN_1586; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1588 = 8'h34 == io_state_in_0 ? 8'h5c : _GEN_1587; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1589 = 8'h35 == io_state_in_0 ? 8'h5f : _GEN_1588; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1590 = 8'h36 == io_state_in_0 ? 8'h5a : _GEN_1589; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1591 = 8'h37 == io_state_in_0 ? 8'h59 : _GEN_1590; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1592 = 8'h38 == io_state_in_0 ? 8'h48 : _GEN_1591; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1593 = 8'h39 == io_state_in_0 ? 8'h4b : _GEN_1592; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1594 = 8'h3a == io_state_in_0 ? 8'h4e : _GEN_1593; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1595 = 8'h3b == io_state_in_0 ? 8'h4d : _GEN_1594; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1596 = 8'h3c == io_state_in_0 ? 8'h44 : _GEN_1595; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1597 = 8'h3d == io_state_in_0 ? 8'h47 : _GEN_1596; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1598 = 8'h3e == io_state_in_0 ? 8'h42 : _GEN_1597; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1599 = 8'h3f == io_state_in_0 ? 8'h41 : _GEN_1598; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1600 = 8'h40 == io_state_in_0 ? 8'hc0 : _GEN_1599; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1601 = 8'h41 == io_state_in_0 ? 8'hc3 : _GEN_1600; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1602 = 8'h42 == io_state_in_0 ? 8'hc6 : _GEN_1601; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1603 = 8'h43 == io_state_in_0 ? 8'hc5 : _GEN_1602; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1604 = 8'h44 == io_state_in_0 ? 8'hcc : _GEN_1603; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1605 = 8'h45 == io_state_in_0 ? 8'hcf : _GEN_1604; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1606 = 8'h46 == io_state_in_0 ? 8'hca : _GEN_1605; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1607 = 8'h47 == io_state_in_0 ? 8'hc9 : _GEN_1606; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1608 = 8'h48 == io_state_in_0 ? 8'hd8 : _GEN_1607; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1609 = 8'h49 == io_state_in_0 ? 8'hdb : _GEN_1608; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1610 = 8'h4a == io_state_in_0 ? 8'hde : _GEN_1609; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1611 = 8'h4b == io_state_in_0 ? 8'hdd : _GEN_1610; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1612 = 8'h4c == io_state_in_0 ? 8'hd4 : _GEN_1611; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1613 = 8'h4d == io_state_in_0 ? 8'hd7 : _GEN_1612; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1614 = 8'h4e == io_state_in_0 ? 8'hd2 : _GEN_1613; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1615 = 8'h4f == io_state_in_0 ? 8'hd1 : _GEN_1614; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1616 = 8'h50 == io_state_in_0 ? 8'hf0 : _GEN_1615; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1617 = 8'h51 == io_state_in_0 ? 8'hf3 : _GEN_1616; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1618 = 8'h52 == io_state_in_0 ? 8'hf6 : _GEN_1617; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1619 = 8'h53 == io_state_in_0 ? 8'hf5 : _GEN_1618; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1620 = 8'h54 == io_state_in_0 ? 8'hfc : _GEN_1619; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1621 = 8'h55 == io_state_in_0 ? 8'hff : _GEN_1620; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1622 = 8'h56 == io_state_in_0 ? 8'hfa : _GEN_1621; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1623 = 8'h57 == io_state_in_0 ? 8'hf9 : _GEN_1622; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1624 = 8'h58 == io_state_in_0 ? 8'he8 : _GEN_1623; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1625 = 8'h59 == io_state_in_0 ? 8'heb : _GEN_1624; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1626 = 8'h5a == io_state_in_0 ? 8'hee : _GEN_1625; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1627 = 8'h5b == io_state_in_0 ? 8'hed : _GEN_1626; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1628 = 8'h5c == io_state_in_0 ? 8'he4 : _GEN_1627; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1629 = 8'h5d == io_state_in_0 ? 8'he7 : _GEN_1628; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1630 = 8'h5e == io_state_in_0 ? 8'he2 : _GEN_1629; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1631 = 8'h5f == io_state_in_0 ? 8'he1 : _GEN_1630; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1632 = 8'h60 == io_state_in_0 ? 8'ha0 : _GEN_1631; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1633 = 8'h61 == io_state_in_0 ? 8'ha3 : _GEN_1632; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1634 = 8'h62 == io_state_in_0 ? 8'ha6 : _GEN_1633; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1635 = 8'h63 == io_state_in_0 ? 8'ha5 : _GEN_1634; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1636 = 8'h64 == io_state_in_0 ? 8'hac : _GEN_1635; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1637 = 8'h65 == io_state_in_0 ? 8'haf : _GEN_1636; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1638 = 8'h66 == io_state_in_0 ? 8'haa : _GEN_1637; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1639 = 8'h67 == io_state_in_0 ? 8'ha9 : _GEN_1638; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1640 = 8'h68 == io_state_in_0 ? 8'hb8 : _GEN_1639; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1641 = 8'h69 == io_state_in_0 ? 8'hbb : _GEN_1640; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1642 = 8'h6a == io_state_in_0 ? 8'hbe : _GEN_1641; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1643 = 8'h6b == io_state_in_0 ? 8'hbd : _GEN_1642; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1644 = 8'h6c == io_state_in_0 ? 8'hb4 : _GEN_1643; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1645 = 8'h6d == io_state_in_0 ? 8'hb7 : _GEN_1644; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1646 = 8'h6e == io_state_in_0 ? 8'hb2 : _GEN_1645; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1647 = 8'h6f == io_state_in_0 ? 8'hb1 : _GEN_1646; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1648 = 8'h70 == io_state_in_0 ? 8'h90 : _GEN_1647; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1649 = 8'h71 == io_state_in_0 ? 8'h93 : _GEN_1648; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1650 = 8'h72 == io_state_in_0 ? 8'h96 : _GEN_1649; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1651 = 8'h73 == io_state_in_0 ? 8'h95 : _GEN_1650; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1652 = 8'h74 == io_state_in_0 ? 8'h9c : _GEN_1651; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1653 = 8'h75 == io_state_in_0 ? 8'h9f : _GEN_1652; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1654 = 8'h76 == io_state_in_0 ? 8'h9a : _GEN_1653; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1655 = 8'h77 == io_state_in_0 ? 8'h99 : _GEN_1654; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1656 = 8'h78 == io_state_in_0 ? 8'h88 : _GEN_1655; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1657 = 8'h79 == io_state_in_0 ? 8'h8b : _GEN_1656; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1658 = 8'h7a == io_state_in_0 ? 8'h8e : _GEN_1657; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1659 = 8'h7b == io_state_in_0 ? 8'h8d : _GEN_1658; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1660 = 8'h7c == io_state_in_0 ? 8'h84 : _GEN_1659; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1661 = 8'h7d == io_state_in_0 ? 8'h87 : _GEN_1660; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1662 = 8'h7e == io_state_in_0 ? 8'h82 : _GEN_1661; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1663 = 8'h7f == io_state_in_0 ? 8'h81 : _GEN_1662; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1664 = 8'h80 == io_state_in_0 ? 8'h9b : _GEN_1663; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1665 = 8'h81 == io_state_in_0 ? 8'h98 : _GEN_1664; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1666 = 8'h82 == io_state_in_0 ? 8'h9d : _GEN_1665; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1667 = 8'h83 == io_state_in_0 ? 8'h9e : _GEN_1666; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1668 = 8'h84 == io_state_in_0 ? 8'h97 : _GEN_1667; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1669 = 8'h85 == io_state_in_0 ? 8'h94 : _GEN_1668; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1670 = 8'h86 == io_state_in_0 ? 8'h91 : _GEN_1669; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1671 = 8'h87 == io_state_in_0 ? 8'h92 : _GEN_1670; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1672 = 8'h88 == io_state_in_0 ? 8'h83 : _GEN_1671; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1673 = 8'h89 == io_state_in_0 ? 8'h80 : _GEN_1672; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1674 = 8'h8a == io_state_in_0 ? 8'h85 : _GEN_1673; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1675 = 8'h8b == io_state_in_0 ? 8'h86 : _GEN_1674; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1676 = 8'h8c == io_state_in_0 ? 8'h8f : _GEN_1675; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1677 = 8'h8d == io_state_in_0 ? 8'h8c : _GEN_1676; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1678 = 8'h8e == io_state_in_0 ? 8'h89 : _GEN_1677; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1679 = 8'h8f == io_state_in_0 ? 8'h8a : _GEN_1678; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1680 = 8'h90 == io_state_in_0 ? 8'hab : _GEN_1679; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1681 = 8'h91 == io_state_in_0 ? 8'ha8 : _GEN_1680; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1682 = 8'h92 == io_state_in_0 ? 8'had : _GEN_1681; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1683 = 8'h93 == io_state_in_0 ? 8'hae : _GEN_1682; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1684 = 8'h94 == io_state_in_0 ? 8'ha7 : _GEN_1683; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1685 = 8'h95 == io_state_in_0 ? 8'ha4 : _GEN_1684; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1686 = 8'h96 == io_state_in_0 ? 8'ha1 : _GEN_1685; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1687 = 8'h97 == io_state_in_0 ? 8'ha2 : _GEN_1686; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1688 = 8'h98 == io_state_in_0 ? 8'hb3 : _GEN_1687; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1689 = 8'h99 == io_state_in_0 ? 8'hb0 : _GEN_1688; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1690 = 8'h9a == io_state_in_0 ? 8'hb5 : _GEN_1689; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1691 = 8'h9b == io_state_in_0 ? 8'hb6 : _GEN_1690; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1692 = 8'h9c == io_state_in_0 ? 8'hbf : _GEN_1691; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1693 = 8'h9d == io_state_in_0 ? 8'hbc : _GEN_1692; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1694 = 8'h9e == io_state_in_0 ? 8'hb9 : _GEN_1693; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1695 = 8'h9f == io_state_in_0 ? 8'hba : _GEN_1694; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1696 = 8'ha0 == io_state_in_0 ? 8'hfb : _GEN_1695; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1697 = 8'ha1 == io_state_in_0 ? 8'hf8 : _GEN_1696; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1698 = 8'ha2 == io_state_in_0 ? 8'hfd : _GEN_1697; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1699 = 8'ha3 == io_state_in_0 ? 8'hfe : _GEN_1698; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1700 = 8'ha4 == io_state_in_0 ? 8'hf7 : _GEN_1699; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1701 = 8'ha5 == io_state_in_0 ? 8'hf4 : _GEN_1700; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1702 = 8'ha6 == io_state_in_0 ? 8'hf1 : _GEN_1701; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1703 = 8'ha7 == io_state_in_0 ? 8'hf2 : _GEN_1702; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1704 = 8'ha8 == io_state_in_0 ? 8'he3 : _GEN_1703; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1705 = 8'ha9 == io_state_in_0 ? 8'he0 : _GEN_1704; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1706 = 8'haa == io_state_in_0 ? 8'he5 : _GEN_1705; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1707 = 8'hab == io_state_in_0 ? 8'he6 : _GEN_1706; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1708 = 8'hac == io_state_in_0 ? 8'hef : _GEN_1707; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1709 = 8'had == io_state_in_0 ? 8'hec : _GEN_1708; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1710 = 8'hae == io_state_in_0 ? 8'he9 : _GEN_1709; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1711 = 8'haf == io_state_in_0 ? 8'hea : _GEN_1710; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1712 = 8'hb0 == io_state_in_0 ? 8'hcb : _GEN_1711; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1713 = 8'hb1 == io_state_in_0 ? 8'hc8 : _GEN_1712; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1714 = 8'hb2 == io_state_in_0 ? 8'hcd : _GEN_1713; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1715 = 8'hb3 == io_state_in_0 ? 8'hce : _GEN_1714; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1716 = 8'hb4 == io_state_in_0 ? 8'hc7 : _GEN_1715; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1717 = 8'hb5 == io_state_in_0 ? 8'hc4 : _GEN_1716; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1718 = 8'hb6 == io_state_in_0 ? 8'hc1 : _GEN_1717; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1719 = 8'hb7 == io_state_in_0 ? 8'hc2 : _GEN_1718; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1720 = 8'hb8 == io_state_in_0 ? 8'hd3 : _GEN_1719; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1721 = 8'hb9 == io_state_in_0 ? 8'hd0 : _GEN_1720; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1722 = 8'hba == io_state_in_0 ? 8'hd5 : _GEN_1721; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1723 = 8'hbb == io_state_in_0 ? 8'hd6 : _GEN_1722; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1724 = 8'hbc == io_state_in_0 ? 8'hdf : _GEN_1723; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1725 = 8'hbd == io_state_in_0 ? 8'hdc : _GEN_1724; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1726 = 8'hbe == io_state_in_0 ? 8'hd9 : _GEN_1725; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1727 = 8'hbf == io_state_in_0 ? 8'hda : _GEN_1726; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1728 = 8'hc0 == io_state_in_0 ? 8'h5b : _GEN_1727; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1729 = 8'hc1 == io_state_in_0 ? 8'h58 : _GEN_1728; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1730 = 8'hc2 == io_state_in_0 ? 8'h5d : _GEN_1729; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1731 = 8'hc3 == io_state_in_0 ? 8'h5e : _GEN_1730; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1732 = 8'hc4 == io_state_in_0 ? 8'h57 : _GEN_1731; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1733 = 8'hc5 == io_state_in_0 ? 8'h54 : _GEN_1732; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1734 = 8'hc6 == io_state_in_0 ? 8'h51 : _GEN_1733; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1735 = 8'hc7 == io_state_in_0 ? 8'h52 : _GEN_1734; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1736 = 8'hc8 == io_state_in_0 ? 8'h43 : _GEN_1735; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1737 = 8'hc9 == io_state_in_0 ? 8'h40 : _GEN_1736; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1738 = 8'hca == io_state_in_0 ? 8'h45 : _GEN_1737; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1739 = 8'hcb == io_state_in_0 ? 8'h46 : _GEN_1738; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1740 = 8'hcc == io_state_in_0 ? 8'h4f : _GEN_1739; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1741 = 8'hcd == io_state_in_0 ? 8'h4c : _GEN_1740; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1742 = 8'hce == io_state_in_0 ? 8'h49 : _GEN_1741; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1743 = 8'hcf == io_state_in_0 ? 8'h4a : _GEN_1742; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1744 = 8'hd0 == io_state_in_0 ? 8'h6b : _GEN_1743; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1745 = 8'hd1 == io_state_in_0 ? 8'h68 : _GEN_1744; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1746 = 8'hd2 == io_state_in_0 ? 8'h6d : _GEN_1745; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1747 = 8'hd3 == io_state_in_0 ? 8'h6e : _GEN_1746; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1748 = 8'hd4 == io_state_in_0 ? 8'h67 : _GEN_1747; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1749 = 8'hd5 == io_state_in_0 ? 8'h64 : _GEN_1748; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1750 = 8'hd6 == io_state_in_0 ? 8'h61 : _GEN_1749; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1751 = 8'hd7 == io_state_in_0 ? 8'h62 : _GEN_1750; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1752 = 8'hd8 == io_state_in_0 ? 8'h73 : _GEN_1751; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1753 = 8'hd9 == io_state_in_0 ? 8'h70 : _GEN_1752; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1754 = 8'hda == io_state_in_0 ? 8'h75 : _GEN_1753; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1755 = 8'hdb == io_state_in_0 ? 8'h76 : _GEN_1754; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1756 = 8'hdc == io_state_in_0 ? 8'h7f : _GEN_1755; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1757 = 8'hdd == io_state_in_0 ? 8'h7c : _GEN_1756; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1758 = 8'hde == io_state_in_0 ? 8'h79 : _GEN_1757; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1759 = 8'hdf == io_state_in_0 ? 8'h7a : _GEN_1758; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1760 = 8'he0 == io_state_in_0 ? 8'h3b : _GEN_1759; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1761 = 8'he1 == io_state_in_0 ? 8'h38 : _GEN_1760; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1762 = 8'he2 == io_state_in_0 ? 8'h3d : _GEN_1761; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1763 = 8'he3 == io_state_in_0 ? 8'h3e : _GEN_1762; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1764 = 8'he4 == io_state_in_0 ? 8'h37 : _GEN_1763; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1765 = 8'he5 == io_state_in_0 ? 8'h34 : _GEN_1764; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1766 = 8'he6 == io_state_in_0 ? 8'h31 : _GEN_1765; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1767 = 8'he7 == io_state_in_0 ? 8'h32 : _GEN_1766; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1768 = 8'he8 == io_state_in_0 ? 8'h23 : _GEN_1767; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1769 = 8'he9 == io_state_in_0 ? 8'h20 : _GEN_1768; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1770 = 8'hea == io_state_in_0 ? 8'h25 : _GEN_1769; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1771 = 8'heb == io_state_in_0 ? 8'h26 : _GEN_1770; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1772 = 8'hec == io_state_in_0 ? 8'h2f : _GEN_1771; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1773 = 8'hed == io_state_in_0 ? 8'h2c : _GEN_1772; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1774 = 8'hee == io_state_in_0 ? 8'h29 : _GEN_1773; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1775 = 8'hef == io_state_in_0 ? 8'h2a : _GEN_1774; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1776 = 8'hf0 == io_state_in_0 ? 8'hb : _GEN_1775; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1777 = 8'hf1 == io_state_in_0 ? 8'h8 : _GEN_1776; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1778 = 8'hf2 == io_state_in_0 ? 8'hd : _GEN_1777; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1779 = 8'hf3 == io_state_in_0 ? 8'he : _GEN_1778; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1780 = 8'hf4 == io_state_in_0 ? 8'h7 : _GEN_1779; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1781 = 8'hf5 == io_state_in_0 ? 8'h4 : _GEN_1780; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1782 = 8'hf6 == io_state_in_0 ? 8'h1 : _GEN_1781; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1783 = 8'hf7 == io_state_in_0 ? 8'h2 : _GEN_1782; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1784 = 8'hf8 == io_state_in_0 ? 8'h13 : _GEN_1783; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1785 = 8'hf9 == io_state_in_0 ? 8'h10 : _GEN_1784; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1786 = 8'hfa == io_state_in_0 ? 8'h15 : _GEN_1785; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1787 = 8'hfb == io_state_in_0 ? 8'h16 : _GEN_1786; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1788 = 8'hfc == io_state_in_0 ? 8'h1f : _GEN_1787; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1789 = 8'hfd == io_state_in_0 ? 8'h1c : _GEN_1788; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1790 = 8'hfe == io_state_in_0 ? 8'h19 : _GEN_1789; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _GEN_1791 = 8'hff == io_state_in_0 ? 8'h1a : _GEN_1790; // @[MixColumns.scala 128:{41,41}]
  wire [7:0] _tmp_state_3_T = _GEN_1791 ^ io_state_in_1; // @[MixColumns.scala 128:41]
  wire [7:0] _tmp_state_3_T_1 = _tmp_state_3_T ^ io_state_in_2; // @[MixColumns.scala 128:58]
  wire [7:0] _GEN_1793 = 8'h1 == io_state_in_3 ? 8'h2 : 8'h0; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1794 = 8'h2 == io_state_in_3 ? 8'h4 : _GEN_1793; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1795 = 8'h3 == io_state_in_3 ? 8'h6 : _GEN_1794; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1796 = 8'h4 == io_state_in_3 ? 8'h8 : _GEN_1795; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1797 = 8'h5 == io_state_in_3 ? 8'ha : _GEN_1796; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1798 = 8'h6 == io_state_in_3 ? 8'hc : _GEN_1797; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1799 = 8'h7 == io_state_in_3 ? 8'he : _GEN_1798; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1800 = 8'h8 == io_state_in_3 ? 8'h10 : _GEN_1799; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1801 = 8'h9 == io_state_in_3 ? 8'h12 : _GEN_1800; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1802 = 8'ha == io_state_in_3 ? 8'h14 : _GEN_1801; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1803 = 8'hb == io_state_in_3 ? 8'h16 : _GEN_1802; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1804 = 8'hc == io_state_in_3 ? 8'h18 : _GEN_1803; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1805 = 8'hd == io_state_in_3 ? 8'h1a : _GEN_1804; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1806 = 8'he == io_state_in_3 ? 8'h1c : _GEN_1805; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1807 = 8'hf == io_state_in_3 ? 8'h1e : _GEN_1806; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1808 = 8'h10 == io_state_in_3 ? 8'h20 : _GEN_1807; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1809 = 8'h11 == io_state_in_3 ? 8'h22 : _GEN_1808; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1810 = 8'h12 == io_state_in_3 ? 8'h24 : _GEN_1809; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1811 = 8'h13 == io_state_in_3 ? 8'h26 : _GEN_1810; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1812 = 8'h14 == io_state_in_3 ? 8'h28 : _GEN_1811; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1813 = 8'h15 == io_state_in_3 ? 8'h2a : _GEN_1812; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1814 = 8'h16 == io_state_in_3 ? 8'h2c : _GEN_1813; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1815 = 8'h17 == io_state_in_3 ? 8'h2e : _GEN_1814; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1816 = 8'h18 == io_state_in_3 ? 8'h30 : _GEN_1815; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1817 = 8'h19 == io_state_in_3 ? 8'h32 : _GEN_1816; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1818 = 8'h1a == io_state_in_3 ? 8'h34 : _GEN_1817; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1819 = 8'h1b == io_state_in_3 ? 8'h36 : _GEN_1818; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1820 = 8'h1c == io_state_in_3 ? 8'h38 : _GEN_1819; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1821 = 8'h1d == io_state_in_3 ? 8'h3a : _GEN_1820; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1822 = 8'h1e == io_state_in_3 ? 8'h3c : _GEN_1821; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1823 = 8'h1f == io_state_in_3 ? 8'h3e : _GEN_1822; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1824 = 8'h20 == io_state_in_3 ? 8'h40 : _GEN_1823; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1825 = 8'h21 == io_state_in_3 ? 8'h42 : _GEN_1824; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1826 = 8'h22 == io_state_in_3 ? 8'h44 : _GEN_1825; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1827 = 8'h23 == io_state_in_3 ? 8'h46 : _GEN_1826; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1828 = 8'h24 == io_state_in_3 ? 8'h48 : _GEN_1827; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1829 = 8'h25 == io_state_in_3 ? 8'h4a : _GEN_1828; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1830 = 8'h26 == io_state_in_3 ? 8'h4c : _GEN_1829; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1831 = 8'h27 == io_state_in_3 ? 8'h4e : _GEN_1830; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1832 = 8'h28 == io_state_in_3 ? 8'h50 : _GEN_1831; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1833 = 8'h29 == io_state_in_3 ? 8'h52 : _GEN_1832; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1834 = 8'h2a == io_state_in_3 ? 8'h54 : _GEN_1833; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1835 = 8'h2b == io_state_in_3 ? 8'h56 : _GEN_1834; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1836 = 8'h2c == io_state_in_3 ? 8'h58 : _GEN_1835; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1837 = 8'h2d == io_state_in_3 ? 8'h5a : _GEN_1836; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1838 = 8'h2e == io_state_in_3 ? 8'h5c : _GEN_1837; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1839 = 8'h2f == io_state_in_3 ? 8'h5e : _GEN_1838; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1840 = 8'h30 == io_state_in_3 ? 8'h60 : _GEN_1839; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1841 = 8'h31 == io_state_in_3 ? 8'h62 : _GEN_1840; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1842 = 8'h32 == io_state_in_3 ? 8'h64 : _GEN_1841; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1843 = 8'h33 == io_state_in_3 ? 8'h66 : _GEN_1842; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1844 = 8'h34 == io_state_in_3 ? 8'h68 : _GEN_1843; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1845 = 8'h35 == io_state_in_3 ? 8'h6a : _GEN_1844; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1846 = 8'h36 == io_state_in_3 ? 8'h6c : _GEN_1845; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1847 = 8'h37 == io_state_in_3 ? 8'h6e : _GEN_1846; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1848 = 8'h38 == io_state_in_3 ? 8'h70 : _GEN_1847; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1849 = 8'h39 == io_state_in_3 ? 8'h72 : _GEN_1848; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1850 = 8'h3a == io_state_in_3 ? 8'h74 : _GEN_1849; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1851 = 8'h3b == io_state_in_3 ? 8'h76 : _GEN_1850; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1852 = 8'h3c == io_state_in_3 ? 8'h78 : _GEN_1851; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1853 = 8'h3d == io_state_in_3 ? 8'h7a : _GEN_1852; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1854 = 8'h3e == io_state_in_3 ? 8'h7c : _GEN_1853; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1855 = 8'h3f == io_state_in_3 ? 8'h7e : _GEN_1854; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1856 = 8'h40 == io_state_in_3 ? 8'h80 : _GEN_1855; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1857 = 8'h41 == io_state_in_3 ? 8'h82 : _GEN_1856; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1858 = 8'h42 == io_state_in_3 ? 8'h84 : _GEN_1857; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1859 = 8'h43 == io_state_in_3 ? 8'h86 : _GEN_1858; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1860 = 8'h44 == io_state_in_3 ? 8'h88 : _GEN_1859; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1861 = 8'h45 == io_state_in_3 ? 8'h8a : _GEN_1860; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1862 = 8'h46 == io_state_in_3 ? 8'h8c : _GEN_1861; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1863 = 8'h47 == io_state_in_3 ? 8'h8e : _GEN_1862; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1864 = 8'h48 == io_state_in_3 ? 8'h90 : _GEN_1863; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1865 = 8'h49 == io_state_in_3 ? 8'h92 : _GEN_1864; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1866 = 8'h4a == io_state_in_3 ? 8'h94 : _GEN_1865; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1867 = 8'h4b == io_state_in_3 ? 8'h96 : _GEN_1866; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1868 = 8'h4c == io_state_in_3 ? 8'h98 : _GEN_1867; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1869 = 8'h4d == io_state_in_3 ? 8'h9a : _GEN_1868; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1870 = 8'h4e == io_state_in_3 ? 8'h9c : _GEN_1869; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1871 = 8'h4f == io_state_in_3 ? 8'h9e : _GEN_1870; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1872 = 8'h50 == io_state_in_3 ? 8'ha0 : _GEN_1871; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1873 = 8'h51 == io_state_in_3 ? 8'ha2 : _GEN_1872; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1874 = 8'h52 == io_state_in_3 ? 8'ha4 : _GEN_1873; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1875 = 8'h53 == io_state_in_3 ? 8'ha6 : _GEN_1874; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1876 = 8'h54 == io_state_in_3 ? 8'ha8 : _GEN_1875; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1877 = 8'h55 == io_state_in_3 ? 8'haa : _GEN_1876; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1878 = 8'h56 == io_state_in_3 ? 8'hac : _GEN_1877; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1879 = 8'h57 == io_state_in_3 ? 8'hae : _GEN_1878; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1880 = 8'h58 == io_state_in_3 ? 8'hb0 : _GEN_1879; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1881 = 8'h59 == io_state_in_3 ? 8'hb2 : _GEN_1880; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1882 = 8'h5a == io_state_in_3 ? 8'hb4 : _GEN_1881; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1883 = 8'h5b == io_state_in_3 ? 8'hb6 : _GEN_1882; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1884 = 8'h5c == io_state_in_3 ? 8'hb8 : _GEN_1883; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1885 = 8'h5d == io_state_in_3 ? 8'hba : _GEN_1884; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1886 = 8'h5e == io_state_in_3 ? 8'hbc : _GEN_1885; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1887 = 8'h5f == io_state_in_3 ? 8'hbe : _GEN_1886; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1888 = 8'h60 == io_state_in_3 ? 8'hc0 : _GEN_1887; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1889 = 8'h61 == io_state_in_3 ? 8'hc2 : _GEN_1888; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1890 = 8'h62 == io_state_in_3 ? 8'hc4 : _GEN_1889; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1891 = 8'h63 == io_state_in_3 ? 8'hc6 : _GEN_1890; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1892 = 8'h64 == io_state_in_3 ? 8'hc8 : _GEN_1891; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1893 = 8'h65 == io_state_in_3 ? 8'hca : _GEN_1892; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1894 = 8'h66 == io_state_in_3 ? 8'hcc : _GEN_1893; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1895 = 8'h67 == io_state_in_3 ? 8'hce : _GEN_1894; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1896 = 8'h68 == io_state_in_3 ? 8'hd0 : _GEN_1895; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1897 = 8'h69 == io_state_in_3 ? 8'hd2 : _GEN_1896; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1898 = 8'h6a == io_state_in_3 ? 8'hd4 : _GEN_1897; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1899 = 8'h6b == io_state_in_3 ? 8'hd6 : _GEN_1898; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1900 = 8'h6c == io_state_in_3 ? 8'hd8 : _GEN_1899; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1901 = 8'h6d == io_state_in_3 ? 8'hda : _GEN_1900; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1902 = 8'h6e == io_state_in_3 ? 8'hdc : _GEN_1901; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1903 = 8'h6f == io_state_in_3 ? 8'hde : _GEN_1902; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1904 = 8'h70 == io_state_in_3 ? 8'he0 : _GEN_1903; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1905 = 8'h71 == io_state_in_3 ? 8'he2 : _GEN_1904; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1906 = 8'h72 == io_state_in_3 ? 8'he4 : _GEN_1905; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1907 = 8'h73 == io_state_in_3 ? 8'he6 : _GEN_1906; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1908 = 8'h74 == io_state_in_3 ? 8'he8 : _GEN_1907; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1909 = 8'h75 == io_state_in_3 ? 8'hea : _GEN_1908; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1910 = 8'h76 == io_state_in_3 ? 8'hec : _GEN_1909; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1911 = 8'h77 == io_state_in_3 ? 8'hee : _GEN_1910; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1912 = 8'h78 == io_state_in_3 ? 8'hf0 : _GEN_1911; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1913 = 8'h79 == io_state_in_3 ? 8'hf2 : _GEN_1912; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1914 = 8'h7a == io_state_in_3 ? 8'hf4 : _GEN_1913; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1915 = 8'h7b == io_state_in_3 ? 8'hf6 : _GEN_1914; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1916 = 8'h7c == io_state_in_3 ? 8'hf8 : _GEN_1915; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1917 = 8'h7d == io_state_in_3 ? 8'hfa : _GEN_1916; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1918 = 8'h7e == io_state_in_3 ? 8'hfc : _GEN_1917; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1919 = 8'h7f == io_state_in_3 ? 8'hfe : _GEN_1918; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1920 = 8'h80 == io_state_in_3 ? 8'h1b : _GEN_1919; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1921 = 8'h81 == io_state_in_3 ? 8'h19 : _GEN_1920; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1922 = 8'h82 == io_state_in_3 ? 8'h1f : _GEN_1921; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1923 = 8'h83 == io_state_in_3 ? 8'h1d : _GEN_1922; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1924 = 8'h84 == io_state_in_3 ? 8'h13 : _GEN_1923; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1925 = 8'h85 == io_state_in_3 ? 8'h11 : _GEN_1924; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1926 = 8'h86 == io_state_in_3 ? 8'h17 : _GEN_1925; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1927 = 8'h87 == io_state_in_3 ? 8'h15 : _GEN_1926; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1928 = 8'h88 == io_state_in_3 ? 8'hb : _GEN_1927; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1929 = 8'h89 == io_state_in_3 ? 8'h9 : _GEN_1928; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1930 = 8'h8a == io_state_in_3 ? 8'hf : _GEN_1929; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1931 = 8'h8b == io_state_in_3 ? 8'hd : _GEN_1930; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1932 = 8'h8c == io_state_in_3 ? 8'h3 : _GEN_1931; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1933 = 8'h8d == io_state_in_3 ? 8'h1 : _GEN_1932; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1934 = 8'h8e == io_state_in_3 ? 8'h7 : _GEN_1933; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1935 = 8'h8f == io_state_in_3 ? 8'h5 : _GEN_1934; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1936 = 8'h90 == io_state_in_3 ? 8'h3b : _GEN_1935; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1937 = 8'h91 == io_state_in_3 ? 8'h39 : _GEN_1936; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1938 = 8'h92 == io_state_in_3 ? 8'h3f : _GEN_1937; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1939 = 8'h93 == io_state_in_3 ? 8'h3d : _GEN_1938; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1940 = 8'h94 == io_state_in_3 ? 8'h33 : _GEN_1939; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1941 = 8'h95 == io_state_in_3 ? 8'h31 : _GEN_1940; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1942 = 8'h96 == io_state_in_3 ? 8'h37 : _GEN_1941; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1943 = 8'h97 == io_state_in_3 ? 8'h35 : _GEN_1942; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1944 = 8'h98 == io_state_in_3 ? 8'h2b : _GEN_1943; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1945 = 8'h99 == io_state_in_3 ? 8'h29 : _GEN_1944; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1946 = 8'h9a == io_state_in_3 ? 8'h2f : _GEN_1945; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1947 = 8'h9b == io_state_in_3 ? 8'h2d : _GEN_1946; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1948 = 8'h9c == io_state_in_3 ? 8'h23 : _GEN_1947; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1949 = 8'h9d == io_state_in_3 ? 8'h21 : _GEN_1948; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1950 = 8'h9e == io_state_in_3 ? 8'h27 : _GEN_1949; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1951 = 8'h9f == io_state_in_3 ? 8'h25 : _GEN_1950; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1952 = 8'ha0 == io_state_in_3 ? 8'h5b : _GEN_1951; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1953 = 8'ha1 == io_state_in_3 ? 8'h59 : _GEN_1952; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1954 = 8'ha2 == io_state_in_3 ? 8'h5f : _GEN_1953; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1955 = 8'ha3 == io_state_in_3 ? 8'h5d : _GEN_1954; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1956 = 8'ha4 == io_state_in_3 ? 8'h53 : _GEN_1955; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1957 = 8'ha5 == io_state_in_3 ? 8'h51 : _GEN_1956; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1958 = 8'ha6 == io_state_in_3 ? 8'h57 : _GEN_1957; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1959 = 8'ha7 == io_state_in_3 ? 8'h55 : _GEN_1958; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1960 = 8'ha8 == io_state_in_3 ? 8'h4b : _GEN_1959; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1961 = 8'ha9 == io_state_in_3 ? 8'h49 : _GEN_1960; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1962 = 8'haa == io_state_in_3 ? 8'h4f : _GEN_1961; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1963 = 8'hab == io_state_in_3 ? 8'h4d : _GEN_1962; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1964 = 8'hac == io_state_in_3 ? 8'h43 : _GEN_1963; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1965 = 8'had == io_state_in_3 ? 8'h41 : _GEN_1964; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1966 = 8'hae == io_state_in_3 ? 8'h47 : _GEN_1965; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1967 = 8'haf == io_state_in_3 ? 8'h45 : _GEN_1966; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1968 = 8'hb0 == io_state_in_3 ? 8'h7b : _GEN_1967; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1969 = 8'hb1 == io_state_in_3 ? 8'h79 : _GEN_1968; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1970 = 8'hb2 == io_state_in_3 ? 8'h7f : _GEN_1969; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1971 = 8'hb3 == io_state_in_3 ? 8'h7d : _GEN_1970; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1972 = 8'hb4 == io_state_in_3 ? 8'h73 : _GEN_1971; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1973 = 8'hb5 == io_state_in_3 ? 8'h71 : _GEN_1972; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1974 = 8'hb6 == io_state_in_3 ? 8'h77 : _GEN_1973; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1975 = 8'hb7 == io_state_in_3 ? 8'h75 : _GEN_1974; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1976 = 8'hb8 == io_state_in_3 ? 8'h6b : _GEN_1975; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1977 = 8'hb9 == io_state_in_3 ? 8'h69 : _GEN_1976; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1978 = 8'hba == io_state_in_3 ? 8'h6f : _GEN_1977; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1979 = 8'hbb == io_state_in_3 ? 8'h6d : _GEN_1978; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1980 = 8'hbc == io_state_in_3 ? 8'h63 : _GEN_1979; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1981 = 8'hbd == io_state_in_3 ? 8'h61 : _GEN_1980; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1982 = 8'hbe == io_state_in_3 ? 8'h67 : _GEN_1981; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1983 = 8'hbf == io_state_in_3 ? 8'h65 : _GEN_1982; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1984 = 8'hc0 == io_state_in_3 ? 8'h9b : _GEN_1983; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1985 = 8'hc1 == io_state_in_3 ? 8'h99 : _GEN_1984; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1986 = 8'hc2 == io_state_in_3 ? 8'h9f : _GEN_1985; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1987 = 8'hc3 == io_state_in_3 ? 8'h9d : _GEN_1986; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1988 = 8'hc4 == io_state_in_3 ? 8'h93 : _GEN_1987; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1989 = 8'hc5 == io_state_in_3 ? 8'h91 : _GEN_1988; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1990 = 8'hc6 == io_state_in_3 ? 8'h97 : _GEN_1989; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1991 = 8'hc7 == io_state_in_3 ? 8'h95 : _GEN_1990; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1992 = 8'hc8 == io_state_in_3 ? 8'h8b : _GEN_1991; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1993 = 8'hc9 == io_state_in_3 ? 8'h89 : _GEN_1992; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1994 = 8'hca == io_state_in_3 ? 8'h8f : _GEN_1993; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1995 = 8'hcb == io_state_in_3 ? 8'h8d : _GEN_1994; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1996 = 8'hcc == io_state_in_3 ? 8'h83 : _GEN_1995; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1997 = 8'hcd == io_state_in_3 ? 8'h81 : _GEN_1996; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1998 = 8'hce == io_state_in_3 ? 8'h87 : _GEN_1997; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_1999 = 8'hcf == io_state_in_3 ? 8'h85 : _GEN_1998; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2000 = 8'hd0 == io_state_in_3 ? 8'hbb : _GEN_1999; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2001 = 8'hd1 == io_state_in_3 ? 8'hb9 : _GEN_2000; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2002 = 8'hd2 == io_state_in_3 ? 8'hbf : _GEN_2001; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2003 = 8'hd3 == io_state_in_3 ? 8'hbd : _GEN_2002; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2004 = 8'hd4 == io_state_in_3 ? 8'hb3 : _GEN_2003; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2005 = 8'hd5 == io_state_in_3 ? 8'hb1 : _GEN_2004; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2006 = 8'hd6 == io_state_in_3 ? 8'hb7 : _GEN_2005; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2007 = 8'hd7 == io_state_in_3 ? 8'hb5 : _GEN_2006; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2008 = 8'hd8 == io_state_in_3 ? 8'hab : _GEN_2007; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2009 = 8'hd9 == io_state_in_3 ? 8'ha9 : _GEN_2008; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2010 = 8'hda == io_state_in_3 ? 8'haf : _GEN_2009; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2011 = 8'hdb == io_state_in_3 ? 8'had : _GEN_2010; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2012 = 8'hdc == io_state_in_3 ? 8'ha3 : _GEN_2011; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2013 = 8'hdd == io_state_in_3 ? 8'ha1 : _GEN_2012; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2014 = 8'hde == io_state_in_3 ? 8'ha7 : _GEN_2013; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2015 = 8'hdf == io_state_in_3 ? 8'ha5 : _GEN_2014; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2016 = 8'he0 == io_state_in_3 ? 8'hdb : _GEN_2015; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2017 = 8'he1 == io_state_in_3 ? 8'hd9 : _GEN_2016; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2018 = 8'he2 == io_state_in_3 ? 8'hdf : _GEN_2017; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2019 = 8'he3 == io_state_in_3 ? 8'hdd : _GEN_2018; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2020 = 8'he4 == io_state_in_3 ? 8'hd3 : _GEN_2019; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2021 = 8'he5 == io_state_in_3 ? 8'hd1 : _GEN_2020; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2022 = 8'he6 == io_state_in_3 ? 8'hd7 : _GEN_2021; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2023 = 8'he7 == io_state_in_3 ? 8'hd5 : _GEN_2022; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2024 = 8'he8 == io_state_in_3 ? 8'hcb : _GEN_2023; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2025 = 8'he9 == io_state_in_3 ? 8'hc9 : _GEN_2024; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2026 = 8'hea == io_state_in_3 ? 8'hcf : _GEN_2025; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2027 = 8'heb == io_state_in_3 ? 8'hcd : _GEN_2026; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2028 = 8'hec == io_state_in_3 ? 8'hc3 : _GEN_2027; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2029 = 8'hed == io_state_in_3 ? 8'hc1 : _GEN_2028; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2030 = 8'hee == io_state_in_3 ? 8'hc7 : _GEN_2029; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2031 = 8'hef == io_state_in_3 ? 8'hc5 : _GEN_2030; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2032 = 8'hf0 == io_state_in_3 ? 8'hfb : _GEN_2031; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2033 = 8'hf1 == io_state_in_3 ? 8'hf9 : _GEN_2032; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2034 = 8'hf2 == io_state_in_3 ? 8'hff : _GEN_2033; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2035 = 8'hf3 == io_state_in_3 ? 8'hfd : _GEN_2034; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2036 = 8'hf4 == io_state_in_3 ? 8'hf3 : _GEN_2035; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2037 = 8'hf5 == io_state_in_3 ? 8'hf1 : _GEN_2036; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2038 = 8'hf6 == io_state_in_3 ? 8'hf7 : _GEN_2037; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2039 = 8'hf7 == io_state_in_3 ? 8'hf5 : _GEN_2038; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2040 = 8'hf8 == io_state_in_3 ? 8'heb : _GEN_2039; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2041 = 8'hf9 == io_state_in_3 ? 8'he9 : _GEN_2040; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2042 = 8'hfa == io_state_in_3 ? 8'hef : _GEN_2041; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2043 = 8'hfb == io_state_in_3 ? 8'hed : _GEN_2042; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2044 = 8'hfc == io_state_in_3 ? 8'he3 : _GEN_2043; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2045 = 8'hfd == io_state_in_3 ? 8'he1 : _GEN_2044; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2046 = 8'hfe == io_state_in_3 ? 8'he7 : _GEN_2045; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2047 = 8'hff == io_state_in_3 ? 8'he5 : _GEN_2046; // @[MixColumns.scala 128:{75,75}]
  wire [7:0] _GEN_2049 = 8'h1 == io_state_in_4 ? 8'h2 : 8'h0; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2050 = 8'h2 == io_state_in_4 ? 8'h4 : _GEN_2049; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2051 = 8'h3 == io_state_in_4 ? 8'h6 : _GEN_2050; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2052 = 8'h4 == io_state_in_4 ? 8'h8 : _GEN_2051; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2053 = 8'h5 == io_state_in_4 ? 8'ha : _GEN_2052; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2054 = 8'h6 == io_state_in_4 ? 8'hc : _GEN_2053; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2055 = 8'h7 == io_state_in_4 ? 8'he : _GEN_2054; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2056 = 8'h8 == io_state_in_4 ? 8'h10 : _GEN_2055; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2057 = 8'h9 == io_state_in_4 ? 8'h12 : _GEN_2056; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2058 = 8'ha == io_state_in_4 ? 8'h14 : _GEN_2057; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2059 = 8'hb == io_state_in_4 ? 8'h16 : _GEN_2058; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2060 = 8'hc == io_state_in_4 ? 8'h18 : _GEN_2059; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2061 = 8'hd == io_state_in_4 ? 8'h1a : _GEN_2060; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2062 = 8'he == io_state_in_4 ? 8'h1c : _GEN_2061; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2063 = 8'hf == io_state_in_4 ? 8'h1e : _GEN_2062; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2064 = 8'h10 == io_state_in_4 ? 8'h20 : _GEN_2063; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2065 = 8'h11 == io_state_in_4 ? 8'h22 : _GEN_2064; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2066 = 8'h12 == io_state_in_4 ? 8'h24 : _GEN_2065; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2067 = 8'h13 == io_state_in_4 ? 8'h26 : _GEN_2066; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2068 = 8'h14 == io_state_in_4 ? 8'h28 : _GEN_2067; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2069 = 8'h15 == io_state_in_4 ? 8'h2a : _GEN_2068; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2070 = 8'h16 == io_state_in_4 ? 8'h2c : _GEN_2069; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2071 = 8'h17 == io_state_in_4 ? 8'h2e : _GEN_2070; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2072 = 8'h18 == io_state_in_4 ? 8'h30 : _GEN_2071; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2073 = 8'h19 == io_state_in_4 ? 8'h32 : _GEN_2072; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2074 = 8'h1a == io_state_in_4 ? 8'h34 : _GEN_2073; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2075 = 8'h1b == io_state_in_4 ? 8'h36 : _GEN_2074; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2076 = 8'h1c == io_state_in_4 ? 8'h38 : _GEN_2075; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2077 = 8'h1d == io_state_in_4 ? 8'h3a : _GEN_2076; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2078 = 8'h1e == io_state_in_4 ? 8'h3c : _GEN_2077; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2079 = 8'h1f == io_state_in_4 ? 8'h3e : _GEN_2078; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2080 = 8'h20 == io_state_in_4 ? 8'h40 : _GEN_2079; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2081 = 8'h21 == io_state_in_4 ? 8'h42 : _GEN_2080; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2082 = 8'h22 == io_state_in_4 ? 8'h44 : _GEN_2081; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2083 = 8'h23 == io_state_in_4 ? 8'h46 : _GEN_2082; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2084 = 8'h24 == io_state_in_4 ? 8'h48 : _GEN_2083; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2085 = 8'h25 == io_state_in_4 ? 8'h4a : _GEN_2084; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2086 = 8'h26 == io_state_in_4 ? 8'h4c : _GEN_2085; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2087 = 8'h27 == io_state_in_4 ? 8'h4e : _GEN_2086; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2088 = 8'h28 == io_state_in_4 ? 8'h50 : _GEN_2087; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2089 = 8'h29 == io_state_in_4 ? 8'h52 : _GEN_2088; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2090 = 8'h2a == io_state_in_4 ? 8'h54 : _GEN_2089; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2091 = 8'h2b == io_state_in_4 ? 8'h56 : _GEN_2090; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2092 = 8'h2c == io_state_in_4 ? 8'h58 : _GEN_2091; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2093 = 8'h2d == io_state_in_4 ? 8'h5a : _GEN_2092; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2094 = 8'h2e == io_state_in_4 ? 8'h5c : _GEN_2093; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2095 = 8'h2f == io_state_in_4 ? 8'h5e : _GEN_2094; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2096 = 8'h30 == io_state_in_4 ? 8'h60 : _GEN_2095; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2097 = 8'h31 == io_state_in_4 ? 8'h62 : _GEN_2096; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2098 = 8'h32 == io_state_in_4 ? 8'h64 : _GEN_2097; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2099 = 8'h33 == io_state_in_4 ? 8'h66 : _GEN_2098; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2100 = 8'h34 == io_state_in_4 ? 8'h68 : _GEN_2099; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2101 = 8'h35 == io_state_in_4 ? 8'h6a : _GEN_2100; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2102 = 8'h36 == io_state_in_4 ? 8'h6c : _GEN_2101; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2103 = 8'h37 == io_state_in_4 ? 8'h6e : _GEN_2102; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2104 = 8'h38 == io_state_in_4 ? 8'h70 : _GEN_2103; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2105 = 8'h39 == io_state_in_4 ? 8'h72 : _GEN_2104; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2106 = 8'h3a == io_state_in_4 ? 8'h74 : _GEN_2105; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2107 = 8'h3b == io_state_in_4 ? 8'h76 : _GEN_2106; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2108 = 8'h3c == io_state_in_4 ? 8'h78 : _GEN_2107; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2109 = 8'h3d == io_state_in_4 ? 8'h7a : _GEN_2108; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2110 = 8'h3e == io_state_in_4 ? 8'h7c : _GEN_2109; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2111 = 8'h3f == io_state_in_4 ? 8'h7e : _GEN_2110; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2112 = 8'h40 == io_state_in_4 ? 8'h80 : _GEN_2111; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2113 = 8'h41 == io_state_in_4 ? 8'h82 : _GEN_2112; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2114 = 8'h42 == io_state_in_4 ? 8'h84 : _GEN_2113; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2115 = 8'h43 == io_state_in_4 ? 8'h86 : _GEN_2114; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2116 = 8'h44 == io_state_in_4 ? 8'h88 : _GEN_2115; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2117 = 8'h45 == io_state_in_4 ? 8'h8a : _GEN_2116; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2118 = 8'h46 == io_state_in_4 ? 8'h8c : _GEN_2117; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2119 = 8'h47 == io_state_in_4 ? 8'h8e : _GEN_2118; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2120 = 8'h48 == io_state_in_4 ? 8'h90 : _GEN_2119; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2121 = 8'h49 == io_state_in_4 ? 8'h92 : _GEN_2120; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2122 = 8'h4a == io_state_in_4 ? 8'h94 : _GEN_2121; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2123 = 8'h4b == io_state_in_4 ? 8'h96 : _GEN_2122; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2124 = 8'h4c == io_state_in_4 ? 8'h98 : _GEN_2123; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2125 = 8'h4d == io_state_in_4 ? 8'h9a : _GEN_2124; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2126 = 8'h4e == io_state_in_4 ? 8'h9c : _GEN_2125; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2127 = 8'h4f == io_state_in_4 ? 8'h9e : _GEN_2126; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2128 = 8'h50 == io_state_in_4 ? 8'ha0 : _GEN_2127; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2129 = 8'h51 == io_state_in_4 ? 8'ha2 : _GEN_2128; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2130 = 8'h52 == io_state_in_4 ? 8'ha4 : _GEN_2129; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2131 = 8'h53 == io_state_in_4 ? 8'ha6 : _GEN_2130; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2132 = 8'h54 == io_state_in_4 ? 8'ha8 : _GEN_2131; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2133 = 8'h55 == io_state_in_4 ? 8'haa : _GEN_2132; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2134 = 8'h56 == io_state_in_4 ? 8'hac : _GEN_2133; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2135 = 8'h57 == io_state_in_4 ? 8'hae : _GEN_2134; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2136 = 8'h58 == io_state_in_4 ? 8'hb0 : _GEN_2135; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2137 = 8'h59 == io_state_in_4 ? 8'hb2 : _GEN_2136; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2138 = 8'h5a == io_state_in_4 ? 8'hb4 : _GEN_2137; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2139 = 8'h5b == io_state_in_4 ? 8'hb6 : _GEN_2138; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2140 = 8'h5c == io_state_in_4 ? 8'hb8 : _GEN_2139; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2141 = 8'h5d == io_state_in_4 ? 8'hba : _GEN_2140; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2142 = 8'h5e == io_state_in_4 ? 8'hbc : _GEN_2141; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2143 = 8'h5f == io_state_in_4 ? 8'hbe : _GEN_2142; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2144 = 8'h60 == io_state_in_4 ? 8'hc0 : _GEN_2143; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2145 = 8'h61 == io_state_in_4 ? 8'hc2 : _GEN_2144; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2146 = 8'h62 == io_state_in_4 ? 8'hc4 : _GEN_2145; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2147 = 8'h63 == io_state_in_4 ? 8'hc6 : _GEN_2146; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2148 = 8'h64 == io_state_in_4 ? 8'hc8 : _GEN_2147; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2149 = 8'h65 == io_state_in_4 ? 8'hca : _GEN_2148; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2150 = 8'h66 == io_state_in_4 ? 8'hcc : _GEN_2149; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2151 = 8'h67 == io_state_in_4 ? 8'hce : _GEN_2150; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2152 = 8'h68 == io_state_in_4 ? 8'hd0 : _GEN_2151; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2153 = 8'h69 == io_state_in_4 ? 8'hd2 : _GEN_2152; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2154 = 8'h6a == io_state_in_4 ? 8'hd4 : _GEN_2153; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2155 = 8'h6b == io_state_in_4 ? 8'hd6 : _GEN_2154; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2156 = 8'h6c == io_state_in_4 ? 8'hd8 : _GEN_2155; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2157 = 8'h6d == io_state_in_4 ? 8'hda : _GEN_2156; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2158 = 8'h6e == io_state_in_4 ? 8'hdc : _GEN_2157; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2159 = 8'h6f == io_state_in_4 ? 8'hde : _GEN_2158; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2160 = 8'h70 == io_state_in_4 ? 8'he0 : _GEN_2159; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2161 = 8'h71 == io_state_in_4 ? 8'he2 : _GEN_2160; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2162 = 8'h72 == io_state_in_4 ? 8'he4 : _GEN_2161; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2163 = 8'h73 == io_state_in_4 ? 8'he6 : _GEN_2162; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2164 = 8'h74 == io_state_in_4 ? 8'he8 : _GEN_2163; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2165 = 8'h75 == io_state_in_4 ? 8'hea : _GEN_2164; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2166 = 8'h76 == io_state_in_4 ? 8'hec : _GEN_2165; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2167 = 8'h77 == io_state_in_4 ? 8'hee : _GEN_2166; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2168 = 8'h78 == io_state_in_4 ? 8'hf0 : _GEN_2167; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2169 = 8'h79 == io_state_in_4 ? 8'hf2 : _GEN_2168; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2170 = 8'h7a == io_state_in_4 ? 8'hf4 : _GEN_2169; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2171 = 8'h7b == io_state_in_4 ? 8'hf6 : _GEN_2170; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2172 = 8'h7c == io_state_in_4 ? 8'hf8 : _GEN_2171; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2173 = 8'h7d == io_state_in_4 ? 8'hfa : _GEN_2172; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2174 = 8'h7e == io_state_in_4 ? 8'hfc : _GEN_2173; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2175 = 8'h7f == io_state_in_4 ? 8'hfe : _GEN_2174; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2176 = 8'h80 == io_state_in_4 ? 8'h1b : _GEN_2175; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2177 = 8'h81 == io_state_in_4 ? 8'h19 : _GEN_2176; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2178 = 8'h82 == io_state_in_4 ? 8'h1f : _GEN_2177; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2179 = 8'h83 == io_state_in_4 ? 8'h1d : _GEN_2178; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2180 = 8'h84 == io_state_in_4 ? 8'h13 : _GEN_2179; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2181 = 8'h85 == io_state_in_4 ? 8'h11 : _GEN_2180; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2182 = 8'h86 == io_state_in_4 ? 8'h17 : _GEN_2181; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2183 = 8'h87 == io_state_in_4 ? 8'h15 : _GEN_2182; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2184 = 8'h88 == io_state_in_4 ? 8'hb : _GEN_2183; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2185 = 8'h89 == io_state_in_4 ? 8'h9 : _GEN_2184; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2186 = 8'h8a == io_state_in_4 ? 8'hf : _GEN_2185; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2187 = 8'h8b == io_state_in_4 ? 8'hd : _GEN_2186; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2188 = 8'h8c == io_state_in_4 ? 8'h3 : _GEN_2187; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2189 = 8'h8d == io_state_in_4 ? 8'h1 : _GEN_2188; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2190 = 8'h8e == io_state_in_4 ? 8'h7 : _GEN_2189; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2191 = 8'h8f == io_state_in_4 ? 8'h5 : _GEN_2190; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2192 = 8'h90 == io_state_in_4 ? 8'h3b : _GEN_2191; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2193 = 8'h91 == io_state_in_4 ? 8'h39 : _GEN_2192; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2194 = 8'h92 == io_state_in_4 ? 8'h3f : _GEN_2193; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2195 = 8'h93 == io_state_in_4 ? 8'h3d : _GEN_2194; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2196 = 8'h94 == io_state_in_4 ? 8'h33 : _GEN_2195; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2197 = 8'h95 == io_state_in_4 ? 8'h31 : _GEN_2196; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2198 = 8'h96 == io_state_in_4 ? 8'h37 : _GEN_2197; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2199 = 8'h97 == io_state_in_4 ? 8'h35 : _GEN_2198; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2200 = 8'h98 == io_state_in_4 ? 8'h2b : _GEN_2199; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2201 = 8'h99 == io_state_in_4 ? 8'h29 : _GEN_2200; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2202 = 8'h9a == io_state_in_4 ? 8'h2f : _GEN_2201; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2203 = 8'h9b == io_state_in_4 ? 8'h2d : _GEN_2202; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2204 = 8'h9c == io_state_in_4 ? 8'h23 : _GEN_2203; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2205 = 8'h9d == io_state_in_4 ? 8'h21 : _GEN_2204; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2206 = 8'h9e == io_state_in_4 ? 8'h27 : _GEN_2205; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2207 = 8'h9f == io_state_in_4 ? 8'h25 : _GEN_2206; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2208 = 8'ha0 == io_state_in_4 ? 8'h5b : _GEN_2207; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2209 = 8'ha1 == io_state_in_4 ? 8'h59 : _GEN_2208; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2210 = 8'ha2 == io_state_in_4 ? 8'h5f : _GEN_2209; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2211 = 8'ha3 == io_state_in_4 ? 8'h5d : _GEN_2210; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2212 = 8'ha4 == io_state_in_4 ? 8'h53 : _GEN_2211; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2213 = 8'ha5 == io_state_in_4 ? 8'h51 : _GEN_2212; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2214 = 8'ha6 == io_state_in_4 ? 8'h57 : _GEN_2213; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2215 = 8'ha7 == io_state_in_4 ? 8'h55 : _GEN_2214; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2216 = 8'ha8 == io_state_in_4 ? 8'h4b : _GEN_2215; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2217 = 8'ha9 == io_state_in_4 ? 8'h49 : _GEN_2216; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2218 = 8'haa == io_state_in_4 ? 8'h4f : _GEN_2217; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2219 = 8'hab == io_state_in_4 ? 8'h4d : _GEN_2218; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2220 = 8'hac == io_state_in_4 ? 8'h43 : _GEN_2219; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2221 = 8'had == io_state_in_4 ? 8'h41 : _GEN_2220; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2222 = 8'hae == io_state_in_4 ? 8'h47 : _GEN_2221; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2223 = 8'haf == io_state_in_4 ? 8'h45 : _GEN_2222; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2224 = 8'hb0 == io_state_in_4 ? 8'h7b : _GEN_2223; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2225 = 8'hb1 == io_state_in_4 ? 8'h79 : _GEN_2224; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2226 = 8'hb2 == io_state_in_4 ? 8'h7f : _GEN_2225; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2227 = 8'hb3 == io_state_in_4 ? 8'h7d : _GEN_2226; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2228 = 8'hb4 == io_state_in_4 ? 8'h73 : _GEN_2227; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2229 = 8'hb5 == io_state_in_4 ? 8'h71 : _GEN_2228; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2230 = 8'hb6 == io_state_in_4 ? 8'h77 : _GEN_2229; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2231 = 8'hb7 == io_state_in_4 ? 8'h75 : _GEN_2230; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2232 = 8'hb8 == io_state_in_4 ? 8'h6b : _GEN_2231; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2233 = 8'hb9 == io_state_in_4 ? 8'h69 : _GEN_2232; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2234 = 8'hba == io_state_in_4 ? 8'h6f : _GEN_2233; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2235 = 8'hbb == io_state_in_4 ? 8'h6d : _GEN_2234; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2236 = 8'hbc == io_state_in_4 ? 8'h63 : _GEN_2235; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2237 = 8'hbd == io_state_in_4 ? 8'h61 : _GEN_2236; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2238 = 8'hbe == io_state_in_4 ? 8'h67 : _GEN_2237; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2239 = 8'hbf == io_state_in_4 ? 8'h65 : _GEN_2238; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2240 = 8'hc0 == io_state_in_4 ? 8'h9b : _GEN_2239; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2241 = 8'hc1 == io_state_in_4 ? 8'h99 : _GEN_2240; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2242 = 8'hc2 == io_state_in_4 ? 8'h9f : _GEN_2241; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2243 = 8'hc3 == io_state_in_4 ? 8'h9d : _GEN_2242; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2244 = 8'hc4 == io_state_in_4 ? 8'h93 : _GEN_2243; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2245 = 8'hc5 == io_state_in_4 ? 8'h91 : _GEN_2244; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2246 = 8'hc6 == io_state_in_4 ? 8'h97 : _GEN_2245; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2247 = 8'hc7 == io_state_in_4 ? 8'h95 : _GEN_2246; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2248 = 8'hc8 == io_state_in_4 ? 8'h8b : _GEN_2247; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2249 = 8'hc9 == io_state_in_4 ? 8'h89 : _GEN_2248; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2250 = 8'hca == io_state_in_4 ? 8'h8f : _GEN_2249; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2251 = 8'hcb == io_state_in_4 ? 8'h8d : _GEN_2250; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2252 = 8'hcc == io_state_in_4 ? 8'h83 : _GEN_2251; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2253 = 8'hcd == io_state_in_4 ? 8'h81 : _GEN_2252; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2254 = 8'hce == io_state_in_4 ? 8'h87 : _GEN_2253; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2255 = 8'hcf == io_state_in_4 ? 8'h85 : _GEN_2254; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2256 = 8'hd0 == io_state_in_4 ? 8'hbb : _GEN_2255; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2257 = 8'hd1 == io_state_in_4 ? 8'hb9 : _GEN_2256; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2258 = 8'hd2 == io_state_in_4 ? 8'hbf : _GEN_2257; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2259 = 8'hd3 == io_state_in_4 ? 8'hbd : _GEN_2258; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2260 = 8'hd4 == io_state_in_4 ? 8'hb3 : _GEN_2259; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2261 = 8'hd5 == io_state_in_4 ? 8'hb1 : _GEN_2260; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2262 = 8'hd6 == io_state_in_4 ? 8'hb7 : _GEN_2261; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2263 = 8'hd7 == io_state_in_4 ? 8'hb5 : _GEN_2262; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2264 = 8'hd8 == io_state_in_4 ? 8'hab : _GEN_2263; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2265 = 8'hd9 == io_state_in_4 ? 8'ha9 : _GEN_2264; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2266 = 8'hda == io_state_in_4 ? 8'haf : _GEN_2265; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2267 = 8'hdb == io_state_in_4 ? 8'had : _GEN_2266; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2268 = 8'hdc == io_state_in_4 ? 8'ha3 : _GEN_2267; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2269 = 8'hdd == io_state_in_4 ? 8'ha1 : _GEN_2268; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2270 = 8'hde == io_state_in_4 ? 8'ha7 : _GEN_2269; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2271 = 8'hdf == io_state_in_4 ? 8'ha5 : _GEN_2270; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2272 = 8'he0 == io_state_in_4 ? 8'hdb : _GEN_2271; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2273 = 8'he1 == io_state_in_4 ? 8'hd9 : _GEN_2272; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2274 = 8'he2 == io_state_in_4 ? 8'hdf : _GEN_2273; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2275 = 8'he3 == io_state_in_4 ? 8'hdd : _GEN_2274; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2276 = 8'he4 == io_state_in_4 ? 8'hd3 : _GEN_2275; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2277 = 8'he5 == io_state_in_4 ? 8'hd1 : _GEN_2276; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2278 = 8'he6 == io_state_in_4 ? 8'hd7 : _GEN_2277; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2279 = 8'he7 == io_state_in_4 ? 8'hd5 : _GEN_2278; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2280 = 8'he8 == io_state_in_4 ? 8'hcb : _GEN_2279; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2281 = 8'he9 == io_state_in_4 ? 8'hc9 : _GEN_2280; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2282 = 8'hea == io_state_in_4 ? 8'hcf : _GEN_2281; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2283 = 8'heb == io_state_in_4 ? 8'hcd : _GEN_2282; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2284 = 8'hec == io_state_in_4 ? 8'hc3 : _GEN_2283; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2285 = 8'hed == io_state_in_4 ? 8'hc1 : _GEN_2284; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2286 = 8'hee == io_state_in_4 ? 8'hc7 : _GEN_2285; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2287 = 8'hef == io_state_in_4 ? 8'hc5 : _GEN_2286; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2288 = 8'hf0 == io_state_in_4 ? 8'hfb : _GEN_2287; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2289 = 8'hf1 == io_state_in_4 ? 8'hf9 : _GEN_2288; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2290 = 8'hf2 == io_state_in_4 ? 8'hff : _GEN_2289; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2291 = 8'hf3 == io_state_in_4 ? 8'hfd : _GEN_2290; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2292 = 8'hf4 == io_state_in_4 ? 8'hf3 : _GEN_2291; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2293 = 8'hf5 == io_state_in_4 ? 8'hf1 : _GEN_2292; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2294 = 8'hf6 == io_state_in_4 ? 8'hf7 : _GEN_2293; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2295 = 8'hf7 == io_state_in_4 ? 8'hf5 : _GEN_2294; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2296 = 8'hf8 == io_state_in_4 ? 8'heb : _GEN_2295; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2297 = 8'hf9 == io_state_in_4 ? 8'he9 : _GEN_2296; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2298 = 8'hfa == io_state_in_4 ? 8'hef : _GEN_2297; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2299 = 8'hfb == io_state_in_4 ? 8'hed : _GEN_2298; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2300 = 8'hfc == io_state_in_4 ? 8'he3 : _GEN_2299; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2301 = 8'hfd == io_state_in_4 ? 8'he1 : _GEN_2300; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2302 = 8'hfe == io_state_in_4 ? 8'he7 : _GEN_2301; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2303 = 8'hff == io_state_in_4 ? 8'he5 : _GEN_2302; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2305 = 8'h1 == io_state_in_5 ? 8'h3 : 8'h0; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2306 = 8'h2 == io_state_in_5 ? 8'h6 : _GEN_2305; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2307 = 8'h3 == io_state_in_5 ? 8'h5 : _GEN_2306; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2308 = 8'h4 == io_state_in_5 ? 8'hc : _GEN_2307; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2309 = 8'h5 == io_state_in_5 ? 8'hf : _GEN_2308; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2310 = 8'h6 == io_state_in_5 ? 8'ha : _GEN_2309; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2311 = 8'h7 == io_state_in_5 ? 8'h9 : _GEN_2310; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2312 = 8'h8 == io_state_in_5 ? 8'h18 : _GEN_2311; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2313 = 8'h9 == io_state_in_5 ? 8'h1b : _GEN_2312; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2314 = 8'ha == io_state_in_5 ? 8'h1e : _GEN_2313; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2315 = 8'hb == io_state_in_5 ? 8'h1d : _GEN_2314; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2316 = 8'hc == io_state_in_5 ? 8'h14 : _GEN_2315; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2317 = 8'hd == io_state_in_5 ? 8'h17 : _GEN_2316; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2318 = 8'he == io_state_in_5 ? 8'h12 : _GEN_2317; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2319 = 8'hf == io_state_in_5 ? 8'h11 : _GEN_2318; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2320 = 8'h10 == io_state_in_5 ? 8'h30 : _GEN_2319; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2321 = 8'h11 == io_state_in_5 ? 8'h33 : _GEN_2320; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2322 = 8'h12 == io_state_in_5 ? 8'h36 : _GEN_2321; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2323 = 8'h13 == io_state_in_5 ? 8'h35 : _GEN_2322; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2324 = 8'h14 == io_state_in_5 ? 8'h3c : _GEN_2323; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2325 = 8'h15 == io_state_in_5 ? 8'h3f : _GEN_2324; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2326 = 8'h16 == io_state_in_5 ? 8'h3a : _GEN_2325; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2327 = 8'h17 == io_state_in_5 ? 8'h39 : _GEN_2326; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2328 = 8'h18 == io_state_in_5 ? 8'h28 : _GEN_2327; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2329 = 8'h19 == io_state_in_5 ? 8'h2b : _GEN_2328; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2330 = 8'h1a == io_state_in_5 ? 8'h2e : _GEN_2329; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2331 = 8'h1b == io_state_in_5 ? 8'h2d : _GEN_2330; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2332 = 8'h1c == io_state_in_5 ? 8'h24 : _GEN_2331; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2333 = 8'h1d == io_state_in_5 ? 8'h27 : _GEN_2332; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2334 = 8'h1e == io_state_in_5 ? 8'h22 : _GEN_2333; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2335 = 8'h1f == io_state_in_5 ? 8'h21 : _GEN_2334; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2336 = 8'h20 == io_state_in_5 ? 8'h60 : _GEN_2335; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2337 = 8'h21 == io_state_in_5 ? 8'h63 : _GEN_2336; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2338 = 8'h22 == io_state_in_5 ? 8'h66 : _GEN_2337; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2339 = 8'h23 == io_state_in_5 ? 8'h65 : _GEN_2338; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2340 = 8'h24 == io_state_in_5 ? 8'h6c : _GEN_2339; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2341 = 8'h25 == io_state_in_5 ? 8'h6f : _GEN_2340; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2342 = 8'h26 == io_state_in_5 ? 8'h6a : _GEN_2341; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2343 = 8'h27 == io_state_in_5 ? 8'h69 : _GEN_2342; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2344 = 8'h28 == io_state_in_5 ? 8'h78 : _GEN_2343; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2345 = 8'h29 == io_state_in_5 ? 8'h7b : _GEN_2344; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2346 = 8'h2a == io_state_in_5 ? 8'h7e : _GEN_2345; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2347 = 8'h2b == io_state_in_5 ? 8'h7d : _GEN_2346; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2348 = 8'h2c == io_state_in_5 ? 8'h74 : _GEN_2347; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2349 = 8'h2d == io_state_in_5 ? 8'h77 : _GEN_2348; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2350 = 8'h2e == io_state_in_5 ? 8'h72 : _GEN_2349; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2351 = 8'h2f == io_state_in_5 ? 8'h71 : _GEN_2350; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2352 = 8'h30 == io_state_in_5 ? 8'h50 : _GEN_2351; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2353 = 8'h31 == io_state_in_5 ? 8'h53 : _GEN_2352; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2354 = 8'h32 == io_state_in_5 ? 8'h56 : _GEN_2353; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2355 = 8'h33 == io_state_in_5 ? 8'h55 : _GEN_2354; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2356 = 8'h34 == io_state_in_5 ? 8'h5c : _GEN_2355; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2357 = 8'h35 == io_state_in_5 ? 8'h5f : _GEN_2356; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2358 = 8'h36 == io_state_in_5 ? 8'h5a : _GEN_2357; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2359 = 8'h37 == io_state_in_5 ? 8'h59 : _GEN_2358; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2360 = 8'h38 == io_state_in_5 ? 8'h48 : _GEN_2359; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2361 = 8'h39 == io_state_in_5 ? 8'h4b : _GEN_2360; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2362 = 8'h3a == io_state_in_5 ? 8'h4e : _GEN_2361; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2363 = 8'h3b == io_state_in_5 ? 8'h4d : _GEN_2362; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2364 = 8'h3c == io_state_in_5 ? 8'h44 : _GEN_2363; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2365 = 8'h3d == io_state_in_5 ? 8'h47 : _GEN_2364; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2366 = 8'h3e == io_state_in_5 ? 8'h42 : _GEN_2365; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2367 = 8'h3f == io_state_in_5 ? 8'h41 : _GEN_2366; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2368 = 8'h40 == io_state_in_5 ? 8'hc0 : _GEN_2367; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2369 = 8'h41 == io_state_in_5 ? 8'hc3 : _GEN_2368; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2370 = 8'h42 == io_state_in_5 ? 8'hc6 : _GEN_2369; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2371 = 8'h43 == io_state_in_5 ? 8'hc5 : _GEN_2370; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2372 = 8'h44 == io_state_in_5 ? 8'hcc : _GEN_2371; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2373 = 8'h45 == io_state_in_5 ? 8'hcf : _GEN_2372; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2374 = 8'h46 == io_state_in_5 ? 8'hca : _GEN_2373; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2375 = 8'h47 == io_state_in_5 ? 8'hc9 : _GEN_2374; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2376 = 8'h48 == io_state_in_5 ? 8'hd8 : _GEN_2375; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2377 = 8'h49 == io_state_in_5 ? 8'hdb : _GEN_2376; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2378 = 8'h4a == io_state_in_5 ? 8'hde : _GEN_2377; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2379 = 8'h4b == io_state_in_5 ? 8'hdd : _GEN_2378; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2380 = 8'h4c == io_state_in_5 ? 8'hd4 : _GEN_2379; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2381 = 8'h4d == io_state_in_5 ? 8'hd7 : _GEN_2380; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2382 = 8'h4e == io_state_in_5 ? 8'hd2 : _GEN_2381; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2383 = 8'h4f == io_state_in_5 ? 8'hd1 : _GEN_2382; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2384 = 8'h50 == io_state_in_5 ? 8'hf0 : _GEN_2383; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2385 = 8'h51 == io_state_in_5 ? 8'hf3 : _GEN_2384; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2386 = 8'h52 == io_state_in_5 ? 8'hf6 : _GEN_2385; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2387 = 8'h53 == io_state_in_5 ? 8'hf5 : _GEN_2386; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2388 = 8'h54 == io_state_in_5 ? 8'hfc : _GEN_2387; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2389 = 8'h55 == io_state_in_5 ? 8'hff : _GEN_2388; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2390 = 8'h56 == io_state_in_5 ? 8'hfa : _GEN_2389; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2391 = 8'h57 == io_state_in_5 ? 8'hf9 : _GEN_2390; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2392 = 8'h58 == io_state_in_5 ? 8'he8 : _GEN_2391; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2393 = 8'h59 == io_state_in_5 ? 8'heb : _GEN_2392; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2394 = 8'h5a == io_state_in_5 ? 8'hee : _GEN_2393; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2395 = 8'h5b == io_state_in_5 ? 8'hed : _GEN_2394; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2396 = 8'h5c == io_state_in_5 ? 8'he4 : _GEN_2395; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2397 = 8'h5d == io_state_in_5 ? 8'he7 : _GEN_2396; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2398 = 8'h5e == io_state_in_5 ? 8'he2 : _GEN_2397; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2399 = 8'h5f == io_state_in_5 ? 8'he1 : _GEN_2398; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2400 = 8'h60 == io_state_in_5 ? 8'ha0 : _GEN_2399; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2401 = 8'h61 == io_state_in_5 ? 8'ha3 : _GEN_2400; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2402 = 8'h62 == io_state_in_5 ? 8'ha6 : _GEN_2401; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2403 = 8'h63 == io_state_in_5 ? 8'ha5 : _GEN_2402; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2404 = 8'h64 == io_state_in_5 ? 8'hac : _GEN_2403; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2405 = 8'h65 == io_state_in_5 ? 8'haf : _GEN_2404; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2406 = 8'h66 == io_state_in_5 ? 8'haa : _GEN_2405; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2407 = 8'h67 == io_state_in_5 ? 8'ha9 : _GEN_2406; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2408 = 8'h68 == io_state_in_5 ? 8'hb8 : _GEN_2407; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2409 = 8'h69 == io_state_in_5 ? 8'hbb : _GEN_2408; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2410 = 8'h6a == io_state_in_5 ? 8'hbe : _GEN_2409; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2411 = 8'h6b == io_state_in_5 ? 8'hbd : _GEN_2410; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2412 = 8'h6c == io_state_in_5 ? 8'hb4 : _GEN_2411; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2413 = 8'h6d == io_state_in_5 ? 8'hb7 : _GEN_2412; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2414 = 8'h6e == io_state_in_5 ? 8'hb2 : _GEN_2413; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2415 = 8'h6f == io_state_in_5 ? 8'hb1 : _GEN_2414; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2416 = 8'h70 == io_state_in_5 ? 8'h90 : _GEN_2415; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2417 = 8'h71 == io_state_in_5 ? 8'h93 : _GEN_2416; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2418 = 8'h72 == io_state_in_5 ? 8'h96 : _GEN_2417; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2419 = 8'h73 == io_state_in_5 ? 8'h95 : _GEN_2418; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2420 = 8'h74 == io_state_in_5 ? 8'h9c : _GEN_2419; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2421 = 8'h75 == io_state_in_5 ? 8'h9f : _GEN_2420; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2422 = 8'h76 == io_state_in_5 ? 8'h9a : _GEN_2421; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2423 = 8'h77 == io_state_in_5 ? 8'h99 : _GEN_2422; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2424 = 8'h78 == io_state_in_5 ? 8'h88 : _GEN_2423; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2425 = 8'h79 == io_state_in_5 ? 8'h8b : _GEN_2424; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2426 = 8'h7a == io_state_in_5 ? 8'h8e : _GEN_2425; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2427 = 8'h7b == io_state_in_5 ? 8'h8d : _GEN_2426; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2428 = 8'h7c == io_state_in_5 ? 8'h84 : _GEN_2427; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2429 = 8'h7d == io_state_in_5 ? 8'h87 : _GEN_2428; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2430 = 8'h7e == io_state_in_5 ? 8'h82 : _GEN_2429; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2431 = 8'h7f == io_state_in_5 ? 8'h81 : _GEN_2430; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2432 = 8'h80 == io_state_in_5 ? 8'h9b : _GEN_2431; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2433 = 8'h81 == io_state_in_5 ? 8'h98 : _GEN_2432; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2434 = 8'h82 == io_state_in_5 ? 8'h9d : _GEN_2433; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2435 = 8'h83 == io_state_in_5 ? 8'h9e : _GEN_2434; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2436 = 8'h84 == io_state_in_5 ? 8'h97 : _GEN_2435; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2437 = 8'h85 == io_state_in_5 ? 8'h94 : _GEN_2436; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2438 = 8'h86 == io_state_in_5 ? 8'h91 : _GEN_2437; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2439 = 8'h87 == io_state_in_5 ? 8'h92 : _GEN_2438; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2440 = 8'h88 == io_state_in_5 ? 8'h83 : _GEN_2439; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2441 = 8'h89 == io_state_in_5 ? 8'h80 : _GEN_2440; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2442 = 8'h8a == io_state_in_5 ? 8'h85 : _GEN_2441; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2443 = 8'h8b == io_state_in_5 ? 8'h86 : _GEN_2442; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2444 = 8'h8c == io_state_in_5 ? 8'h8f : _GEN_2443; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2445 = 8'h8d == io_state_in_5 ? 8'h8c : _GEN_2444; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2446 = 8'h8e == io_state_in_5 ? 8'h89 : _GEN_2445; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2447 = 8'h8f == io_state_in_5 ? 8'h8a : _GEN_2446; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2448 = 8'h90 == io_state_in_5 ? 8'hab : _GEN_2447; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2449 = 8'h91 == io_state_in_5 ? 8'ha8 : _GEN_2448; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2450 = 8'h92 == io_state_in_5 ? 8'had : _GEN_2449; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2451 = 8'h93 == io_state_in_5 ? 8'hae : _GEN_2450; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2452 = 8'h94 == io_state_in_5 ? 8'ha7 : _GEN_2451; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2453 = 8'h95 == io_state_in_5 ? 8'ha4 : _GEN_2452; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2454 = 8'h96 == io_state_in_5 ? 8'ha1 : _GEN_2453; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2455 = 8'h97 == io_state_in_5 ? 8'ha2 : _GEN_2454; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2456 = 8'h98 == io_state_in_5 ? 8'hb3 : _GEN_2455; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2457 = 8'h99 == io_state_in_5 ? 8'hb0 : _GEN_2456; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2458 = 8'h9a == io_state_in_5 ? 8'hb5 : _GEN_2457; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2459 = 8'h9b == io_state_in_5 ? 8'hb6 : _GEN_2458; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2460 = 8'h9c == io_state_in_5 ? 8'hbf : _GEN_2459; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2461 = 8'h9d == io_state_in_5 ? 8'hbc : _GEN_2460; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2462 = 8'h9e == io_state_in_5 ? 8'hb9 : _GEN_2461; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2463 = 8'h9f == io_state_in_5 ? 8'hba : _GEN_2462; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2464 = 8'ha0 == io_state_in_5 ? 8'hfb : _GEN_2463; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2465 = 8'ha1 == io_state_in_5 ? 8'hf8 : _GEN_2464; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2466 = 8'ha2 == io_state_in_5 ? 8'hfd : _GEN_2465; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2467 = 8'ha3 == io_state_in_5 ? 8'hfe : _GEN_2466; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2468 = 8'ha4 == io_state_in_5 ? 8'hf7 : _GEN_2467; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2469 = 8'ha5 == io_state_in_5 ? 8'hf4 : _GEN_2468; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2470 = 8'ha6 == io_state_in_5 ? 8'hf1 : _GEN_2469; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2471 = 8'ha7 == io_state_in_5 ? 8'hf2 : _GEN_2470; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2472 = 8'ha8 == io_state_in_5 ? 8'he3 : _GEN_2471; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2473 = 8'ha9 == io_state_in_5 ? 8'he0 : _GEN_2472; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2474 = 8'haa == io_state_in_5 ? 8'he5 : _GEN_2473; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2475 = 8'hab == io_state_in_5 ? 8'he6 : _GEN_2474; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2476 = 8'hac == io_state_in_5 ? 8'hef : _GEN_2475; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2477 = 8'had == io_state_in_5 ? 8'hec : _GEN_2476; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2478 = 8'hae == io_state_in_5 ? 8'he9 : _GEN_2477; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2479 = 8'haf == io_state_in_5 ? 8'hea : _GEN_2478; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2480 = 8'hb0 == io_state_in_5 ? 8'hcb : _GEN_2479; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2481 = 8'hb1 == io_state_in_5 ? 8'hc8 : _GEN_2480; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2482 = 8'hb2 == io_state_in_5 ? 8'hcd : _GEN_2481; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2483 = 8'hb3 == io_state_in_5 ? 8'hce : _GEN_2482; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2484 = 8'hb4 == io_state_in_5 ? 8'hc7 : _GEN_2483; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2485 = 8'hb5 == io_state_in_5 ? 8'hc4 : _GEN_2484; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2486 = 8'hb6 == io_state_in_5 ? 8'hc1 : _GEN_2485; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2487 = 8'hb7 == io_state_in_5 ? 8'hc2 : _GEN_2486; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2488 = 8'hb8 == io_state_in_5 ? 8'hd3 : _GEN_2487; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2489 = 8'hb9 == io_state_in_5 ? 8'hd0 : _GEN_2488; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2490 = 8'hba == io_state_in_5 ? 8'hd5 : _GEN_2489; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2491 = 8'hbb == io_state_in_5 ? 8'hd6 : _GEN_2490; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2492 = 8'hbc == io_state_in_5 ? 8'hdf : _GEN_2491; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2493 = 8'hbd == io_state_in_5 ? 8'hdc : _GEN_2492; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2494 = 8'hbe == io_state_in_5 ? 8'hd9 : _GEN_2493; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2495 = 8'hbf == io_state_in_5 ? 8'hda : _GEN_2494; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2496 = 8'hc0 == io_state_in_5 ? 8'h5b : _GEN_2495; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2497 = 8'hc1 == io_state_in_5 ? 8'h58 : _GEN_2496; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2498 = 8'hc2 == io_state_in_5 ? 8'h5d : _GEN_2497; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2499 = 8'hc3 == io_state_in_5 ? 8'h5e : _GEN_2498; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2500 = 8'hc4 == io_state_in_5 ? 8'h57 : _GEN_2499; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2501 = 8'hc5 == io_state_in_5 ? 8'h54 : _GEN_2500; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2502 = 8'hc6 == io_state_in_5 ? 8'h51 : _GEN_2501; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2503 = 8'hc7 == io_state_in_5 ? 8'h52 : _GEN_2502; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2504 = 8'hc8 == io_state_in_5 ? 8'h43 : _GEN_2503; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2505 = 8'hc9 == io_state_in_5 ? 8'h40 : _GEN_2504; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2506 = 8'hca == io_state_in_5 ? 8'h45 : _GEN_2505; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2507 = 8'hcb == io_state_in_5 ? 8'h46 : _GEN_2506; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2508 = 8'hcc == io_state_in_5 ? 8'h4f : _GEN_2507; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2509 = 8'hcd == io_state_in_5 ? 8'h4c : _GEN_2508; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2510 = 8'hce == io_state_in_5 ? 8'h49 : _GEN_2509; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2511 = 8'hcf == io_state_in_5 ? 8'h4a : _GEN_2510; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2512 = 8'hd0 == io_state_in_5 ? 8'h6b : _GEN_2511; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2513 = 8'hd1 == io_state_in_5 ? 8'h68 : _GEN_2512; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2514 = 8'hd2 == io_state_in_5 ? 8'h6d : _GEN_2513; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2515 = 8'hd3 == io_state_in_5 ? 8'h6e : _GEN_2514; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2516 = 8'hd4 == io_state_in_5 ? 8'h67 : _GEN_2515; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2517 = 8'hd5 == io_state_in_5 ? 8'h64 : _GEN_2516; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2518 = 8'hd6 == io_state_in_5 ? 8'h61 : _GEN_2517; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2519 = 8'hd7 == io_state_in_5 ? 8'h62 : _GEN_2518; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2520 = 8'hd8 == io_state_in_5 ? 8'h73 : _GEN_2519; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2521 = 8'hd9 == io_state_in_5 ? 8'h70 : _GEN_2520; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2522 = 8'hda == io_state_in_5 ? 8'h75 : _GEN_2521; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2523 = 8'hdb == io_state_in_5 ? 8'h76 : _GEN_2522; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2524 = 8'hdc == io_state_in_5 ? 8'h7f : _GEN_2523; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2525 = 8'hdd == io_state_in_5 ? 8'h7c : _GEN_2524; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2526 = 8'hde == io_state_in_5 ? 8'h79 : _GEN_2525; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2527 = 8'hdf == io_state_in_5 ? 8'h7a : _GEN_2526; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2528 = 8'he0 == io_state_in_5 ? 8'h3b : _GEN_2527; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2529 = 8'he1 == io_state_in_5 ? 8'h38 : _GEN_2528; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2530 = 8'he2 == io_state_in_5 ? 8'h3d : _GEN_2529; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2531 = 8'he3 == io_state_in_5 ? 8'h3e : _GEN_2530; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2532 = 8'he4 == io_state_in_5 ? 8'h37 : _GEN_2531; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2533 = 8'he5 == io_state_in_5 ? 8'h34 : _GEN_2532; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2534 = 8'he6 == io_state_in_5 ? 8'h31 : _GEN_2533; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2535 = 8'he7 == io_state_in_5 ? 8'h32 : _GEN_2534; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2536 = 8'he8 == io_state_in_5 ? 8'h23 : _GEN_2535; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2537 = 8'he9 == io_state_in_5 ? 8'h20 : _GEN_2536; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2538 = 8'hea == io_state_in_5 ? 8'h25 : _GEN_2537; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2539 = 8'heb == io_state_in_5 ? 8'h26 : _GEN_2538; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2540 = 8'hec == io_state_in_5 ? 8'h2f : _GEN_2539; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2541 = 8'hed == io_state_in_5 ? 8'h2c : _GEN_2540; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2542 = 8'hee == io_state_in_5 ? 8'h29 : _GEN_2541; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2543 = 8'hef == io_state_in_5 ? 8'h2a : _GEN_2542; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2544 = 8'hf0 == io_state_in_5 ? 8'hb : _GEN_2543; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2545 = 8'hf1 == io_state_in_5 ? 8'h8 : _GEN_2544; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2546 = 8'hf2 == io_state_in_5 ? 8'hd : _GEN_2545; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2547 = 8'hf3 == io_state_in_5 ? 8'he : _GEN_2546; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2548 = 8'hf4 == io_state_in_5 ? 8'h7 : _GEN_2547; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2549 = 8'hf5 == io_state_in_5 ? 8'h4 : _GEN_2548; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2550 = 8'hf6 == io_state_in_5 ? 8'h1 : _GEN_2549; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2551 = 8'hf7 == io_state_in_5 ? 8'h2 : _GEN_2550; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2552 = 8'hf8 == io_state_in_5 ? 8'h13 : _GEN_2551; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2553 = 8'hf9 == io_state_in_5 ? 8'h10 : _GEN_2552; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2554 = 8'hfa == io_state_in_5 ? 8'h15 : _GEN_2553; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2555 = 8'hfb == io_state_in_5 ? 8'h16 : _GEN_2554; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2556 = 8'hfc == io_state_in_5 ? 8'h1f : _GEN_2555; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2557 = 8'hfd == io_state_in_5 ? 8'h1c : _GEN_2556; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2558 = 8'hfe == io_state_in_5 ? 8'h19 : _GEN_2557; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _GEN_2559 = 8'hff == io_state_in_5 ? 8'h1a : _GEN_2558; // @[MixColumns.scala 130:{41,41}]
  wire [7:0] _tmp_state_4_T = _GEN_2303 ^ _GEN_2559; // @[MixColumns.scala 130:41]
  wire [7:0] _tmp_state_4_T_1 = _tmp_state_4_T ^ io_state_in_6; // @[MixColumns.scala 130:65]
  wire [7:0] _GEN_2561 = 8'h1 == io_state_in_5 ? 8'h2 : 8'h0; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2562 = 8'h2 == io_state_in_5 ? 8'h4 : _GEN_2561; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2563 = 8'h3 == io_state_in_5 ? 8'h6 : _GEN_2562; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2564 = 8'h4 == io_state_in_5 ? 8'h8 : _GEN_2563; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2565 = 8'h5 == io_state_in_5 ? 8'ha : _GEN_2564; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2566 = 8'h6 == io_state_in_5 ? 8'hc : _GEN_2565; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2567 = 8'h7 == io_state_in_5 ? 8'he : _GEN_2566; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2568 = 8'h8 == io_state_in_5 ? 8'h10 : _GEN_2567; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2569 = 8'h9 == io_state_in_5 ? 8'h12 : _GEN_2568; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2570 = 8'ha == io_state_in_5 ? 8'h14 : _GEN_2569; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2571 = 8'hb == io_state_in_5 ? 8'h16 : _GEN_2570; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2572 = 8'hc == io_state_in_5 ? 8'h18 : _GEN_2571; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2573 = 8'hd == io_state_in_5 ? 8'h1a : _GEN_2572; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2574 = 8'he == io_state_in_5 ? 8'h1c : _GEN_2573; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2575 = 8'hf == io_state_in_5 ? 8'h1e : _GEN_2574; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2576 = 8'h10 == io_state_in_5 ? 8'h20 : _GEN_2575; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2577 = 8'h11 == io_state_in_5 ? 8'h22 : _GEN_2576; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2578 = 8'h12 == io_state_in_5 ? 8'h24 : _GEN_2577; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2579 = 8'h13 == io_state_in_5 ? 8'h26 : _GEN_2578; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2580 = 8'h14 == io_state_in_5 ? 8'h28 : _GEN_2579; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2581 = 8'h15 == io_state_in_5 ? 8'h2a : _GEN_2580; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2582 = 8'h16 == io_state_in_5 ? 8'h2c : _GEN_2581; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2583 = 8'h17 == io_state_in_5 ? 8'h2e : _GEN_2582; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2584 = 8'h18 == io_state_in_5 ? 8'h30 : _GEN_2583; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2585 = 8'h19 == io_state_in_5 ? 8'h32 : _GEN_2584; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2586 = 8'h1a == io_state_in_5 ? 8'h34 : _GEN_2585; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2587 = 8'h1b == io_state_in_5 ? 8'h36 : _GEN_2586; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2588 = 8'h1c == io_state_in_5 ? 8'h38 : _GEN_2587; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2589 = 8'h1d == io_state_in_5 ? 8'h3a : _GEN_2588; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2590 = 8'h1e == io_state_in_5 ? 8'h3c : _GEN_2589; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2591 = 8'h1f == io_state_in_5 ? 8'h3e : _GEN_2590; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2592 = 8'h20 == io_state_in_5 ? 8'h40 : _GEN_2591; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2593 = 8'h21 == io_state_in_5 ? 8'h42 : _GEN_2592; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2594 = 8'h22 == io_state_in_5 ? 8'h44 : _GEN_2593; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2595 = 8'h23 == io_state_in_5 ? 8'h46 : _GEN_2594; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2596 = 8'h24 == io_state_in_5 ? 8'h48 : _GEN_2595; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2597 = 8'h25 == io_state_in_5 ? 8'h4a : _GEN_2596; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2598 = 8'h26 == io_state_in_5 ? 8'h4c : _GEN_2597; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2599 = 8'h27 == io_state_in_5 ? 8'h4e : _GEN_2598; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2600 = 8'h28 == io_state_in_5 ? 8'h50 : _GEN_2599; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2601 = 8'h29 == io_state_in_5 ? 8'h52 : _GEN_2600; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2602 = 8'h2a == io_state_in_5 ? 8'h54 : _GEN_2601; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2603 = 8'h2b == io_state_in_5 ? 8'h56 : _GEN_2602; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2604 = 8'h2c == io_state_in_5 ? 8'h58 : _GEN_2603; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2605 = 8'h2d == io_state_in_5 ? 8'h5a : _GEN_2604; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2606 = 8'h2e == io_state_in_5 ? 8'h5c : _GEN_2605; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2607 = 8'h2f == io_state_in_5 ? 8'h5e : _GEN_2606; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2608 = 8'h30 == io_state_in_5 ? 8'h60 : _GEN_2607; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2609 = 8'h31 == io_state_in_5 ? 8'h62 : _GEN_2608; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2610 = 8'h32 == io_state_in_5 ? 8'h64 : _GEN_2609; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2611 = 8'h33 == io_state_in_5 ? 8'h66 : _GEN_2610; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2612 = 8'h34 == io_state_in_5 ? 8'h68 : _GEN_2611; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2613 = 8'h35 == io_state_in_5 ? 8'h6a : _GEN_2612; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2614 = 8'h36 == io_state_in_5 ? 8'h6c : _GEN_2613; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2615 = 8'h37 == io_state_in_5 ? 8'h6e : _GEN_2614; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2616 = 8'h38 == io_state_in_5 ? 8'h70 : _GEN_2615; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2617 = 8'h39 == io_state_in_5 ? 8'h72 : _GEN_2616; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2618 = 8'h3a == io_state_in_5 ? 8'h74 : _GEN_2617; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2619 = 8'h3b == io_state_in_5 ? 8'h76 : _GEN_2618; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2620 = 8'h3c == io_state_in_5 ? 8'h78 : _GEN_2619; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2621 = 8'h3d == io_state_in_5 ? 8'h7a : _GEN_2620; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2622 = 8'h3e == io_state_in_5 ? 8'h7c : _GEN_2621; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2623 = 8'h3f == io_state_in_5 ? 8'h7e : _GEN_2622; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2624 = 8'h40 == io_state_in_5 ? 8'h80 : _GEN_2623; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2625 = 8'h41 == io_state_in_5 ? 8'h82 : _GEN_2624; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2626 = 8'h42 == io_state_in_5 ? 8'h84 : _GEN_2625; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2627 = 8'h43 == io_state_in_5 ? 8'h86 : _GEN_2626; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2628 = 8'h44 == io_state_in_5 ? 8'h88 : _GEN_2627; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2629 = 8'h45 == io_state_in_5 ? 8'h8a : _GEN_2628; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2630 = 8'h46 == io_state_in_5 ? 8'h8c : _GEN_2629; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2631 = 8'h47 == io_state_in_5 ? 8'h8e : _GEN_2630; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2632 = 8'h48 == io_state_in_5 ? 8'h90 : _GEN_2631; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2633 = 8'h49 == io_state_in_5 ? 8'h92 : _GEN_2632; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2634 = 8'h4a == io_state_in_5 ? 8'h94 : _GEN_2633; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2635 = 8'h4b == io_state_in_5 ? 8'h96 : _GEN_2634; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2636 = 8'h4c == io_state_in_5 ? 8'h98 : _GEN_2635; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2637 = 8'h4d == io_state_in_5 ? 8'h9a : _GEN_2636; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2638 = 8'h4e == io_state_in_5 ? 8'h9c : _GEN_2637; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2639 = 8'h4f == io_state_in_5 ? 8'h9e : _GEN_2638; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2640 = 8'h50 == io_state_in_5 ? 8'ha0 : _GEN_2639; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2641 = 8'h51 == io_state_in_5 ? 8'ha2 : _GEN_2640; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2642 = 8'h52 == io_state_in_5 ? 8'ha4 : _GEN_2641; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2643 = 8'h53 == io_state_in_5 ? 8'ha6 : _GEN_2642; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2644 = 8'h54 == io_state_in_5 ? 8'ha8 : _GEN_2643; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2645 = 8'h55 == io_state_in_5 ? 8'haa : _GEN_2644; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2646 = 8'h56 == io_state_in_5 ? 8'hac : _GEN_2645; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2647 = 8'h57 == io_state_in_5 ? 8'hae : _GEN_2646; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2648 = 8'h58 == io_state_in_5 ? 8'hb0 : _GEN_2647; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2649 = 8'h59 == io_state_in_5 ? 8'hb2 : _GEN_2648; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2650 = 8'h5a == io_state_in_5 ? 8'hb4 : _GEN_2649; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2651 = 8'h5b == io_state_in_5 ? 8'hb6 : _GEN_2650; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2652 = 8'h5c == io_state_in_5 ? 8'hb8 : _GEN_2651; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2653 = 8'h5d == io_state_in_5 ? 8'hba : _GEN_2652; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2654 = 8'h5e == io_state_in_5 ? 8'hbc : _GEN_2653; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2655 = 8'h5f == io_state_in_5 ? 8'hbe : _GEN_2654; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2656 = 8'h60 == io_state_in_5 ? 8'hc0 : _GEN_2655; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2657 = 8'h61 == io_state_in_5 ? 8'hc2 : _GEN_2656; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2658 = 8'h62 == io_state_in_5 ? 8'hc4 : _GEN_2657; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2659 = 8'h63 == io_state_in_5 ? 8'hc6 : _GEN_2658; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2660 = 8'h64 == io_state_in_5 ? 8'hc8 : _GEN_2659; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2661 = 8'h65 == io_state_in_5 ? 8'hca : _GEN_2660; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2662 = 8'h66 == io_state_in_5 ? 8'hcc : _GEN_2661; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2663 = 8'h67 == io_state_in_5 ? 8'hce : _GEN_2662; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2664 = 8'h68 == io_state_in_5 ? 8'hd0 : _GEN_2663; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2665 = 8'h69 == io_state_in_5 ? 8'hd2 : _GEN_2664; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2666 = 8'h6a == io_state_in_5 ? 8'hd4 : _GEN_2665; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2667 = 8'h6b == io_state_in_5 ? 8'hd6 : _GEN_2666; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2668 = 8'h6c == io_state_in_5 ? 8'hd8 : _GEN_2667; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2669 = 8'h6d == io_state_in_5 ? 8'hda : _GEN_2668; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2670 = 8'h6e == io_state_in_5 ? 8'hdc : _GEN_2669; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2671 = 8'h6f == io_state_in_5 ? 8'hde : _GEN_2670; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2672 = 8'h70 == io_state_in_5 ? 8'he0 : _GEN_2671; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2673 = 8'h71 == io_state_in_5 ? 8'he2 : _GEN_2672; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2674 = 8'h72 == io_state_in_5 ? 8'he4 : _GEN_2673; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2675 = 8'h73 == io_state_in_5 ? 8'he6 : _GEN_2674; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2676 = 8'h74 == io_state_in_5 ? 8'he8 : _GEN_2675; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2677 = 8'h75 == io_state_in_5 ? 8'hea : _GEN_2676; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2678 = 8'h76 == io_state_in_5 ? 8'hec : _GEN_2677; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2679 = 8'h77 == io_state_in_5 ? 8'hee : _GEN_2678; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2680 = 8'h78 == io_state_in_5 ? 8'hf0 : _GEN_2679; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2681 = 8'h79 == io_state_in_5 ? 8'hf2 : _GEN_2680; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2682 = 8'h7a == io_state_in_5 ? 8'hf4 : _GEN_2681; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2683 = 8'h7b == io_state_in_5 ? 8'hf6 : _GEN_2682; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2684 = 8'h7c == io_state_in_5 ? 8'hf8 : _GEN_2683; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2685 = 8'h7d == io_state_in_5 ? 8'hfa : _GEN_2684; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2686 = 8'h7e == io_state_in_5 ? 8'hfc : _GEN_2685; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2687 = 8'h7f == io_state_in_5 ? 8'hfe : _GEN_2686; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2688 = 8'h80 == io_state_in_5 ? 8'h1b : _GEN_2687; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2689 = 8'h81 == io_state_in_5 ? 8'h19 : _GEN_2688; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2690 = 8'h82 == io_state_in_5 ? 8'h1f : _GEN_2689; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2691 = 8'h83 == io_state_in_5 ? 8'h1d : _GEN_2690; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2692 = 8'h84 == io_state_in_5 ? 8'h13 : _GEN_2691; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2693 = 8'h85 == io_state_in_5 ? 8'h11 : _GEN_2692; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2694 = 8'h86 == io_state_in_5 ? 8'h17 : _GEN_2693; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2695 = 8'h87 == io_state_in_5 ? 8'h15 : _GEN_2694; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2696 = 8'h88 == io_state_in_5 ? 8'hb : _GEN_2695; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2697 = 8'h89 == io_state_in_5 ? 8'h9 : _GEN_2696; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2698 = 8'h8a == io_state_in_5 ? 8'hf : _GEN_2697; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2699 = 8'h8b == io_state_in_5 ? 8'hd : _GEN_2698; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2700 = 8'h8c == io_state_in_5 ? 8'h3 : _GEN_2699; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2701 = 8'h8d == io_state_in_5 ? 8'h1 : _GEN_2700; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2702 = 8'h8e == io_state_in_5 ? 8'h7 : _GEN_2701; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2703 = 8'h8f == io_state_in_5 ? 8'h5 : _GEN_2702; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2704 = 8'h90 == io_state_in_5 ? 8'h3b : _GEN_2703; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2705 = 8'h91 == io_state_in_5 ? 8'h39 : _GEN_2704; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2706 = 8'h92 == io_state_in_5 ? 8'h3f : _GEN_2705; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2707 = 8'h93 == io_state_in_5 ? 8'h3d : _GEN_2706; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2708 = 8'h94 == io_state_in_5 ? 8'h33 : _GEN_2707; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2709 = 8'h95 == io_state_in_5 ? 8'h31 : _GEN_2708; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2710 = 8'h96 == io_state_in_5 ? 8'h37 : _GEN_2709; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2711 = 8'h97 == io_state_in_5 ? 8'h35 : _GEN_2710; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2712 = 8'h98 == io_state_in_5 ? 8'h2b : _GEN_2711; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2713 = 8'h99 == io_state_in_5 ? 8'h29 : _GEN_2712; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2714 = 8'h9a == io_state_in_5 ? 8'h2f : _GEN_2713; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2715 = 8'h9b == io_state_in_5 ? 8'h2d : _GEN_2714; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2716 = 8'h9c == io_state_in_5 ? 8'h23 : _GEN_2715; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2717 = 8'h9d == io_state_in_5 ? 8'h21 : _GEN_2716; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2718 = 8'h9e == io_state_in_5 ? 8'h27 : _GEN_2717; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2719 = 8'h9f == io_state_in_5 ? 8'h25 : _GEN_2718; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2720 = 8'ha0 == io_state_in_5 ? 8'h5b : _GEN_2719; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2721 = 8'ha1 == io_state_in_5 ? 8'h59 : _GEN_2720; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2722 = 8'ha2 == io_state_in_5 ? 8'h5f : _GEN_2721; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2723 = 8'ha3 == io_state_in_5 ? 8'h5d : _GEN_2722; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2724 = 8'ha4 == io_state_in_5 ? 8'h53 : _GEN_2723; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2725 = 8'ha5 == io_state_in_5 ? 8'h51 : _GEN_2724; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2726 = 8'ha6 == io_state_in_5 ? 8'h57 : _GEN_2725; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2727 = 8'ha7 == io_state_in_5 ? 8'h55 : _GEN_2726; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2728 = 8'ha8 == io_state_in_5 ? 8'h4b : _GEN_2727; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2729 = 8'ha9 == io_state_in_5 ? 8'h49 : _GEN_2728; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2730 = 8'haa == io_state_in_5 ? 8'h4f : _GEN_2729; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2731 = 8'hab == io_state_in_5 ? 8'h4d : _GEN_2730; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2732 = 8'hac == io_state_in_5 ? 8'h43 : _GEN_2731; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2733 = 8'had == io_state_in_5 ? 8'h41 : _GEN_2732; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2734 = 8'hae == io_state_in_5 ? 8'h47 : _GEN_2733; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2735 = 8'haf == io_state_in_5 ? 8'h45 : _GEN_2734; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2736 = 8'hb0 == io_state_in_5 ? 8'h7b : _GEN_2735; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2737 = 8'hb1 == io_state_in_5 ? 8'h79 : _GEN_2736; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2738 = 8'hb2 == io_state_in_5 ? 8'h7f : _GEN_2737; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2739 = 8'hb3 == io_state_in_5 ? 8'h7d : _GEN_2738; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2740 = 8'hb4 == io_state_in_5 ? 8'h73 : _GEN_2739; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2741 = 8'hb5 == io_state_in_5 ? 8'h71 : _GEN_2740; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2742 = 8'hb6 == io_state_in_5 ? 8'h77 : _GEN_2741; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2743 = 8'hb7 == io_state_in_5 ? 8'h75 : _GEN_2742; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2744 = 8'hb8 == io_state_in_5 ? 8'h6b : _GEN_2743; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2745 = 8'hb9 == io_state_in_5 ? 8'h69 : _GEN_2744; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2746 = 8'hba == io_state_in_5 ? 8'h6f : _GEN_2745; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2747 = 8'hbb == io_state_in_5 ? 8'h6d : _GEN_2746; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2748 = 8'hbc == io_state_in_5 ? 8'h63 : _GEN_2747; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2749 = 8'hbd == io_state_in_5 ? 8'h61 : _GEN_2748; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2750 = 8'hbe == io_state_in_5 ? 8'h67 : _GEN_2749; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2751 = 8'hbf == io_state_in_5 ? 8'h65 : _GEN_2750; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2752 = 8'hc0 == io_state_in_5 ? 8'h9b : _GEN_2751; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2753 = 8'hc1 == io_state_in_5 ? 8'h99 : _GEN_2752; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2754 = 8'hc2 == io_state_in_5 ? 8'h9f : _GEN_2753; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2755 = 8'hc3 == io_state_in_5 ? 8'h9d : _GEN_2754; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2756 = 8'hc4 == io_state_in_5 ? 8'h93 : _GEN_2755; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2757 = 8'hc5 == io_state_in_5 ? 8'h91 : _GEN_2756; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2758 = 8'hc6 == io_state_in_5 ? 8'h97 : _GEN_2757; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2759 = 8'hc7 == io_state_in_5 ? 8'h95 : _GEN_2758; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2760 = 8'hc8 == io_state_in_5 ? 8'h8b : _GEN_2759; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2761 = 8'hc9 == io_state_in_5 ? 8'h89 : _GEN_2760; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2762 = 8'hca == io_state_in_5 ? 8'h8f : _GEN_2761; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2763 = 8'hcb == io_state_in_5 ? 8'h8d : _GEN_2762; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2764 = 8'hcc == io_state_in_5 ? 8'h83 : _GEN_2763; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2765 = 8'hcd == io_state_in_5 ? 8'h81 : _GEN_2764; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2766 = 8'hce == io_state_in_5 ? 8'h87 : _GEN_2765; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2767 = 8'hcf == io_state_in_5 ? 8'h85 : _GEN_2766; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2768 = 8'hd0 == io_state_in_5 ? 8'hbb : _GEN_2767; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2769 = 8'hd1 == io_state_in_5 ? 8'hb9 : _GEN_2768; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2770 = 8'hd2 == io_state_in_5 ? 8'hbf : _GEN_2769; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2771 = 8'hd3 == io_state_in_5 ? 8'hbd : _GEN_2770; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2772 = 8'hd4 == io_state_in_5 ? 8'hb3 : _GEN_2771; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2773 = 8'hd5 == io_state_in_5 ? 8'hb1 : _GEN_2772; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2774 = 8'hd6 == io_state_in_5 ? 8'hb7 : _GEN_2773; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2775 = 8'hd7 == io_state_in_5 ? 8'hb5 : _GEN_2774; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2776 = 8'hd8 == io_state_in_5 ? 8'hab : _GEN_2775; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2777 = 8'hd9 == io_state_in_5 ? 8'ha9 : _GEN_2776; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2778 = 8'hda == io_state_in_5 ? 8'haf : _GEN_2777; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2779 = 8'hdb == io_state_in_5 ? 8'had : _GEN_2778; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2780 = 8'hdc == io_state_in_5 ? 8'ha3 : _GEN_2779; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2781 = 8'hdd == io_state_in_5 ? 8'ha1 : _GEN_2780; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2782 = 8'hde == io_state_in_5 ? 8'ha7 : _GEN_2781; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2783 = 8'hdf == io_state_in_5 ? 8'ha5 : _GEN_2782; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2784 = 8'he0 == io_state_in_5 ? 8'hdb : _GEN_2783; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2785 = 8'he1 == io_state_in_5 ? 8'hd9 : _GEN_2784; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2786 = 8'he2 == io_state_in_5 ? 8'hdf : _GEN_2785; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2787 = 8'he3 == io_state_in_5 ? 8'hdd : _GEN_2786; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2788 = 8'he4 == io_state_in_5 ? 8'hd3 : _GEN_2787; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2789 = 8'he5 == io_state_in_5 ? 8'hd1 : _GEN_2788; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2790 = 8'he6 == io_state_in_5 ? 8'hd7 : _GEN_2789; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2791 = 8'he7 == io_state_in_5 ? 8'hd5 : _GEN_2790; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2792 = 8'he8 == io_state_in_5 ? 8'hcb : _GEN_2791; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2793 = 8'he9 == io_state_in_5 ? 8'hc9 : _GEN_2792; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2794 = 8'hea == io_state_in_5 ? 8'hcf : _GEN_2793; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2795 = 8'heb == io_state_in_5 ? 8'hcd : _GEN_2794; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2796 = 8'hec == io_state_in_5 ? 8'hc3 : _GEN_2795; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2797 = 8'hed == io_state_in_5 ? 8'hc1 : _GEN_2796; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2798 = 8'hee == io_state_in_5 ? 8'hc7 : _GEN_2797; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2799 = 8'hef == io_state_in_5 ? 8'hc5 : _GEN_2798; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2800 = 8'hf0 == io_state_in_5 ? 8'hfb : _GEN_2799; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2801 = 8'hf1 == io_state_in_5 ? 8'hf9 : _GEN_2800; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2802 = 8'hf2 == io_state_in_5 ? 8'hff : _GEN_2801; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2803 = 8'hf3 == io_state_in_5 ? 8'hfd : _GEN_2802; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2804 = 8'hf4 == io_state_in_5 ? 8'hf3 : _GEN_2803; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2805 = 8'hf5 == io_state_in_5 ? 8'hf1 : _GEN_2804; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2806 = 8'hf6 == io_state_in_5 ? 8'hf7 : _GEN_2805; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2807 = 8'hf7 == io_state_in_5 ? 8'hf5 : _GEN_2806; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2808 = 8'hf8 == io_state_in_5 ? 8'heb : _GEN_2807; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2809 = 8'hf9 == io_state_in_5 ? 8'he9 : _GEN_2808; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2810 = 8'hfa == io_state_in_5 ? 8'hef : _GEN_2809; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2811 = 8'hfb == io_state_in_5 ? 8'hed : _GEN_2810; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2812 = 8'hfc == io_state_in_5 ? 8'he3 : _GEN_2811; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2813 = 8'hfd == io_state_in_5 ? 8'he1 : _GEN_2812; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2814 = 8'hfe == io_state_in_5 ? 8'he7 : _GEN_2813; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _GEN_2815 = 8'hff == io_state_in_5 ? 8'he5 : _GEN_2814; // @[MixColumns.scala 131:{34,34}]
  wire [7:0] _tmp_state_5_T = io_state_in_4 ^ _GEN_2815; // @[MixColumns.scala 131:34]
  wire [7:0] _GEN_2817 = 8'h1 == io_state_in_6 ? 8'h3 : 8'h0; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2818 = 8'h2 == io_state_in_6 ? 8'h6 : _GEN_2817; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2819 = 8'h3 == io_state_in_6 ? 8'h5 : _GEN_2818; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2820 = 8'h4 == io_state_in_6 ? 8'hc : _GEN_2819; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2821 = 8'h5 == io_state_in_6 ? 8'hf : _GEN_2820; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2822 = 8'h6 == io_state_in_6 ? 8'ha : _GEN_2821; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2823 = 8'h7 == io_state_in_6 ? 8'h9 : _GEN_2822; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2824 = 8'h8 == io_state_in_6 ? 8'h18 : _GEN_2823; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2825 = 8'h9 == io_state_in_6 ? 8'h1b : _GEN_2824; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2826 = 8'ha == io_state_in_6 ? 8'h1e : _GEN_2825; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2827 = 8'hb == io_state_in_6 ? 8'h1d : _GEN_2826; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2828 = 8'hc == io_state_in_6 ? 8'h14 : _GEN_2827; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2829 = 8'hd == io_state_in_6 ? 8'h17 : _GEN_2828; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2830 = 8'he == io_state_in_6 ? 8'h12 : _GEN_2829; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2831 = 8'hf == io_state_in_6 ? 8'h11 : _GEN_2830; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2832 = 8'h10 == io_state_in_6 ? 8'h30 : _GEN_2831; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2833 = 8'h11 == io_state_in_6 ? 8'h33 : _GEN_2832; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2834 = 8'h12 == io_state_in_6 ? 8'h36 : _GEN_2833; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2835 = 8'h13 == io_state_in_6 ? 8'h35 : _GEN_2834; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2836 = 8'h14 == io_state_in_6 ? 8'h3c : _GEN_2835; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2837 = 8'h15 == io_state_in_6 ? 8'h3f : _GEN_2836; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2838 = 8'h16 == io_state_in_6 ? 8'h3a : _GEN_2837; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2839 = 8'h17 == io_state_in_6 ? 8'h39 : _GEN_2838; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2840 = 8'h18 == io_state_in_6 ? 8'h28 : _GEN_2839; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2841 = 8'h19 == io_state_in_6 ? 8'h2b : _GEN_2840; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2842 = 8'h1a == io_state_in_6 ? 8'h2e : _GEN_2841; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2843 = 8'h1b == io_state_in_6 ? 8'h2d : _GEN_2842; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2844 = 8'h1c == io_state_in_6 ? 8'h24 : _GEN_2843; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2845 = 8'h1d == io_state_in_6 ? 8'h27 : _GEN_2844; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2846 = 8'h1e == io_state_in_6 ? 8'h22 : _GEN_2845; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2847 = 8'h1f == io_state_in_6 ? 8'h21 : _GEN_2846; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2848 = 8'h20 == io_state_in_6 ? 8'h60 : _GEN_2847; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2849 = 8'h21 == io_state_in_6 ? 8'h63 : _GEN_2848; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2850 = 8'h22 == io_state_in_6 ? 8'h66 : _GEN_2849; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2851 = 8'h23 == io_state_in_6 ? 8'h65 : _GEN_2850; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2852 = 8'h24 == io_state_in_6 ? 8'h6c : _GEN_2851; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2853 = 8'h25 == io_state_in_6 ? 8'h6f : _GEN_2852; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2854 = 8'h26 == io_state_in_6 ? 8'h6a : _GEN_2853; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2855 = 8'h27 == io_state_in_6 ? 8'h69 : _GEN_2854; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2856 = 8'h28 == io_state_in_6 ? 8'h78 : _GEN_2855; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2857 = 8'h29 == io_state_in_6 ? 8'h7b : _GEN_2856; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2858 = 8'h2a == io_state_in_6 ? 8'h7e : _GEN_2857; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2859 = 8'h2b == io_state_in_6 ? 8'h7d : _GEN_2858; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2860 = 8'h2c == io_state_in_6 ? 8'h74 : _GEN_2859; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2861 = 8'h2d == io_state_in_6 ? 8'h77 : _GEN_2860; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2862 = 8'h2e == io_state_in_6 ? 8'h72 : _GEN_2861; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2863 = 8'h2f == io_state_in_6 ? 8'h71 : _GEN_2862; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2864 = 8'h30 == io_state_in_6 ? 8'h50 : _GEN_2863; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2865 = 8'h31 == io_state_in_6 ? 8'h53 : _GEN_2864; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2866 = 8'h32 == io_state_in_6 ? 8'h56 : _GEN_2865; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2867 = 8'h33 == io_state_in_6 ? 8'h55 : _GEN_2866; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2868 = 8'h34 == io_state_in_6 ? 8'h5c : _GEN_2867; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2869 = 8'h35 == io_state_in_6 ? 8'h5f : _GEN_2868; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2870 = 8'h36 == io_state_in_6 ? 8'h5a : _GEN_2869; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2871 = 8'h37 == io_state_in_6 ? 8'h59 : _GEN_2870; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2872 = 8'h38 == io_state_in_6 ? 8'h48 : _GEN_2871; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2873 = 8'h39 == io_state_in_6 ? 8'h4b : _GEN_2872; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2874 = 8'h3a == io_state_in_6 ? 8'h4e : _GEN_2873; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2875 = 8'h3b == io_state_in_6 ? 8'h4d : _GEN_2874; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2876 = 8'h3c == io_state_in_6 ? 8'h44 : _GEN_2875; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2877 = 8'h3d == io_state_in_6 ? 8'h47 : _GEN_2876; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2878 = 8'h3e == io_state_in_6 ? 8'h42 : _GEN_2877; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2879 = 8'h3f == io_state_in_6 ? 8'h41 : _GEN_2878; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2880 = 8'h40 == io_state_in_6 ? 8'hc0 : _GEN_2879; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2881 = 8'h41 == io_state_in_6 ? 8'hc3 : _GEN_2880; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2882 = 8'h42 == io_state_in_6 ? 8'hc6 : _GEN_2881; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2883 = 8'h43 == io_state_in_6 ? 8'hc5 : _GEN_2882; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2884 = 8'h44 == io_state_in_6 ? 8'hcc : _GEN_2883; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2885 = 8'h45 == io_state_in_6 ? 8'hcf : _GEN_2884; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2886 = 8'h46 == io_state_in_6 ? 8'hca : _GEN_2885; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2887 = 8'h47 == io_state_in_6 ? 8'hc9 : _GEN_2886; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2888 = 8'h48 == io_state_in_6 ? 8'hd8 : _GEN_2887; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2889 = 8'h49 == io_state_in_6 ? 8'hdb : _GEN_2888; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2890 = 8'h4a == io_state_in_6 ? 8'hde : _GEN_2889; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2891 = 8'h4b == io_state_in_6 ? 8'hdd : _GEN_2890; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2892 = 8'h4c == io_state_in_6 ? 8'hd4 : _GEN_2891; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2893 = 8'h4d == io_state_in_6 ? 8'hd7 : _GEN_2892; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2894 = 8'h4e == io_state_in_6 ? 8'hd2 : _GEN_2893; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2895 = 8'h4f == io_state_in_6 ? 8'hd1 : _GEN_2894; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2896 = 8'h50 == io_state_in_6 ? 8'hf0 : _GEN_2895; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2897 = 8'h51 == io_state_in_6 ? 8'hf3 : _GEN_2896; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2898 = 8'h52 == io_state_in_6 ? 8'hf6 : _GEN_2897; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2899 = 8'h53 == io_state_in_6 ? 8'hf5 : _GEN_2898; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2900 = 8'h54 == io_state_in_6 ? 8'hfc : _GEN_2899; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2901 = 8'h55 == io_state_in_6 ? 8'hff : _GEN_2900; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2902 = 8'h56 == io_state_in_6 ? 8'hfa : _GEN_2901; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2903 = 8'h57 == io_state_in_6 ? 8'hf9 : _GEN_2902; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2904 = 8'h58 == io_state_in_6 ? 8'he8 : _GEN_2903; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2905 = 8'h59 == io_state_in_6 ? 8'heb : _GEN_2904; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2906 = 8'h5a == io_state_in_6 ? 8'hee : _GEN_2905; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2907 = 8'h5b == io_state_in_6 ? 8'hed : _GEN_2906; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2908 = 8'h5c == io_state_in_6 ? 8'he4 : _GEN_2907; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2909 = 8'h5d == io_state_in_6 ? 8'he7 : _GEN_2908; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2910 = 8'h5e == io_state_in_6 ? 8'he2 : _GEN_2909; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2911 = 8'h5f == io_state_in_6 ? 8'he1 : _GEN_2910; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2912 = 8'h60 == io_state_in_6 ? 8'ha0 : _GEN_2911; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2913 = 8'h61 == io_state_in_6 ? 8'ha3 : _GEN_2912; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2914 = 8'h62 == io_state_in_6 ? 8'ha6 : _GEN_2913; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2915 = 8'h63 == io_state_in_6 ? 8'ha5 : _GEN_2914; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2916 = 8'h64 == io_state_in_6 ? 8'hac : _GEN_2915; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2917 = 8'h65 == io_state_in_6 ? 8'haf : _GEN_2916; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2918 = 8'h66 == io_state_in_6 ? 8'haa : _GEN_2917; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2919 = 8'h67 == io_state_in_6 ? 8'ha9 : _GEN_2918; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2920 = 8'h68 == io_state_in_6 ? 8'hb8 : _GEN_2919; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2921 = 8'h69 == io_state_in_6 ? 8'hbb : _GEN_2920; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2922 = 8'h6a == io_state_in_6 ? 8'hbe : _GEN_2921; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2923 = 8'h6b == io_state_in_6 ? 8'hbd : _GEN_2922; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2924 = 8'h6c == io_state_in_6 ? 8'hb4 : _GEN_2923; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2925 = 8'h6d == io_state_in_6 ? 8'hb7 : _GEN_2924; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2926 = 8'h6e == io_state_in_6 ? 8'hb2 : _GEN_2925; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2927 = 8'h6f == io_state_in_6 ? 8'hb1 : _GEN_2926; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2928 = 8'h70 == io_state_in_6 ? 8'h90 : _GEN_2927; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2929 = 8'h71 == io_state_in_6 ? 8'h93 : _GEN_2928; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2930 = 8'h72 == io_state_in_6 ? 8'h96 : _GEN_2929; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2931 = 8'h73 == io_state_in_6 ? 8'h95 : _GEN_2930; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2932 = 8'h74 == io_state_in_6 ? 8'h9c : _GEN_2931; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2933 = 8'h75 == io_state_in_6 ? 8'h9f : _GEN_2932; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2934 = 8'h76 == io_state_in_6 ? 8'h9a : _GEN_2933; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2935 = 8'h77 == io_state_in_6 ? 8'h99 : _GEN_2934; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2936 = 8'h78 == io_state_in_6 ? 8'h88 : _GEN_2935; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2937 = 8'h79 == io_state_in_6 ? 8'h8b : _GEN_2936; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2938 = 8'h7a == io_state_in_6 ? 8'h8e : _GEN_2937; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2939 = 8'h7b == io_state_in_6 ? 8'h8d : _GEN_2938; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2940 = 8'h7c == io_state_in_6 ? 8'h84 : _GEN_2939; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2941 = 8'h7d == io_state_in_6 ? 8'h87 : _GEN_2940; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2942 = 8'h7e == io_state_in_6 ? 8'h82 : _GEN_2941; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2943 = 8'h7f == io_state_in_6 ? 8'h81 : _GEN_2942; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2944 = 8'h80 == io_state_in_6 ? 8'h9b : _GEN_2943; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2945 = 8'h81 == io_state_in_6 ? 8'h98 : _GEN_2944; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2946 = 8'h82 == io_state_in_6 ? 8'h9d : _GEN_2945; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2947 = 8'h83 == io_state_in_6 ? 8'h9e : _GEN_2946; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2948 = 8'h84 == io_state_in_6 ? 8'h97 : _GEN_2947; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2949 = 8'h85 == io_state_in_6 ? 8'h94 : _GEN_2948; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2950 = 8'h86 == io_state_in_6 ? 8'h91 : _GEN_2949; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2951 = 8'h87 == io_state_in_6 ? 8'h92 : _GEN_2950; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2952 = 8'h88 == io_state_in_6 ? 8'h83 : _GEN_2951; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2953 = 8'h89 == io_state_in_6 ? 8'h80 : _GEN_2952; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2954 = 8'h8a == io_state_in_6 ? 8'h85 : _GEN_2953; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2955 = 8'h8b == io_state_in_6 ? 8'h86 : _GEN_2954; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2956 = 8'h8c == io_state_in_6 ? 8'h8f : _GEN_2955; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2957 = 8'h8d == io_state_in_6 ? 8'h8c : _GEN_2956; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2958 = 8'h8e == io_state_in_6 ? 8'h89 : _GEN_2957; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2959 = 8'h8f == io_state_in_6 ? 8'h8a : _GEN_2958; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2960 = 8'h90 == io_state_in_6 ? 8'hab : _GEN_2959; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2961 = 8'h91 == io_state_in_6 ? 8'ha8 : _GEN_2960; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2962 = 8'h92 == io_state_in_6 ? 8'had : _GEN_2961; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2963 = 8'h93 == io_state_in_6 ? 8'hae : _GEN_2962; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2964 = 8'h94 == io_state_in_6 ? 8'ha7 : _GEN_2963; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2965 = 8'h95 == io_state_in_6 ? 8'ha4 : _GEN_2964; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2966 = 8'h96 == io_state_in_6 ? 8'ha1 : _GEN_2965; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2967 = 8'h97 == io_state_in_6 ? 8'ha2 : _GEN_2966; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2968 = 8'h98 == io_state_in_6 ? 8'hb3 : _GEN_2967; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2969 = 8'h99 == io_state_in_6 ? 8'hb0 : _GEN_2968; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2970 = 8'h9a == io_state_in_6 ? 8'hb5 : _GEN_2969; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2971 = 8'h9b == io_state_in_6 ? 8'hb6 : _GEN_2970; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2972 = 8'h9c == io_state_in_6 ? 8'hbf : _GEN_2971; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2973 = 8'h9d == io_state_in_6 ? 8'hbc : _GEN_2972; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2974 = 8'h9e == io_state_in_6 ? 8'hb9 : _GEN_2973; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2975 = 8'h9f == io_state_in_6 ? 8'hba : _GEN_2974; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2976 = 8'ha0 == io_state_in_6 ? 8'hfb : _GEN_2975; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2977 = 8'ha1 == io_state_in_6 ? 8'hf8 : _GEN_2976; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2978 = 8'ha2 == io_state_in_6 ? 8'hfd : _GEN_2977; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2979 = 8'ha3 == io_state_in_6 ? 8'hfe : _GEN_2978; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2980 = 8'ha4 == io_state_in_6 ? 8'hf7 : _GEN_2979; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2981 = 8'ha5 == io_state_in_6 ? 8'hf4 : _GEN_2980; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2982 = 8'ha6 == io_state_in_6 ? 8'hf1 : _GEN_2981; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2983 = 8'ha7 == io_state_in_6 ? 8'hf2 : _GEN_2982; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2984 = 8'ha8 == io_state_in_6 ? 8'he3 : _GEN_2983; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2985 = 8'ha9 == io_state_in_6 ? 8'he0 : _GEN_2984; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2986 = 8'haa == io_state_in_6 ? 8'he5 : _GEN_2985; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2987 = 8'hab == io_state_in_6 ? 8'he6 : _GEN_2986; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2988 = 8'hac == io_state_in_6 ? 8'hef : _GEN_2987; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2989 = 8'had == io_state_in_6 ? 8'hec : _GEN_2988; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2990 = 8'hae == io_state_in_6 ? 8'he9 : _GEN_2989; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2991 = 8'haf == io_state_in_6 ? 8'hea : _GEN_2990; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2992 = 8'hb0 == io_state_in_6 ? 8'hcb : _GEN_2991; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2993 = 8'hb1 == io_state_in_6 ? 8'hc8 : _GEN_2992; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2994 = 8'hb2 == io_state_in_6 ? 8'hcd : _GEN_2993; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2995 = 8'hb3 == io_state_in_6 ? 8'hce : _GEN_2994; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2996 = 8'hb4 == io_state_in_6 ? 8'hc7 : _GEN_2995; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2997 = 8'hb5 == io_state_in_6 ? 8'hc4 : _GEN_2996; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2998 = 8'hb6 == io_state_in_6 ? 8'hc1 : _GEN_2997; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_2999 = 8'hb7 == io_state_in_6 ? 8'hc2 : _GEN_2998; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3000 = 8'hb8 == io_state_in_6 ? 8'hd3 : _GEN_2999; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3001 = 8'hb9 == io_state_in_6 ? 8'hd0 : _GEN_3000; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3002 = 8'hba == io_state_in_6 ? 8'hd5 : _GEN_3001; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3003 = 8'hbb == io_state_in_6 ? 8'hd6 : _GEN_3002; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3004 = 8'hbc == io_state_in_6 ? 8'hdf : _GEN_3003; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3005 = 8'hbd == io_state_in_6 ? 8'hdc : _GEN_3004; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3006 = 8'hbe == io_state_in_6 ? 8'hd9 : _GEN_3005; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3007 = 8'hbf == io_state_in_6 ? 8'hda : _GEN_3006; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3008 = 8'hc0 == io_state_in_6 ? 8'h5b : _GEN_3007; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3009 = 8'hc1 == io_state_in_6 ? 8'h58 : _GEN_3008; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3010 = 8'hc2 == io_state_in_6 ? 8'h5d : _GEN_3009; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3011 = 8'hc3 == io_state_in_6 ? 8'h5e : _GEN_3010; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3012 = 8'hc4 == io_state_in_6 ? 8'h57 : _GEN_3011; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3013 = 8'hc5 == io_state_in_6 ? 8'h54 : _GEN_3012; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3014 = 8'hc6 == io_state_in_6 ? 8'h51 : _GEN_3013; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3015 = 8'hc7 == io_state_in_6 ? 8'h52 : _GEN_3014; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3016 = 8'hc8 == io_state_in_6 ? 8'h43 : _GEN_3015; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3017 = 8'hc9 == io_state_in_6 ? 8'h40 : _GEN_3016; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3018 = 8'hca == io_state_in_6 ? 8'h45 : _GEN_3017; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3019 = 8'hcb == io_state_in_6 ? 8'h46 : _GEN_3018; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3020 = 8'hcc == io_state_in_6 ? 8'h4f : _GEN_3019; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3021 = 8'hcd == io_state_in_6 ? 8'h4c : _GEN_3020; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3022 = 8'hce == io_state_in_6 ? 8'h49 : _GEN_3021; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3023 = 8'hcf == io_state_in_6 ? 8'h4a : _GEN_3022; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3024 = 8'hd0 == io_state_in_6 ? 8'h6b : _GEN_3023; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3025 = 8'hd1 == io_state_in_6 ? 8'h68 : _GEN_3024; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3026 = 8'hd2 == io_state_in_6 ? 8'h6d : _GEN_3025; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3027 = 8'hd3 == io_state_in_6 ? 8'h6e : _GEN_3026; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3028 = 8'hd4 == io_state_in_6 ? 8'h67 : _GEN_3027; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3029 = 8'hd5 == io_state_in_6 ? 8'h64 : _GEN_3028; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3030 = 8'hd6 == io_state_in_6 ? 8'h61 : _GEN_3029; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3031 = 8'hd7 == io_state_in_6 ? 8'h62 : _GEN_3030; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3032 = 8'hd8 == io_state_in_6 ? 8'h73 : _GEN_3031; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3033 = 8'hd9 == io_state_in_6 ? 8'h70 : _GEN_3032; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3034 = 8'hda == io_state_in_6 ? 8'h75 : _GEN_3033; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3035 = 8'hdb == io_state_in_6 ? 8'h76 : _GEN_3034; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3036 = 8'hdc == io_state_in_6 ? 8'h7f : _GEN_3035; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3037 = 8'hdd == io_state_in_6 ? 8'h7c : _GEN_3036; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3038 = 8'hde == io_state_in_6 ? 8'h79 : _GEN_3037; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3039 = 8'hdf == io_state_in_6 ? 8'h7a : _GEN_3038; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3040 = 8'he0 == io_state_in_6 ? 8'h3b : _GEN_3039; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3041 = 8'he1 == io_state_in_6 ? 8'h38 : _GEN_3040; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3042 = 8'he2 == io_state_in_6 ? 8'h3d : _GEN_3041; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3043 = 8'he3 == io_state_in_6 ? 8'h3e : _GEN_3042; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3044 = 8'he4 == io_state_in_6 ? 8'h37 : _GEN_3043; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3045 = 8'he5 == io_state_in_6 ? 8'h34 : _GEN_3044; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3046 = 8'he6 == io_state_in_6 ? 8'h31 : _GEN_3045; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3047 = 8'he7 == io_state_in_6 ? 8'h32 : _GEN_3046; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3048 = 8'he8 == io_state_in_6 ? 8'h23 : _GEN_3047; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3049 = 8'he9 == io_state_in_6 ? 8'h20 : _GEN_3048; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3050 = 8'hea == io_state_in_6 ? 8'h25 : _GEN_3049; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3051 = 8'heb == io_state_in_6 ? 8'h26 : _GEN_3050; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3052 = 8'hec == io_state_in_6 ? 8'h2f : _GEN_3051; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3053 = 8'hed == io_state_in_6 ? 8'h2c : _GEN_3052; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3054 = 8'hee == io_state_in_6 ? 8'h29 : _GEN_3053; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3055 = 8'hef == io_state_in_6 ? 8'h2a : _GEN_3054; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3056 = 8'hf0 == io_state_in_6 ? 8'hb : _GEN_3055; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3057 = 8'hf1 == io_state_in_6 ? 8'h8 : _GEN_3056; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3058 = 8'hf2 == io_state_in_6 ? 8'hd : _GEN_3057; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3059 = 8'hf3 == io_state_in_6 ? 8'he : _GEN_3058; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3060 = 8'hf4 == io_state_in_6 ? 8'h7 : _GEN_3059; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3061 = 8'hf5 == io_state_in_6 ? 8'h4 : _GEN_3060; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3062 = 8'hf6 == io_state_in_6 ? 8'h1 : _GEN_3061; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3063 = 8'hf7 == io_state_in_6 ? 8'h2 : _GEN_3062; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3064 = 8'hf8 == io_state_in_6 ? 8'h13 : _GEN_3063; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3065 = 8'hf9 == io_state_in_6 ? 8'h10 : _GEN_3064; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3066 = 8'hfa == io_state_in_6 ? 8'h15 : _GEN_3065; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3067 = 8'hfb == io_state_in_6 ? 8'h16 : _GEN_3066; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3068 = 8'hfc == io_state_in_6 ? 8'h1f : _GEN_3067; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3069 = 8'hfd == io_state_in_6 ? 8'h1c : _GEN_3068; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3070 = 8'hfe == io_state_in_6 ? 8'h19 : _GEN_3069; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _GEN_3071 = 8'hff == io_state_in_6 ? 8'h1a : _GEN_3070; // @[MixColumns.scala 131:{58,58}]
  wire [7:0] _tmp_state_5_T_1 = _tmp_state_5_T ^ _GEN_3071; // @[MixColumns.scala 131:58]
  wire [7:0] _tmp_state_6_T = io_state_in_4 ^ io_state_in_5; // @[MixColumns.scala 132:34]
  wire [7:0] _GEN_3073 = 8'h1 == io_state_in_6 ? 8'h2 : 8'h0; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3074 = 8'h2 == io_state_in_6 ? 8'h4 : _GEN_3073; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3075 = 8'h3 == io_state_in_6 ? 8'h6 : _GEN_3074; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3076 = 8'h4 == io_state_in_6 ? 8'h8 : _GEN_3075; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3077 = 8'h5 == io_state_in_6 ? 8'ha : _GEN_3076; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3078 = 8'h6 == io_state_in_6 ? 8'hc : _GEN_3077; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3079 = 8'h7 == io_state_in_6 ? 8'he : _GEN_3078; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3080 = 8'h8 == io_state_in_6 ? 8'h10 : _GEN_3079; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3081 = 8'h9 == io_state_in_6 ? 8'h12 : _GEN_3080; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3082 = 8'ha == io_state_in_6 ? 8'h14 : _GEN_3081; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3083 = 8'hb == io_state_in_6 ? 8'h16 : _GEN_3082; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3084 = 8'hc == io_state_in_6 ? 8'h18 : _GEN_3083; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3085 = 8'hd == io_state_in_6 ? 8'h1a : _GEN_3084; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3086 = 8'he == io_state_in_6 ? 8'h1c : _GEN_3085; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3087 = 8'hf == io_state_in_6 ? 8'h1e : _GEN_3086; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3088 = 8'h10 == io_state_in_6 ? 8'h20 : _GEN_3087; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3089 = 8'h11 == io_state_in_6 ? 8'h22 : _GEN_3088; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3090 = 8'h12 == io_state_in_6 ? 8'h24 : _GEN_3089; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3091 = 8'h13 == io_state_in_6 ? 8'h26 : _GEN_3090; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3092 = 8'h14 == io_state_in_6 ? 8'h28 : _GEN_3091; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3093 = 8'h15 == io_state_in_6 ? 8'h2a : _GEN_3092; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3094 = 8'h16 == io_state_in_6 ? 8'h2c : _GEN_3093; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3095 = 8'h17 == io_state_in_6 ? 8'h2e : _GEN_3094; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3096 = 8'h18 == io_state_in_6 ? 8'h30 : _GEN_3095; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3097 = 8'h19 == io_state_in_6 ? 8'h32 : _GEN_3096; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3098 = 8'h1a == io_state_in_6 ? 8'h34 : _GEN_3097; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3099 = 8'h1b == io_state_in_6 ? 8'h36 : _GEN_3098; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3100 = 8'h1c == io_state_in_6 ? 8'h38 : _GEN_3099; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3101 = 8'h1d == io_state_in_6 ? 8'h3a : _GEN_3100; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3102 = 8'h1e == io_state_in_6 ? 8'h3c : _GEN_3101; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3103 = 8'h1f == io_state_in_6 ? 8'h3e : _GEN_3102; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3104 = 8'h20 == io_state_in_6 ? 8'h40 : _GEN_3103; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3105 = 8'h21 == io_state_in_6 ? 8'h42 : _GEN_3104; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3106 = 8'h22 == io_state_in_6 ? 8'h44 : _GEN_3105; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3107 = 8'h23 == io_state_in_6 ? 8'h46 : _GEN_3106; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3108 = 8'h24 == io_state_in_6 ? 8'h48 : _GEN_3107; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3109 = 8'h25 == io_state_in_6 ? 8'h4a : _GEN_3108; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3110 = 8'h26 == io_state_in_6 ? 8'h4c : _GEN_3109; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3111 = 8'h27 == io_state_in_6 ? 8'h4e : _GEN_3110; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3112 = 8'h28 == io_state_in_6 ? 8'h50 : _GEN_3111; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3113 = 8'h29 == io_state_in_6 ? 8'h52 : _GEN_3112; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3114 = 8'h2a == io_state_in_6 ? 8'h54 : _GEN_3113; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3115 = 8'h2b == io_state_in_6 ? 8'h56 : _GEN_3114; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3116 = 8'h2c == io_state_in_6 ? 8'h58 : _GEN_3115; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3117 = 8'h2d == io_state_in_6 ? 8'h5a : _GEN_3116; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3118 = 8'h2e == io_state_in_6 ? 8'h5c : _GEN_3117; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3119 = 8'h2f == io_state_in_6 ? 8'h5e : _GEN_3118; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3120 = 8'h30 == io_state_in_6 ? 8'h60 : _GEN_3119; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3121 = 8'h31 == io_state_in_6 ? 8'h62 : _GEN_3120; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3122 = 8'h32 == io_state_in_6 ? 8'h64 : _GEN_3121; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3123 = 8'h33 == io_state_in_6 ? 8'h66 : _GEN_3122; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3124 = 8'h34 == io_state_in_6 ? 8'h68 : _GEN_3123; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3125 = 8'h35 == io_state_in_6 ? 8'h6a : _GEN_3124; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3126 = 8'h36 == io_state_in_6 ? 8'h6c : _GEN_3125; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3127 = 8'h37 == io_state_in_6 ? 8'h6e : _GEN_3126; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3128 = 8'h38 == io_state_in_6 ? 8'h70 : _GEN_3127; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3129 = 8'h39 == io_state_in_6 ? 8'h72 : _GEN_3128; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3130 = 8'h3a == io_state_in_6 ? 8'h74 : _GEN_3129; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3131 = 8'h3b == io_state_in_6 ? 8'h76 : _GEN_3130; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3132 = 8'h3c == io_state_in_6 ? 8'h78 : _GEN_3131; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3133 = 8'h3d == io_state_in_6 ? 8'h7a : _GEN_3132; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3134 = 8'h3e == io_state_in_6 ? 8'h7c : _GEN_3133; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3135 = 8'h3f == io_state_in_6 ? 8'h7e : _GEN_3134; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3136 = 8'h40 == io_state_in_6 ? 8'h80 : _GEN_3135; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3137 = 8'h41 == io_state_in_6 ? 8'h82 : _GEN_3136; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3138 = 8'h42 == io_state_in_6 ? 8'h84 : _GEN_3137; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3139 = 8'h43 == io_state_in_6 ? 8'h86 : _GEN_3138; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3140 = 8'h44 == io_state_in_6 ? 8'h88 : _GEN_3139; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3141 = 8'h45 == io_state_in_6 ? 8'h8a : _GEN_3140; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3142 = 8'h46 == io_state_in_6 ? 8'h8c : _GEN_3141; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3143 = 8'h47 == io_state_in_6 ? 8'h8e : _GEN_3142; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3144 = 8'h48 == io_state_in_6 ? 8'h90 : _GEN_3143; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3145 = 8'h49 == io_state_in_6 ? 8'h92 : _GEN_3144; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3146 = 8'h4a == io_state_in_6 ? 8'h94 : _GEN_3145; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3147 = 8'h4b == io_state_in_6 ? 8'h96 : _GEN_3146; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3148 = 8'h4c == io_state_in_6 ? 8'h98 : _GEN_3147; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3149 = 8'h4d == io_state_in_6 ? 8'h9a : _GEN_3148; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3150 = 8'h4e == io_state_in_6 ? 8'h9c : _GEN_3149; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3151 = 8'h4f == io_state_in_6 ? 8'h9e : _GEN_3150; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3152 = 8'h50 == io_state_in_6 ? 8'ha0 : _GEN_3151; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3153 = 8'h51 == io_state_in_6 ? 8'ha2 : _GEN_3152; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3154 = 8'h52 == io_state_in_6 ? 8'ha4 : _GEN_3153; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3155 = 8'h53 == io_state_in_6 ? 8'ha6 : _GEN_3154; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3156 = 8'h54 == io_state_in_6 ? 8'ha8 : _GEN_3155; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3157 = 8'h55 == io_state_in_6 ? 8'haa : _GEN_3156; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3158 = 8'h56 == io_state_in_6 ? 8'hac : _GEN_3157; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3159 = 8'h57 == io_state_in_6 ? 8'hae : _GEN_3158; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3160 = 8'h58 == io_state_in_6 ? 8'hb0 : _GEN_3159; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3161 = 8'h59 == io_state_in_6 ? 8'hb2 : _GEN_3160; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3162 = 8'h5a == io_state_in_6 ? 8'hb4 : _GEN_3161; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3163 = 8'h5b == io_state_in_6 ? 8'hb6 : _GEN_3162; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3164 = 8'h5c == io_state_in_6 ? 8'hb8 : _GEN_3163; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3165 = 8'h5d == io_state_in_6 ? 8'hba : _GEN_3164; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3166 = 8'h5e == io_state_in_6 ? 8'hbc : _GEN_3165; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3167 = 8'h5f == io_state_in_6 ? 8'hbe : _GEN_3166; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3168 = 8'h60 == io_state_in_6 ? 8'hc0 : _GEN_3167; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3169 = 8'h61 == io_state_in_6 ? 8'hc2 : _GEN_3168; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3170 = 8'h62 == io_state_in_6 ? 8'hc4 : _GEN_3169; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3171 = 8'h63 == io_state_in_6 ? 8'hc6 : _GEN_3170; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3172 = 8'h64 == io_state_in_6 ? 8'hc8 : _GEN_3171; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3173 = 8'h65 == io_state_in_6 ? 8'hca : _GEN_3172; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3174 = 8'h66 == io_state_in_6 ? 8'hcc : _GEN_3173; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3175 = 8'h67 == io_state_in_6 ? 8'hce : _GEN_3174; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3176 = 8'h68 == io_state_in_6 ? 8'hd0 : _GEN_3175; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3177 = 8'h69 == io_state_in_6 ? 8'hd2 : _GEN_3176; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3178 = 8'h6a == io_state_in_6 ? 8'hd4 : _GEN_3177; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3179 = 8'h6b == io_state_in_6 ? 8'hd6 : _GEN_3178; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3180 = 8'h6c == io_state_in_6 ? 8'hd8 : _GEN_3179; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3181 = 8'h6d == io_state_in_6 ? 8'hda : _GEN_3180; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3182 = 8'h6e == io_state_in_6 ? 8'hdc : _GEN_3181; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3183 = 8'h6f == io_state_in_6 ? 8'hde : _GEN_3182; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3184 = 8'h70 == io_state_in_6 ? 8'he0 : _GEN_3183; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3185 = 8'h71 == io_state_in_6 ? 8'he2 : _GEN_3184; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3186 = 8'h72 == io_state_in_6 ? 8'he4 : _GEN_3185; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3187 = 8'h73 == io_state_in_6 ? 8'he6 : _GEN_3186; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3188 = 8'h74 == io_state_in_6 ? 8'he8 : _GEN_3187; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3189 = 8'h75 == io_state_in_6 ? 8'hea : _GEN_3188; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3190 = 8'h76 == io_state_in_6 ? 8'hec : _GEN_3189; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3191 = 8'h77 == io_state_in_6 ? 8'hee : _GEN_3190; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3192 = 8'h78 == io_state_in_6 ? 8'hf0 : _GEN_3191; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3193 = 8'h79 == io_state_in_6 ? 8'hf2 : _GEN_3192; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3194 = 8'h7a == io_state_in_6 ? 8'hf4 : _GEN_3193; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3195 = 8'h7b == io_state_in_6 ? 8'hf6 : _GEN_3194; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3196 = 8'h7c == io_state_in_6 ? 8'hf8 : _GEN_3195; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3197 = 8'h7d == io_state_in_6 ? 8'hfa : _GEN_3196; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3198 = 8'h7e == io_state_in_6 ? 8'hfc : _GEN_3197; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3199 = 8'h7f == io_state_in_6 ? 8'hfe : _GEN_3198; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3200 = 8'h80 == io_state_in_6 ? 8'h1b : _GEN_3199; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3201 = 8'h81 == io_state_in_6 ? 8'h19 : _GEN_3200; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3202 = 8'h82 == io_state_in_6 ? 8'h1f : _GEN_3201; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3203 = 8'h83 == io_state_in_6 ? 8'h1d : _GEN_3202; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3204 = 8'h84 == io_state_in_6 ? 8'h13 : _GEN_3203; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3205 = 8'h85 == io_state_in_6 ? 8'h11 : _GEN_3204; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3206 = 8'h86 == io_state_in_6 ? 8'h17 : _GEN_3205; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3207 = 8'h87 == io_state_in_6 ? 8'h15 : _GEN_3206; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3208 = 8'h88 == io_state_in_6 ? 8'hb : _GEN_3207; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3209 = 8'h89 == io_state_in_6 ? 8'h9 : _GEN_3208; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3210 = 8'h8a == io_state_in_6 ? 8'hf : _GEN_3209; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3211 = 8'h8b == io_state_in_6 ? 8'hd : _GEN_3210; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3212 = 8'h8c == io_state_in_6 ? 8'h3 : _GEN_3211; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3213 = 8'h8d == io_state_in_6 ? 8'h1 : _GEN_3212; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3214 = 8'h8e == io_state_in_6 ? 8'h7 : _GEN_3213; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3215 = 8'h8f == io_state_in_6 ? 8'h5 : _GEN_3214; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3216 = 8'h90 == io_state_in_6 ? 8'h3b : _GEN_3215; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3217 = 8'h91 == io_state_in_6 ? 8'h39 : _GEN_3216; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3218 = 8'h92 == io_state_in_6 ? 8'h3f : _GEN_3217; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3219 = 8'h93 == io_state_in_6 ? 8'h3d : _GEN_3218; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3220 = 8'h94 == io_state_in_6 ? 8'h33 : _GEN_3219; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3221 = 8'h95 == io_state_in_6 ? 8'h31 : _GEN_3220; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3222 = 8'h96 == io_state_in_6 ? 8'h37 : _GEN_3221; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3223 = 8'h97 == io_state_in_6 ? 8'h35 : _GEN_3222; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3224 = 8'h98 == io_state_in_6 ? 8'h2b : _GEN_3223; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3225 = 8'h99 == io_state_in_6 ? 8'h29 : _GEN_3224; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3226 = 8'h9a == io_state_in_6 ? 8'h2f : _GEN_3225; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3227 = 8'h9b == io_state_in_6 ? 8'h2d : _GEN_3226; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3228 = 8'h9c == io_state_in_6 ? 8'h23 : _GEN_3227; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3229 = 8'h9d == io_state_in_6 ? 8'h21 : _GEN_3228; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3230 = 8'h9e == io_state_in_6 ? 8'h27 : _GEN_3229; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3231 = 8'h9f == io_state_in_6 ? 8'h25 : _GEN_3230; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3232 = 8'ha0 == io_state_in_6 ? 8'h5b : _GEN_3231; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3233 = 8'ha1 == io_state_in_6 ? 8'h59 : _GEN_3232; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3234 = 8'ha2 == io_state_in_6 ? 8'h5f : _GEN_3233; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3235 = 8'ha3 == io_state_in_6 ? 8'h5d : _GEN_3234; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3236 = 8'ha4 == io_state_in_6 ? 8'h53 : _GEN_3235; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3237 = 8'ha5 == io_state_in_6 ? 8'h51 : _GEN_3236; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3238 = 8'ha6 == io_state_in_6 ? 8'h57 : _GEN_3237; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3239 = 8'ha7 == io_state_in_6 ? 8'h55 : _GEN_3238; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3240 = 8'ha8 == io_state_in_6 ? 8'h4b : _GEN_3239; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3241 = 8'ha9 == io_state_in_6 ? 8'h49 : _GEN_3240; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3242 = 8'haa == io_state_in_6 ? 8'h4f : _GEN_3241; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3243 = 8'hab == io_state_in_6 ? 8'h4d : _GEN_3242; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3244 = 8'hac == io_state_in_6 ? 8'h43 : _GEN_3243; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3245 = 8'had == io_state_in_6 ? 8'h41 : _GEN_3244; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3246 = 8'hae == io_state_in_6 ? 8'h47 : _GEN_3245; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3247 = 8'haf == io_state_in_6 ? 8'h45 : _GEN_3246; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3248 = 8'hb0 == io_state_in_6 ? 8'h7b : _GEN_3247; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3249 = 8'hb1 == io_state_in_6 ? 8'h79 : _GEN_3248; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3250 = 8'hb2 == io_state_in_6 ? 8'h7f : _GEN_3249; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3251 = 8'hb3 == io_state_in_6 ? 8'h7d : _GEN_3250; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3252 = 8'hb4 == io_state_in_6 ? 8'h73 : _GEN_3251; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3253 = 8'hb5 == io_state_in_6 ? 8'h71 : _GEN_3252; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3254 = 8'hb6 == io_state_in_6 ? 8'h77 : _GEN_3253; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3255 = 8'hb7 == io_state_in_6 ? 8'h75 : _GEN_3254; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3256 = 8'hb8 == io_state_in_6 ? 8'h6b : _GEN_3255; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3257 = 8'hb9 == io_state_in_6 ? 8'h69 : _GEN_3256; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3258 = 8'hba == io_state_in_6 ? 8'h6f : _GEN_3257; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3259 = 8'hbb == io_state_in_6 ? 8'h6d : _GEN_3258; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3260 = 8'hbc == io_state_in_6 ? 8'h63 : _GEN_3259; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3261 = 8'hbd == io_state_in_6 ? 8'h61 : _GEN_3260; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3262 = 8'hbe == io_state_in_6 ? 8'h67 : _GEN_3261; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3263 = 8'hbf == io_state_in_6 ? 8'h65 : _GEN_3262; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3264 = 8'hc0 == io_state_in_6 ? 8'h9b : _GEN_3263; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3265 = 8'hc1 == io_state_in_6 ? 8'h99 : _GEN_3264; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3266 = 8'hc2 == io_state_in_6 ? 8'h9f : _GEN_3265; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3267 = 8'hc3 == io_state_in_6 ? 8'h9d : _GEN_3266; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3268 = 8'hc4 == io_state_in_6 ? 8'h93 : _GEN_3267; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3269 = 8'hc5 == io_state_in_6 ? 8'h91 : _GEN_3268; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3270 = 8'hc6 == io_state_in_6 ? 8'h97 : _GEN_3269; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3271 = 8'hc7 == io_state_in_6 ? 8'h95 : _GEN_3270; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3272 = 8'hc8 == io_state_in_6 ? 8'h8b : _GEN_3271; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3273 = 8'hc9 == io_state_in_6 ? 8'h89 : _GEN_3272; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3274 = 8'hca == io_state_in_6 ? 8'h8f : _GEN_3273; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3275 = 8'hcb == io_state_in_6 ? 8'h8d : _GEN_3274; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3276 = 8'hcc == io_state_in_6 ? 8'h83 : _GEN_3275; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3277 = 8'hcd == io_state_in_6 ? 8'h81 : _GEN_3276; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3278 = 8'hce == io_state_in_6 ? 8'h87 : _GEN_3277; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3279 = 8'hcf == io_state_in_6 ? 8'h85 : _GEN_3278; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3280 = 8'hd0 == io_state_in_6 ? 8'hbb : _GEN_3279; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3281 = 8'hd1 == io_state_in_6 ? 8'hb9 : _GEN_3280; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3282 = 8'hd2 == io_state_in_6 ? 8'hbf : _GEN_3281; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3283 = 8'hd3 == io_state_in_6 ? 8'hbd : _GEN_3282; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3284 = 8'hd4 == io_state_in_6 ? 8'hb3 : _GEN_3283; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3285 = 8'hd5 == io_state_in_6 ? 8'hb1 : _GEN_3284; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3286 = 8'hd6 == io_state_in_6 ? 8'hb7 : _GEN_3285; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3287 = 8'hd7 == io_state_in_6 ? 8'hb5 : _GEN_3286; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3288 = 8'hd8 == io_state_in_6 ? 8'hab : _GEN_3287; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3289 = 8'hd9 == io_state_in_6 ? 8'ha9 : _GEN_3288; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3290 = 8'hda == io_state_in_6 ? 8'haf : _GEN_3289; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3291 = 8'hdb == io_state_in_6 ? 8'had : _GEN_3290; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3292 = 8'hdc == io_state_in_6 ? 8'ha3 : _GEN_3291; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3293 = 8'hdd == io_state_in_6 ? 8'ha1 : _GEN_3292; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3294 = 8'hde == io_state_in_6 ? 8'ha7 : _GEN_3293; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3295 = 8'hdf == io_state_in_6 ? 8'ha5 : _GEN_3294; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3296 = 8'he0 == io_state_in_6 ? 8'hdb : _GEN_3295; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3297 = 8'he1 == io_state_in_6 ? 8'hd9 : _GEN_3296; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3298 = 8'he2 == io_state_in_6 ? 8'hdf : _GEN_3297; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3299 = 8'he3 == io_state_in_6 ? 8'hdd : _GEN_3298; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3300 = 8'he4 == io_state_in_6 ? 8'hd3 : _GEN_3299; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3301 = 8'he5 == io_state_in_6 ? 8'hd1 : _GEN_3300; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3302 = 8'he6 == io_state_in_6 ? 8'hd7 : _GEN_3301; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3303 = 8'he7 == io_state_in_6 ? 8'hd5 : _GEN_3302; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3304 = 8'he8 == io_state_in_6 ? 8'hcb : _GEN_3303; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3305 = 8'he9 == io_state_in_6 ? 8'hc9 : _GEN_3304; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3306 = 8'hea == io_state_in_6 ? 8'hcf : _GEN_3305; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3307 = 8'heb == io_state_in_6 ? 8'hcd : _GEN_3306; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3308 = 8'hec == io_state_in_6 ? 8'hc3 : _GEN_3307; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3309 = 8'hed == io_state_in_6 ? 8'hc1 : _GEN_3308; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3310 = 8'hee == io_state_in_6 ? 8'hc7 : _GEN_3309; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3311 = 8'hef == io_state_in_6 ? 8'hc5 : _GEN_3310; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3312 = 8'hf0 == io_state_in_6 ? 8'hfb : _GEN_3311; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3313 = 8'hf1 == io_state_in_6 ? 8'hf9 : _GEN_3312; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3314 = 8'hf2 == io_state_in_6 ? 8'hff : _GEN_3313; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3315 = 8'hf3 == io_state_in_6 ? 8'hfd : _GEN_3314; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3316 = 8'hf4 == io_state_in_6 ? 8'hf3 : _GEN_3315; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3317 = 8'hf5 == io_state_in_6 ? 8'hf1 : _GEN_3316; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3318 = 8'hf6 == io_state_in_6 ? 8'hf7 : _GEN_3317; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3319 = 8'hf7 == io_state_in_6 ? 8'hf5 : _GEN_3318; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3320 = 8'hf8 == io_state_in_6 ? 8'heb : _GEN_3319; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3321 = 8'hf9 == io_state_in_6 ? 8'he9 : _GEN_3320; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3322 = 8'hfa == io_state_in_6 ? 8'hef : _GEN_3321; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3323 = 8'hfb == io_state_in_6 ? 8'hed : _GEN_3322; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3324 = 8'hfc == io_state_in_6 ? 8'he3 : _GEN_3323; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3325 = 8'hfd == io_state_in_6 ? 8'he1 : _GEN_3324; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3326 = 8'hfe == io_state_in_6 ? 8'he7 : _GEN_3325; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _GEN_3327 = 8'hff == io_state_in_6 ? 8'he5 : _GEN_3326; // @[MixColumns.scala 132:{51,51}]
  wire [7:0] _tmp_state_6_T_1 = _tmp_state_6_T ^ _GEN_3327; // @[MixColumns.scala 132:51]
  wire [7:0] _GEN_3329 = 8'h1 == io_state_in_7 ? 8'h3 : 8'h0; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3330 = 8'h2 == io_state_in_7 ? 8'h6 : _GEN_3329; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3331 = 8'h3 == io_state_in_7 ? 8'h5 : _GEN_3330; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3332 = 8'h4 == io_state_in_7 ? 8'hc : _GEN_3331; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3333 = 8'h5 == io_state_in_7 ? 8'hf : _GEN_3332; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3334 = 8'h6 == io_state_in_7 ? 8'ha : _GEN_3333; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3335 = 8'h7 == io_state_in_7 ? 8'h9 : _GEN_3334; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3336 = 8'h8 == io_state_in_7 ? 8'h18 : _GEN_3335; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3337 = 8'h9 == io_state_in_7 ? 8'h1b : _GEN_3336; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3338 = 8'ha == io_state_in_7 ? 8'h1e : _GEN_3337; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3339 = 8'hb == io_state_in_7 ? 8'h1d : _GEN_3338; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3340 = 8'hc == io_state_in_7 ? 8'h14 : _GEN_3339; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3341 = 8'hd == io_state_in_7 ? 8'h17 : _GEN_3340; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3342 = 8'he == io_state_in_7 ? 8'h12 : _GEN_3341; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3343 = 8'hf == io_state_in_7 ? 8'h11 : _GEN_3342; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3344 = 8'h10 == io_state_in_7 ? 8'h30 : _GEN_3343; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3345 = 8'h11 == io_state_in_7 ? 8'h33 : _GEN_3344; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3346 = 8'h12 == io_state_in_7 ? 8'h36 : _GEN_3345; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3347 = 8'h13 == io_state_in_7 ? 8'h35 : _GEN_3346; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3348 = 8'h14 == io_state_in_7 ? 8'h3c : _GEN_3347; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3349 = 8'h15 == io_state_in_7 ? 8'h3f : _GEN_3348; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3350 = 8'h16 == io_state_in_7 ? 8'h3a : _GEN_3349; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3351 = 8'h17 == io_state_in_7 ? 8'h39 : _GEN_3350; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3352 = 8'h18 == io_state_in_7 ? 8'h28 : _GEN_3351; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3353 = 8'h19 == io_state_in_7 ? 8'h2b : _GEN_3352; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3354 = 8'h1a == io_state_in_7 ? 8'h2e : _GEN_3353; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3355 = 8'h1b == io_state_in_7 ? 8'h2d : _GEN_3354; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3356 = 8'h1c == io_state_in_7 ? 8'h24 : _GEN_3355; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3357 = 8'h1d == io_state_in_7 ? 8'h27 : _GEN_3356; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3358 = 8'h1e == io_state_in_7 ? 8'h22 : _GEN_3357; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3359 = 8'h1f == io_state_in_7 ? 8'h21 : _GEN_3358; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3360 = 8'h20 == io_state_in_7 ? 8'h60 : _GEN_3359; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3361 = 8'h21 == io_state_in_7 ? 8'h63 : _GEN_3360; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3362 = 8'h22 == io_state_in_7 ? 8'h66 : _GEN_3361; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3363 = 8'h23 == io_state_in_7 ? 8'h65 : _GEN_3362; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3364 = 8'h24 == io_state_in_7 ? 8'h6c : _GEN_3363; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3365 = 8'h25 == io_state_in_7 ? 8'h6f : _GEN_3364; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3366 = 8'h26 == io_state_in_7 ? 8'h6a : _GEN_3365; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3367 = 8'h27 == io_state_in_7 ? 8'h69 : _GEN_3366; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3368 = 8'h28 == io_state_in_7 ? 8'h78 : _GEN_3367; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3369 = 8'h29 == io_state_in_7 ? 8'h7b : _GEN_3368; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3370 = 8'h2a == io_state_in_7 ? 8'h7e : _GEN_3369; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3371 = 8'h2b == io_state_in_7 ? 8'h7d : _GEN_3370; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3372 = 8'h2c == io_state_in_7 ? 8'h74 : _GEN_3371; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3373 = 8'h2d == io_state_in_7 ? 8'h77 : _GEN_3372; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3374 = 8'h2e == io_state_in_7 ? 8'h72 : _GEN_3373; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3375 = 8'h2f == io_state_in_7 ? 8'h71 : _GEN_3374; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3376 = 8'h30 == io_state_in_7 ? 8'h50 : _GEN_3375; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3377 = 8'h31 == io_state_in_7 ? 8'h53 : _GEN_3376; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3378 = 8'h32 == io_state_in_7 ? 8'h56 : _GEN_3377; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3379 = 8'h33 == io_state_in_7 ? 8'h55 : _GEN_3378; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3380 = 8'h34 == io_state_in_7 ? 8'h5c : _GEN_3379; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3381 = 8'h35 == io_state_in_7 ? 8'h5f : _GEN_3380; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3382 = 8'h36 == io_state_in_7 ? 8'h5a : _GEN_3381; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3383 = 8'h37 == io_state_in_7 ? 8'h59 : _GEN_3382; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3384 = 8'h38 == io_state_in_7 ? 8'h48 : _GEN_3383; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3385 = 8'h39 == io_state_in_7 ? 8'h4b : _GEN_3384; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3386 = 8'h3a == io_state_in_7 ? 8'h4e : _GEN_3385; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3387 = 8'h3b == io_state_in_7 ? 8'h4d : _GEN_3386; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3388 = 8'h3c == io_state_in_7 ? 8'h44 : _GEN_3387; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3389 = 8'h3d == io_state_in_7 ? 8'h47 : _GEN_3388; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3390 = 8'h3e == io_state_in_7 ? 8'h42 : _GEN_3389; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3391 = 8'h3f == io_state_in_7 ? 8'h41 : _GEN_3390; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3392 = 8'h40 == io_state_in_7 ? 8'hc0 : _GEN_3391; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3393 = 8'h41 == io_state_in_7 ? 8'hc3 : _GEN_3392; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3394 = 8'h42 == io_state_in_7 ? 8'hc6 : _GEN_3393; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3395 = 8'h43 == io_state_in_7 ? 8'hc5 : _GEN_3394; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3396 = 8'h44 == io_state_in_7 ? 8'hcc : _GEN_3395; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3397 = 8'h45 == io_state_in_7 ? 8'hcf : _GEN_3396; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3398 = 8'h46 == io_state_in_7 ? 8'hca : _GEN_3397; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3399 = 8'h47 == io_state_in_7 ? 8'hc9 : _GEN_3398; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3400 = 8'h48 == io_state_in_7 ? 8'hd8 : _GEN_3399; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3401 = 8'h49 == io_state_in_7 ? 8'hdb : _GEN_3400; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3402 = 8'h4a == io_state_in_7 ? 8'hde : _GEN_3401; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3403 = 8'h4b == io_state_in_7 ? 8'hdd : _GEN_3402; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3404 = 8'h4c == io_state_in_7 ? 8'hd4 : _GEN_3403; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3405 = 8'h4d == io_state_in_7 ? 8'hd7 : _GEN_3404; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3406 = 8'h4e == io_state_in_7 ? 8'hd2 : _GEN_3405; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3407 = 8'h4f == io_state_in_7 ? 8'hd1 : _GEN_3406; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3408 = 8'h50 == io_state_in_7 ? 8'hf0 : _GEN_3407; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3409 = 8'h51 == io_state_in_7 ? 8'hf3 : _GEN_3408; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3410 = 8'h52 == io_state_in_7 ? 8'hf6 : _GEN_3409; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3411 = 8'h53 == io_state_in_7 ? 8'hf5 : _GEN_3410; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3412 = 8'h54 == io_state_in_7 ? 8'hfc : _GEN_3411; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3413 = 8'h55 == io_state_in_7 ? 8'hff : _GEN_3412; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3414 = 8'h56 == io_state_in_7 ? 8'hfa : _GEN_3413; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3415 = 8'h57 == io_state_in_7 ? 8'hf9 : _GEN_3414; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3416 = 8'h58 == io_state_in_7 ? 8'he8 : _GEN_3415; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3417 = 8'h59 == io_state_in_7 ? 8'heb : _GEN_3416; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3418 = 8'h5a == io_state_in_7 ? 8'hee : _GEN_3417; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3419 = 8'h5b == io_state_in_7 ? 8'hed : _GEN_3418; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3420 = 8'h5c == io_state_in_7 ? 8'he4 : _GEN_3419; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3421 = 8'h5d == io_state_in_7 ? 8'he7 : _GEN_3420; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3422 = 8'h5e == io_state_in_7 ? 8'he2 : _GEN_3421; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3423 = 8'h5f == io_state_in_7 ? 8'he1 : _GEN_3422; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3424 = 8'h60 == io_state_in_7 ? 8'ha0 : _GEN_3423; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3425 = 8'h61 == io_state_in_7 ? 8'ha3 : _GEN_3424; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3426 = 8'h62 == io_state_in_7 ? 8'ha6 : _GEN_3425; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3427 = 8'h63 == io_state_in_7 ? 8'ha5 : _GEN_3426; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3428 = 8'h64 == io_state_in_7 ? 8'hac : _GEN_3427; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3429 = 8'h65 == io_state_in_7 ? 8'haf : _GEN_3428; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3430 = 8'h66 == io_state_in_7 ? 8'haa : _GEN_3429; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3431 = 8'h67 == io_state_in_7 ? 8'ha9 : _GEN_3430; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3432 = 8'h68 == io_state_in_7 ? 8'hb8 : _GEN_3431; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3433 = 8'h69 == io_state_in_7 ? 8'hbb : _GEN_3432; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3434 = 8'h6a == io_state_in_7 ? 8'hbe : _GEN_3433; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3435 = 8'h6b == io_state_in_7 ? 8'hbd : _GEN_3434; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3436 = 8'h6c == io_state_in_7 ? 8'hb4 : _GEN_3435; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3437 = 8'h6d == io_state_in_7 ? 8'hb7 : _GEN_3436; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3438 = 8'h6e == io_state_in_7 ? 8'hb2 : _GEN_3437; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3439 = 8'h6f == io_state_in_7 ? 8'hb1 : _GEN_3438; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3440 = 8'h70 == io_state_in_7 ? 8'h90 : _GEN_3439; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3441 = 8'h71 == io_state_in_7 ? 8'h93 : _GEN_3440; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3442 = 8'h72 == io_state_in_7 ? 8'h96 : _GEN_3441; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3443 = 8'h73 == io_state_in_7 ? 8'h95 : _GEN_3442; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3444 = 8'h74 == io_state_in_7 ? 8'h9c : _GEN_3443; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3445 = 8'h75 == io_state_in_7 ? 8'h9f : _GEN_3444; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3446 = 8'h76 == io_state_in_7 ? 8'h9a : _GEN_3445; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3447 = 8'h77 == io_state_in_7 ? 8'h99 : _GEN_3446; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3448 = 8'h78 == io_state_in_7 ? 8'h88 : _GEN_3447; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3449 = 8'h79 == io_state_in_7 ? 8'h8b : _GEN_3448; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3450 = 8'h7a == io_state_in_7 ? 8'h8e : _GEN_3449; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3451 = 8'h7b == io_state_in_7 ? 8'h8d : _GEN_3450; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3452 = 8'h7c == io_state_in_7 ? 8'h84 : _GEN_3451; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3453 = 8'h7d == io_state_in_7 ? 8'h87 : _GEN_3452; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3454 = 8'h7e == io_state_in_7 ? 8'h82 : _GEN_3453; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3455 = 8'h7f == io_state_in_7 ? 8'h81 : _GEN_3454; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3456 = 8'h80 == io_state_in_7 ? 8'h9b : _GEN_3455; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3457 = 8'h81 == io_state_in_7 ? 8'h98 : _GEN_3456; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3458 = 8'h82 == io_state_in_7 ? 8'h9d : _GEN_3457; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3459 = 8'h83 == io_state_in_7 ? 8'h9e : _GEN_3458; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3460 = 8'h84 == io_state_in_7 ? 8'h97 : _GEN_3459; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3461 = 8'h85 == io_state_in_7 ? 8'h94 : _GEN_3460; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3462 = 8'h86 == io_state_in_7 ? 8'h91 : _GEN_3461; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3463 = 8'h87 == io_state_in_7 ? 8'h92 : _GEN_3462; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3464 = 8'h88 == io_state_in_7 ? 8'h83 : _GEN_3463; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3465 = 8'h89 == io_state_in_7 ? 8'h80 : _GEN_3464; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3466 = 8'h8a == io_state_in_7 ? 8'h85 : _GEN_3465; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3467 = 8'h8b == io_state_in_7 ? 8'h86 : _GEN_3466; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3468 = 8'h8c == io_state_in_7 ? 8'h8f : _GEN_3467; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3469 = 8'h8d == io_state_in_7 ? 8'h8c : _GEN_3468; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3470 = 8'h8e == io_state_in_7 ? 8'h89 : _GEN_3469; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3471 = 8'h8f == io_state_in_7 ? 8'h8a : _GEN_3470; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3472 = 8'h90 == io_state_in_7 ? 8'hab : _GEN_3471; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3473 = 8'h91 == io_state_in_7 ? 8'ha8 : _GEN_3472; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3474 = 8'h92 == io_state_in_7 ? 8'had : _GEN_3473; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3475 = 8'h93 == io_state_in_7 ? 8'hae : _GEN_3474; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3476 = 8'h94 == io_state_in_7 ? 8'ha7 : _GEN_3475; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3477 = 8'h95 == io_state_in_7 ? 8'ha4 : _GEN_3476; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3478 = 8'h96 == io_state_in_7 ? 8'ha1 : _GEN_3477; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3479 = 8'h97 == io_state_in_7 ? 8'ha2 : _GEN_3478; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3480 = 8'h98 == io_state_in_7 ? 8'hb3 : _GEN_3479; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3481 = 8'h99 == io_state_in_7 ? 8'hb0 : _GEN_3480; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3482 = 8'h9a == io_state_in_7 ? 8'hb5 : _GEN_3481; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3483 = 8'h9b == io_state_in_7 ? 8'hb6 : _GEN_3482; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3484 = 8'h9c == io_state_in_7 ? 8'hbf : _GEN_3483; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3485 = 8'h9d == io_state_in_7 ? 8'hbc : _GEN_3484; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3486 = 8'h9e == io_state_in_7 ? 8'hb9 : _GEN_3485; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3487 = 8'h9f == io_state_in_7 ? 8'hba : _GEN_3486; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3488 = 8'ha0 == io_state_in_7 ? 8'hfb : _GEN_3487; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3489 = 8'ha1 == io_state_in_7 ? 8'hf8 : _GEN_3488; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3490 = 8'ha2 == io_state_in_7 ? 8'hfd : _GEN_3489; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3491 = 8'ha3 == io_state_in_7 ? 8'hfe : _GEN_3490; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3492 = 8'ha4 == io_state_in_7 ? 8'hf7 : _GEN_3491; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3493 = 8'ha5 == io_state_in_7 ? 8'hf4 : _GEN_3492; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3494 = 8'ha6 == io_state_in_7 ? 8'hf1 : _GEN_3493; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3495 = 8'ha7 == io_state_in_7 ? 8'hf2 : _GEN_3494; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3496 = 8'ha8 == io_state_in_7 ? 8'he3 : _GEN_3495; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3497 = 8'ha9 == io_state_in_7 ? 8'he0 : _GEN_3496; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3498 = 8'haa == io_state_in_7 ? 8'he5 : _GEN_3497; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3499 = 8'hab == io_state_in_7 ? 8'he6 : _GEN_3498; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3500 = 8'hac == io_state_in_7 ? 8'hef : _GEN_3499; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3501 = 8'had == io_state_in_7 ? 8'hec : _GEN_3500; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3502 = 8'hae == io_state_in_7 ? 8'he9 : _GEN_3501; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3503 = 8'haf == io_state_in_7 ? 8'hea : _GEN_3502; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3504 = 8'hb0 == io_state_in_7 ? 8'hcb : _GEN_3503; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3505 = 8'hb1 == io_state_in_7 ? 8'hc8 : _GEN_3504; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3506 = 8'hb2 == io_state_in_7 ? 8'hcd : _GEN_3505; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3507 = 8'hb3 == io_state_in_7 ? 8'hce : _GEN_3506; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3508 = 8'hb4 == io_state_in_7 ? 8'hc7 : _GEN_3507; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3509 = 8'hb5 == io_state_in_7 ? 8'hc4 : _GEN_3508; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3510 = 8'hb6 == io_state_in_7 ? 8'hc1 : _GEN_3509; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3511 = 8'hb7 == io_state_in_7 ? 8'hc2 : _GEN_3510; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3512 = 8'hb8 == io_state_in_7 ? 8'hd3 : _GEN_3511; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3513 = 8'hb9 == io_state_in_7 ? 8'hd0 : _GEN_3512; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3514 = 8'hba == io_state_in_7 ? 8'hd5 : _GEN_3513; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3515 = 8'hbb == io_state_in_7 ? 8'hd6 : _GEN_3514; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3516 = 8'hbc == io_state_in_7 ? 8'hdf : _GEN_3515; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3517 = 8'hbd == io_state_in_7 ? 8'hdc : _GEN_3516; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3518 = 8'hbe == io_state_in_7 ? 8'hd9 : _GEN_3517; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3519 = 8'hbf == io_state_in_7 ? 8'hda : _GEN_3518; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3520 = 8'hc0 == io_state_in_7 ? 8'h5b : _GEN_3519; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3521 = 8'hc1 == io_state_in_7 ? 8'h58 : _GEN_3520; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3522 = 8'hc2 == io_state_in_7 ? 8'h5d : _GEN_3521; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3523 = 8'hc3 == io_state_in_7 ? 8'h5e : _GEN_3522; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3524 = 8'hc4 == io_state_in_7 ? 8'h57 : _GEN_3523; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3525 = 8'hc5 == io_state_in_7 ? 8'h54 : _GEN_3524; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3526 = 8'hc6 == io_state_in_7 ? 8'h51 : _GEN_3525; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3527 = 8'hc7 == io_state_in_7 ? 8'h52 : _GEN_3526; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3528 = 8'hc8 == io_state_in_7 ? 8'h43 : _GEN_3527; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3529 = 8'hc9 == io_state_in_7 ? 8'h40 : _GEN_3528; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3530 = 8'hca == io_state_in_7 ? 8'h45 : _GEN_3529; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3531 = 8'hcb == io_state_in_7 ? 8'h46 : _GEN_3530; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3532 = 8'hcc == io_state_in_7 ? 8'h4f : _GEN_3531; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3533 = 8'hcd == io_state_in_7 ? 8'h4c : _GEN_3532; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3534 = 8'hce == io_state_in_7 ? 8'h49 : _GEN_3533; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3535 = 8'hcf == io_state_in_7 ? 8'h4a : _GEN_3534; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3536 = 8'hd0 == io_state_in_7 ? 8'h6b : _GEN_3535; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3537 = 8'hd1 == io_state_in_7 ? 8'h68 : _GEN_3536; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3538 = 8'hd2 == io_state_in_7 ? 8'h6d : _GEN_3537; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3539 = 8'hd3 == io_state_in_7 ? 8'h6e : _GEN_3538; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3540 = 8'hd4 == io_state_in_7 ? 8'h67 : _GEN_3539; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3541 = 8'hd5 == io_state_in_7 ? 8'h64 : _GEN_3540; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3542 = 8'hd6 == io_state_in_7 ? 8'h61 : _GEN_3541; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3543 = 8'hd7 == io_state_in_7 ? 8'h62 : _GEN_3542; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3544 = 8'hd8 == io_state_in_7 ? 8'h73 : _GEN_3543; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3545 = 8'hd9 == io_state_in_7 ? 8'h70 : _GEN_3544; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3546 = 8'hda == io_state_in_7 ? 8'h75 : _GEN_3545; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3547 = 8'hdb == io_state_in_7 ? 8'h76 : _GEN_3546; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3548 = 8'hdc == io_state_in_7 ? 8'h7f : _GEN_3547; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3549 = 8'hdd == io_state_in_7 ? 8'h7c : _GEN_3548; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3550 = 8'hde == io_state_in_7 ? 8'h79 : _GEN_3549; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3551 = 8'hdf == io_state_in_7 ? 8'h7a : _GEN_3550; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3552 = 8'he0 == io_state_in_7 ? 8'h3b : _GEN_3551; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3553 = 8'he1 == io_state_in_7 ? 8'h38 : _GEN_3552; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3554 = 8'he2 == io_state_in_7 ? 8'h3d : _GEN_3553; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3555 = 8'he3 == io_state_in_7 ? 8'h3e : _GEN_3554; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3556 = 8'he4 == io_state_in_7 ? 8'h37 : _GEN_3555; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3557 = 8'he5 == io_state_in_7 ? 8'h34 : _GEN_3556; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3558 = 8'he6 == io_state_in_7 ? 8'h31 : _GEN_3557; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3559 = 8'he7 == io_state_in_7 ? 8'h32 : _GEN_3558; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3560 = 8'he8 == io_state_in_7 ? 8'h23 : _GEN_3559; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3561 = 8'he9 == io_state_in_7 ? 8'h20 : _GEN_3560; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3562 = 8'hea == io_state_in_7 ? 8'h25 : _GEN_3561; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3563 = 8'heb == io_state_in_7 ? 8'h26 : _GEN_3562; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3564 = 8'hec == io_state_in_7 ? 8'h2f : _GEN_3563; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3565 = 8'hed == io_state_in_7 ? 8'h2c : _GEN_3564; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3566 = 8'hee == io_state_in_7 ? 8'h29 : _GEN_3565; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3567 = 8'hef == io_state_in_7 ? 8'h2a : _GEN_3566; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3568 = 8'hf0 == io_state_in_7 ? 8'hb : _GEN_3567; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3569 = 8'hf1 == io_state_in_7 ? 8'h8 : _GEN_3568; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3570 = 8'hf2 == io_state_in_7 ? 8'hd : _GEN_3569; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3571 = 8'hf3 == io_state_in_7 ? 8'he : _GEN_3570; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3572 = 8'hf4 == io_state_in_7 ? 8'h7 : _GEN_3571; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3573 = 8'hf5 == io_state_in_7 ? 8'h4 : _GEN_3572; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3574 = 8'hf6 == io_state_in_7 ? 8'h1 : _GEN_3573; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3575 = 8'hf7 == io_state_in_7 ? 8'h2 : _GEN_3574; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3576 = 8'hf8 == io_state_in_7 ? 8'h13 : _GEN_3575; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3577 = 8'hf9 == io_state_in_7 ? 8'h10 : _GEN_3576; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3578 = 8'hfa == io_state_in_7 ? 8'h15 : _GEN_3577; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3579 = 8'hfb == io_state_in_7 ? 8'h16 : _GEN_3578; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3580 = 8'hfc == io_state_in_7 ? 8'h1f : _GEN_3579; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3581 = 8'hfd == io_state_in_7 ? 8'h1c : _GEN_3580; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3582 = 8'hfe == io_state_in_7 ? 8'h19 : _GEN_3581; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3583 = 8'hff == io_state_in_7 ? 8'h1a : _GEN_3582; // @[MixColumns.scala 132:{75,75}]
  wire [7:0] _GEN_3585 = 8'h1 == io_state_in_4 ? 8'h3 : 8'h0; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3586 = 8'h2 == io_state_in_4 ? 8'h6 : _GEN_3585; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3587 = 8'h3 == io_state_in_4 ? 8'h5 : _GEN_3586; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3588 = 8'h4 == io_state_in_4 ? 8'hc : _GEN_3587; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3589 = 8'h5 == io_state_in_4 ? 8'hf : _GEN_3588; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3590 = 8'h6 == io_state_in_4 ? 8'ha : _GEN_3589; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3591 = 8'h7 == io_state_in_4 ? 8'h9 : _GEN_3590; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3592 = 8'h8 == io_state_in_4 ? 8'h18 : _GEN_3591; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3593 = 8'h9 == io_state_in_4 ? 8'h1b : _GEN_3592; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3594 = 8'ha == io_state_in_4 ? 8'h1e : _GEN_3593; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3595 = 8'hb == io_state_in_4 ? 8'h1d : _GEN_3594; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3596 = 8'hc == io_state_in_4 ? 8'h14 : _GEN_3595; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3597 = 8'hd == io_state_in_4 ? 8'h17 : _GEN_3596; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3598 = 8'he == io_state_in_4 ? 8'h12 : _GEN_3597; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3599 = 8'hf == io_state_in_4 ? 8'h11 : _GEN_3598; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3600 = 8'h10 == io_state_in_4 ? 8'h30 : _GEN_3599; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3601 = 8'h11 == io_state_in_4 ? 8'h33 : _GEN_3600; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3602 = 8'h12 == io_state_in_4 ? 8'h36 : _GEN_3601; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3603 = 8'h13 == io_state_in_4 ? 8'h35 : _GEN_3602; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3604 = 8'h14 == io_state_in_4 ? 8'h3c : _GEN_3603; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3605 = 8'h15 == io_state_in_4 ? 8'h3f : _GEN_3604; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3606 = 8'h16 == io_state_in_4 ? 8'h3a : _GEN_3605; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3607 = 8'h17 == io_state_in_4 ? 8'h39 : _GEN_3606; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3608 = 8'h18 == io_state_in_4 ? 8'h28 : _GEN_3607; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3609 = 8'h19 == io_state_in_4 ? 8'h2b : _GEN_3608; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3610 = 8'h1a == io_state_in_4 ? 8'h2e : _GEN_3609; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3611 = 8'h1b == io_state_in_4 ? 8'h2d : _GEN_3610; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3612 = 8'h1c == io_state_in_4 ? 8'h24 : _GEN_3611; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3613 = 8'h1d == io_state_in_4 ? 8'h27 : _GEN_3612; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3614 = 8'h1e == io_state_in_4 ? 8'h22 : _GEN_3613; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3615 = 8'h1f == io_state_in_4 ? 8'h21 : _GEN_3614; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3616 = 8'h20 == io_state_in_4 ? 8'h60 : _GEN_3615; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3617 = 8'h21 == io_state_in_4 ? 8'h63 : _GEN_3616; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3618 = 8'h22 == io_state_in_4 ? 8'h66 : _GEN_3617; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3619 = 8'h23 == io_state_in_4 ? 8'h65 : _GEN_3618; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3620 = 8'h24 == io_state_in_4 ? 8'h6c : _GEN_3619; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3621 = 8'h25 == io_state_in_4 ? 8'h6f : _GEN_3620; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3622 = 8'h26 == io_state_in_4 ? 8'h6a : _GEN_3621; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3623 = 8'h27 == io_state_in_4 ? 8'h69 : _GEN_3622; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3624 = 8'h28 == io_state_in_4 ? 8'h78 : _GEN_3623; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3625 = 8'h29 == io_state_in_4 ? 8'h7b : _GEN_3624; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3626 = 8'h2a == io_state_in_4 ? 8'h7e : _GEN_3625; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3627 = 8'h2b == io_state_in_4 ? 8'h7d : _GEN_3626; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3628 = 8'h2c == io_state_in_4 ? 8'h74 : _GEN_3627; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3629 = 8'h2d == io_state_in_4 ? 8'h77 : _GEN_3628; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3630 = 8'h2e == io_state_in_4 ? 8'h72 : _GEN_3629; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3631 = 8'h2f == io_state_in_4 ? 8'h71 : _GEN_3630; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3632 = 8'h30 == io_state_in_4 ? 8'h50 : _GEN_3631; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3633 = 8'h31 == io_state_in_4 ? 8'h53 : _GEN_3632; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3634 = 8'h32 == io_state_in_4 ? 8'h56 : _GEN_3633; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3635 = 8'h33 == io_state_in_4 ? 8'h55 : _GEN_3634; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3636 = 8'h34 == io_state_in_4 ? 8'h5c : _GEN_3635; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3637 = 8'h35 == io_state_in_4 ? 8'h5f : _GEN_3636; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3638 = 8'h36 == io_state_in_4 ? 8'h5a : _GEN_3637; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3639 = 8'h37 == io_state_in_4 ? 8'h59 : _GEN_3638; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3640 = 8'h38 == io_state_in_4 ? 8'h48 : _GEN_3639; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3641 = 8'h39 == io_state_in_4 ? 8'h4b : _GEN_3640; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3642 = 8'h3a == io_state_in_4 ? 8'h4e : _GEN_3641; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3643 = 8'h3b == io_state_in_4 ? 8'h4d : _GEN_3642; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3644 = 8'h3c == io_state_in_4 ? 8'h44 : _GEN_3643; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3645 = 8'h3d == io_state_in_4 ? 8'h47 : _GEN_3644; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3646 = 8'h3e == io_state_in_4 ? 8'h42 : _GEN_3645; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3647 = 8'h3f == io_state_in_4 ? 8'h41 : _GEN_3646; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3648 = 8'h40 == io_state_in_4 ? 8'hc0 : _GEN_3647; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3649 = 8'h41 == io_state_in_4 ? 8'hc3 : _GEN_3648; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3650 = 8'h42 == io_state_in_4 ? 8'hc6 : _GEN_3649; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3651 = 8'h43 == io_state_in_4 ? 8'hc5 : _GEN_3650; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3652 = 8'h44 == io_state_in_4 ? 8'hcc : _GEN_3651; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3653 = 8'h45 == io_state_in_4 ? 8'hcf : _GEN_3652; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3654 = 8'h46 == io_state_in_4 ? 8'hca : _GEN_3653; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3655 = 8'h47 == io_state_in_4 ? 8'hc9 : _GEN_3654; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3656 = 8'h48 == io_state_in_4 ? 8'hd8 : _GEN_3655; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3657 = 8'h49 == io_state_in_4 ? 8'hdb : _GEN_3656; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3658 = 8'h4a == io_state_in_4 ? 8'hde : _GEN_3657; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3659 = 8'h4b == io_state_in_4 ? 8'hdd : _GEN_3658; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3660 = 8'h4c == io_state_in_4 ? 8'hd4 : _GEN_3659; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3661 = 8'h4d == io_state_in_4 ? 8'hd7 : _GEN_3660; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3662 = 8'h4e == io_state_in_4 ? 8'hd2 : _GEN_3661; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3663 = 8'h4f == io_state_in_4 ? 8'hd1 : _GEN_3662; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3664 = 8'h50 == io_state_in_4 ? 8'hf0 : _GEN_3663; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3665 = 8'h51 == io_state_in_4 ? 8'hf3 : _GEN_3664; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3666 = 8'h52 == io_state_in_4 ? 8'hf6 : _GEN_3665; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3667 = 8'h53 == io_state_in_4 ? 8'hf5 : _GEN_3666; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3668 = 8'h54 == io_state_in_4 ? 8'hfc : _GEN_3667; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3669 = 8'h55 == io_state_in_4 ? 8'hff : _GEN_3668; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3670 = 8'h56 == io_state_in_4 ? 8'hfa : _GEN_3669; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3671 = 8'h57 == io_state_in_4 ? 8'hf9 : _GEN_3670; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3672 = 8'h58 == io_state_in_4 ? 8'he8 : _GEN_3671; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3673 = 8'h59 == io_state_in_4 ? 8'heb : _GEN_3672; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3674 = 8'h5a == io_state_in_4 ? 8'hee : _GEN_3673; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3675 = 8'h5b == io_state_in_4 ? 8'hed : _GEN_3674; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3676 = 8'h5c == io_state_in_4 ? 8'he4 : _GEN_3675; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3677 = 8'h5d == io_state_in_4 ? 8'he7 : _GEN_3676; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3678 = 8'h5e == io_state_in_4 ? 8'he2 : _GEN_3677; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3679 = 8'h5f == io_state_in_4 ? 8'he1 : _GEN_3678; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3680 = 8'h60 == io_state_in_4 ? 8'ha0 : _GEN_3679; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3681 = 8'h61 == io_state_in_4 ? 8'ha3 : _GEN_3680; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3682 = 8'h62 == io_state_in_4 ? 8'ha6 : _GEN_3681; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3683 = 8'h63 == io_state_in_4 ? 8'ha5 : _GEN_3682; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3684 = 8'h64 == io_state_in_4 ? 8'hac : _GEN_3683; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3685 = 8'h65 == io_state_in_4 ? 8'haf : _GEN_3684; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3686 = 8'h66 == io_state_in_4 ? 8'haa : _GEN_3685; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3687 = 8'h67 == io_state_in_4 ? 8'ha9 : _GEN_3686; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3688 = 8'h68 == io_state_in_4 ? 8'hb8 : _GEN_3687; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3689 = 8'h69 == io_state_in_4 ? 8'hbb : _GEN_3688; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3690 = 8'h6a == io_state_in_4 ? 8'hbe : _GEN_3689; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3691 = 8'h6b == io_state_in_4 ? 8'hbd : _GEN_3690; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3692 = 8'h6c == io_state_in_4 ? 8'hb4 : _GEN_3691; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3693 = 8'h6d == io_state_in_4 ? 8'hb7 : _GEN_3692; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3694 = 8'h6e == io_state_in_4 ? 8'hb2 : _GEN_3693; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3695 = 8'h6f == io_state_in_4 ? 8'hb1 : _GEN_3694; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3696 = 8'h70 == io_state_in_4 ? 8'h90 : _GEN_3695; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3697 = 8'h71 == io_state_in_4 ? 8'h93 : _GEN_3696; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3698 = 8'h72 == io_state_in_4 ? 8'h96 : _GEN_3697; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3699 = 8'h73 == io_state_in_4 ? 8'h95 : _GEN_3698; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3700 = 8'h74 == io_state_in_4 ? 8'h9c : _GEN_3699; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3701 = 8'h75 == io_state_in_4 ? 8'h9f : _GEN_3700; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3702 = 8'h76 == io_state_in_4 ? 8'h9a : _GEN_3701; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3703 = 8'h77 == io_state_in_4 ? 8'h99 : _GEN_3702; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3704 = 8'h78 == io_state_in_4 ? 8'h88 : _GEN_3703; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3705 = 8'h79 == io_state_in_4 ? 8'h8b : _GEN_3704; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3706 = 8'h7a == io_state_in_4 ? 8'h8e : _GEN_3705; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3707 = 8'h7b == io_state_in_4 ? 8'h8d : _GEN_3706; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3708 = 8'h7c == io_state_in_4 ? 8'h84 : _GEN_3707; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3709 = 8'h7d == io_state_in_4 ? 8'h87 : _GEN_3708; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3710 = 8'h7e == io_state_in_4 ? 8'h82 : _GEN_3709; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3711 = 8'h7f == io_state_in_4 ? 8'h81 : _GEN_3710; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3712 = 8'h80 == io_state_in_4 ? 8'h9b : _GEN_3711; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3713 = 8'h81 == io_state_in_4 ? 8'h98 : _GEN_3712; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3714 = 8'h82 == io_state_in_4 ? 8'h9d : _GEN_3713; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3715 = 8'h83 == io_state_in_4 ? 8'h9e : _GEN_3714; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3716 = 8'h84 == io_state_in_4 ? 8'h97 : _GEN_3715; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3717 = 8'h85 == io_state_in_4 ? 8'h94 : _GEN_3716; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3718 = 8'h86 == io_state_in_4 ? 8'h91 : _GEN_3717; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3719 = 8'h87 == io_state_in_4 ? 8'h92 : _GEN_3718; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3720 = 8'h88 == io_state_in_4 ? 8'h83 : _GEN_3719; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3721 = 8'h89 == io_state_in_4 ? 8'h80 : _GEN_3720; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3722 = 8'h8a == io_state_in_4 ? 8'h85 : _GEN_3721; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3723 = 8'h8b == io_state_in_4 ? 8'h86 : _GEN_3722; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3724 = 8'h8c == io_state_in_4 ? 8'h8f : _GEN_3723; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3725 = 8'h8d == io_state_in_4 ? 8'h8c : _GEN_3724; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3726 = 8'h8e == io_state_in_4 ? 8'h89 : _GEN_3725; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3727 = 8'h8f == io_state_in_4 ? 8'h8a : _GEN_3726; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3728 = 8'h90 == io_state_in_4 ? 8'hab : _GEN_3727; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3729 = 8'h91 == io_state_in_4 ? 8'ha8 : _GEN_3728; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3730 = 8'h92 == io_state_in_4 ? 8'had : _GEN_3729; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3731 = 8'h93 == io_state_in_4 ? 8'hae : _GEN_3730; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3732 = 8'h94 == io_state_in_4 ? 8'ha7 : _GEN_3731; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3733 = 8'h95 == io_state_in_4 ? 8'ha4 : _GEN_3732; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3734 = 8'h96 == io_state_in_4 ? 8'ha1 : _GEN_3733; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3735 = 8'h97 == io_state_in_4 ? 8'ha2 : _GEN_3734; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3736 = 8'h98 == io_state_in_4 ? 8'hb3 : _GEN_3735; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3737 = 8'h99 == io_state_in_4 ? 8'hb0 : _GEN_3736; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3738 = 8'h9a == io_state_in_4 ? 8'hb5 : _GEN_3737; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3739 = 8'h9b == io_state_in_4 ? 8'hb6 : _GEN_3738; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3740 = 8'h9c == io_state_in_4 ? 8'hbf : _GEN_3739; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3741 = 8'h9d == io_state_in_4 ? 8'hbc : _GEN_3740; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3742 = 8'h9e == io_state_in_4 ? 8'hb9 : _GEN_3741; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3743 = 8'h9f == io_state_in_4 ? 8'hba : _GEN_3742; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3744 = 8'ha0 == io_state_in_4 ? 8'hfb : _GEN_3743; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3745 = 8'ha1 == io_state_in_4 ? 8'hf8 : _GEN_3744; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3746 = 8'ha2 == io_state_in_4 ? 8'hfd : _GEN_3745; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3747 = 8'ha3 == io_state_in_4 ? 8'hfe : _GEN_3746; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3748 = 8'ha4 == io_state_in_4 ? 8'hf7 : _GEN_3747; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3749 = 8'ha5 == io_state_in_4 ? 8'hf4 : _GEN_3748; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3750 = 8'ha6 == io_state_in_4 ? 8'hf1 : _GEN_3749; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3751 = 8'ha7 == io_state_in_4 ? 8'hf2 : _GEN_3750; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3752 = 8'ha8 == io_state_in_4 ? 8'he3 : _GEN_3751; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3753 = 8'ha9 == io_state_in_4 ? 8'he0 : _GEN_3752; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3754 = 8'haa == io_state_in_4 ? 8'he5 : _GEN_3753; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3755 = 8'hab == io_state_in_4 ? 8'he6 : _GEN_3754; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3756 = 8'hac == io_state_in_4 ? 8'hef : _GEN_3755; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3757 = 8'had == io_state_in_4 ? 8'hec : _GEN_3756; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3758 = 8'hae == io_state_in_4 ? 8'he9 : _GEN_3757; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3759 = 8'haf == io_state_in_4 ? 8'hea : _GEN_3758; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3760 = 8'hb0 == io_state_in_4 ? 8'hcb : _GEN_3759; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3761 = 8'hb1 == io_state_in_4 ? 8'hc8 : _GEN_3760; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3762 = 8'hb2 == io_state_in_4 ? 8'hcd : _GEN_3761; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3763 = 8'hb3 == io_state_in_4 ? 8'hce : _GEN_3762; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3764 = 8'hb4 == io_state_in_4 ? 8'hc7 : _GEN_3763; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3765 = 8'hb5 == io_state_in_4 ? 8'hc4 : _GEN_3764; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3766 = 8'hb6 == io_state_in_4 ? 8'hc1 : _GEN_3765; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3767 = 8'hb7 == io_state_in_4 ? 8'hc2 : _GEN_3766; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3768 = 8'hb8 == io_state_in_4 ? 8'hd3 : _GEN_3767; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3769 = 8'hb9 == io_state_in_4 ? 8'hd0 : _GEN_3768; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3770 = 8'hba == io_state_in_4 ? 8'hd5 : _GEN_3769; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3771 = 8'hbb == io_state_in_4 ? 8'hd6 : _GEN_3770; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3772 = 8'hbc == io_state_in_4 ? 8'hdf : _GEN_3771; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3773 = 8'hbd == io_state_in_4 ? 8'hdc : _GEN_3772; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3774 = 8'hbe == io_state_in_4 ? 8'hd9 : _GEN_3773; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3775 = 8'hbf == io_state_in_4 ? 8'hda : _GEN_3774; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3776 = 8'hc0 == io_state_in_4 ? 8'h5b : _GEN_3775; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3777 = 8'hc1 == io_state_in_4 ? 8'h58 : _GEN_3776; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3778 = 8'hc2 == io_state_in_4 ? 8'h5d : _GEN_3777; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3779 = 8'hc3 == io_state_in_4 ? 8'h5e : _GEN_3778; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3780 = 8'hc4 == io_state_in_4 ? 8'h57 : _GEN_3779; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3781 = 8'hc5 == io_state_in_4 ? 8'h54 : _GEN_3780; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3782 = 8'hc6 == io_state_in_4 ? 8'h51 : _GEN_3781; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3783 = 8'hc7 == io_state_in_4 ? 8'h52 : _GEN_3782; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3784 = 8'hc8 == io_state_in_4 ? 8'h43 : _GEN_3783; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3785 = 8'hc9 == io_state_in_4 ? 8'h40 : _GEN_3784; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3786 = 8'hca == io_state_in_4 ? 8'h45 : _GEN_3785; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3787 = 8'hcb == io_state_in_4 ? 8'h46 : _GEN_3786; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3788 = 8'hcc == io_state_in_4 ? 8'h4f : _GEN_3787; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3789 = 8'hcd == io_state_in_4 ? 8'h4c : _GEN_3788; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3790 = 8'hce == io_state_in_4 ? 8'h49 : _GEN_3789; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3791 = 8'hcf == io_state_in_4 ? 8'h4a : _GEN_3790; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3792 = 8'hd0 == io_state_in_4 ? 8'h6b : _GEN_3791; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3793 = 8'hd1 == io_state_in_4 ? 8'h68 : _GEN_3792; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3794 = 8'hd2 == io_state_in_4 ? 8'h6d : _GEN_3793; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3795 = 8'hd3 == io_state_in_4 ? 8'h6e : _GEN_3794; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3796 = 8'hd4 == io_state_in_4 ? 8'h67 : _GEN_3795; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3797 = 8'hd5 == io_state_in_4 ? 8'h64 : _GEN_3796; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3798 = 8'hd6 == io_state_in_4 ? 8'h61 : _GEN_3797; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3799 = 8'hd7 == io_state_in_4 ? 8'h62 : _GEN_3798; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3800 = 8'hd8 == io_state_in_4 ? 8'h73 : _GEN_3799; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3801 = 8'hd9 == io_state_in_4 ? 8'h70 : _GEN_3800; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3802 = 8'hda == io_state_in_4 ? 8'h75 : _GEN_3801; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3803 = 8'hdb == io_state_in_4 ? 8'h76 : _GEN_3802; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3804 = 8'hdc == io_state_in_4 ? 8'h7f : _GEN_3803; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3805 = 8'hdd == io_state_in_4 ? 8'h7c : _GEN_3804; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3806 = 8'hde == io_state_in_4 ? 8'h79 : _GEN_3805; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3807 = 8'hdf == io_state_in_4 ? 8'h7a : _GEN_3806; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3808 = 8'he0 == io_state_in_4 ? 8'h3b : _GEN_3807; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3809 = 8'he1 == io_state_in_4 ? 8'h38 : _GEN_3808; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3810 = 8'he2 == io_state_in_4 ? 8'h3d : _GEN_3809; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3811 = 8'he3 == io_state_in_4 ? 8'h3e : _GEN_3810; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3812 = 8'he4 == io_state_in_4 ? 8'h37 : _GEN_3811; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3813 = 8'he5 == io_state_in_4 ? 8'h34 : _GEN_3812; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3814 = 8'he6 == io_state_in_4 ? 8'h31 : _GEN_3813; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3815 = 8'he7 == io_state_in_4 ? 8'h32 : _GEN_3814; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3816 = 8'he8 == io_state_in_4 ? 8'h23 : _GEN_3815; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3817 = 8'he9 == io_state_in_4 ? 8'h20 : _GEN_3816; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3818 = 8'hea == io_state_in_4 ? 8'h25 : _GEN_3817; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3819 = 8'heb == io_state_in_4 ? 8'h26 : _GEN_3818; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3820 = 8'hec == io_state_in_4 ? 8'h2f : _GEN_3819; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3821 = 8'hed == io_state_in_4 ? 8'h2c : _GEN_3820; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3822 = 8'hee == io_state_in_4 ? 8'h29 : _GEN_3821; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3823 = 8'hef == io_state_in_4 ? 8'h2a : _GEN_3822; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3824 = 8'hf0 == io_state_in_4 ? 8'hb : _GEN_3823; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3825 = 8'hf1 == io_state_in_4 ? 8'h8 : _GEN_3824; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3826 = 8'hf2 == io_state_in_4 ? 8'hd : _GEN_3825; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3827 = 8'hf3 == io_state_in_4 ? 8'he : _GEN_3826; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3828 = 8'hf4 == io_state_in_4 ? 8'h7 : _GEN_3827; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3829 = 8'hf5 == io_state_in_4 ? 8'h4 : _GEN_3828; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3830 = 8'hf6 == io_state_in_4 ? 8'h1 : _GEN_3829; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3831 = 8'hf7 == io_state_in_4 ? 8'h2 : _GEN_3830; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3832 = 8'hf8 == io_state_in_4 ? 8'h13 : _GEN_3831; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3833 = 8'hf9 == io_state_in_4 ? 8'h10 : _GEN_3832; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3834 = 8'hfa == io_state_in_4 ? 8'h15 : _GEN_3833; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3835 = 8'hfb == io_state_in_4 ? 8'h16 : _GEN_3834; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3836 = 8'hfc == io_state_in_4 ? 8'h1f : _GEN_3835; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3837 = 8'hfd == io_state_in_4 ? 8'h1c : _GEN_3836; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3838 = 8'hfe == io_state_in_4 ? 8'h19 : _GEN_3837; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _GEN_3839 = 8'hff == io_state_in_4 ? 8'h1a : _GEN_3838; // @[MixColumns.scala 133:{41,41}]
  wire [7:0] _tmp_state_7_T = _GEN_3839 ^ io_state_in_5; // @[MixColumns.scala 133:41]
  wire [7:0] _tmp_state_7_T_1 = _tmp_state_7_T ^ io_state_in_6; // @[MixColumns.scala 133:58]
  wire [7:0] _GEN_3841 = 8'h1 == io_state_in_7 ? 8'h2 : 8'h0; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3842 = 8'h2 == io_state_in_7 ? 8'h4 : _GEN_3841; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3843 = 8'h3 == io_state_in_7 ? 8'h6 : _GEN_3842; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3844 = 8'h4 == io_state_in_7 ? 8'h8 : _GEN_3843; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3845 = 8'h5 == io_state_in_7 ? 8'ha : _GEN_3844; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3846 = 8'h6 == io_state_in_7 ? 8'hc : _GEN_3845; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3847 = 8'h7 == io_state_in_7 ? 8'he : _GEN_3846; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3848 = 8'h8 == io_state_in_7 ? 8'h10 : _GEN_3847; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3849 = 8'h9 == io_state_in_7 ? 8'h12 : _GEN_3848; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3850 = 8'ha == io_state_in_7 ? 8'h14 : _GEN_3849; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3851 = 8'hb == io_state_in_7 ? 8'h16 : _GEN_3850; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3852 = 8'hc == io_state_in_7 ? 8'h18 : _GEN_3851; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3853 = 8'hd == io_state_in_7 ? 8'h1a : _GEN_3852; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3854 = 8'he == io_state_in_7 ? 8'h1c : _GEN_3853; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3855 = 8'hf == io_state_in_7 ? 8'h1e : _GEN_3854; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3856 = 8'h10 == io_state_in_7 ? 8'h20 : _GEN_3855; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3857 = 8'h11 == io_state_in_7 ? 8'h22 : _GEN_3856; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3858 = 8'h12 == io_state_in_7 ? 8'h24 : _GEN_3857; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3859 = 8'h13 == io_state_in_7 ? 8'h26 : _GEN_3858; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3860 = 8'h14 == io_state_in_7 ? 8'h28 : _GEN_3859; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3861 = 8'h15 == io_state_in_7 ? 8'h2a : _GEN_3860; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3862 = 8'h16 == io_state_in_7 ? 8'h2c : _GEN_3861; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3863 = 8'h17 == io_state_in_7 ? 8'h2e : _GEN_3862; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3864 = 8'h18 == io_state_in_7 ? 8'h30 : _GEN_3863; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3865 = 8'h19 == io_state_in_7 ? 8'h32 : _GEN_3864; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3866 = 8'h1a == io_state_in_7 ? 8'h34 : _GEN_3865; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3867 = 8'h1b == io_state_in_7 ? 8'h36 : _GEN_3866; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3868 = 8'h1c == io_state_in_7 ? 8'h38 : _GEN_3867; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3869 = 8'h1d == io_state_in_7 ? 8'h3a : _GEN_3868; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3870 = 8'h1e == io_state_in_7 ? 8'h3c : _GEN_3869; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3871 = 8'h1f == io_state_in_7 ? 8'h3e : _GEN_3870; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3872 = 8'h20 == io_state_in_7 ? 8'h40 : _GEN_3871; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3873 = 8'h21 == io_state_in_7 ? 8'h42 : _GEN_3872; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3874 = 8'h22 == io_state_in_7 ? 8'h44 : _GEN_3873; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3875 = 8'h23 == io_state_in_7 ? 8'h46 : _GEN_3874; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3876 = 8'h24 == io_state_in_7 ? 8'h48 : _GEN_3875; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3877 = 8'h25 == io_state_in_7 ? 8'h4a : _GEN_3876; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3878 = 8'h26 == io_state_in_7 ? 8'h4c : _GEN_3877; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3879 = 8'h27 == io_state_in_7 ? 8'h4e : _GEN_3878; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3880 = 8'h28 == io_state_in_7 ? 8'h50 : _GEN_3879; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3881 = 8'h29 == io_state_in_7 ? 8'h52 : _GEN_3880; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3882 = 8'h2a == io_state_in_7 ? 8'h54 : _GEN_3881; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3883 = 8'h2b == io_state_in_7 ? 8'h56 : _GEN_3882; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3884 = 8'h2c == io_state_in_7 ? 8'h58 : _GEN_3883; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3885 = 8'h2d == io_state_in_7 ? 8'h5a : _GEN_3884; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3886 = 8'h2e == io_state_in_7 ? 8'h5c : _GEN_3885; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3887 = 8'h2f == io_state_in_7 ? 8'h5e : _GEN_3886; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3888 = 8'h30 == io_state_in_7 ? 8'h60 : _GEN_3887; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3889 = 8'h31 == io_state_in_7 ? 8'h62 : _GEN_3888; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3890 = 8'h32 == io_state_in_7 ? 8'h64 : _GEN_3889; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3891 = 8'h33 == io_state_in_7 ? 8'h66 : _GEN_3890; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3892 = 8'h34 == io_state_in_7 ? 8'h68 : _GEN_3891; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3893 = 8'h35 == io_state_in_7 ? 8'h6a : _GEN_3892; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3894 = 8'h36 == io_state_in_7 ? 8'h6c : _GEN_3893; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3895 = 8'h37 == io_state_in_7 ? 8'h6e : _GEN_3894; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3896 = 8'h38 == io_state_in_7 ? 8'h70 : _GEN_3895; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3897 = 8'h39 == io_state_in_7 ? 8'h72 : _GEN_3896; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3898 = 8'h3a == io_state_in_7 ? 8'h74 : _GEN_3897; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3899 = 8'h3b == io_state_in_7 ? 8'h76 : _GEN_3898; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3900 = 8'h3c == io_state_in_7 ? 8'h78 : _GEN_3899; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3901 = 8'h3d == io_state_in_7 ? 8'h7a : _GEN_3900; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3902 = 8'h3e == io_state_in_7 ? 8'h7c : _GEN_3901; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3903 = 8'h3f == io_state_in_7 ? 8'h7e : _GEN_3902; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3904 = 8'h40 == io_state_in_7 ? 8'h80 : _GEN_3903; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3905 = 8'h41 == io_state_in_7 ? 8'h82 : _GEN_3904; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3906 = 8'h42 == io_state_in_7 ? 8'h84 : _GEN_3905; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3907 = 8'h43 == io_state_in_7 ? 8'h86 : _GEN_3906; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3908 = 8'h44 == io_state_in_7 ? 8'h88 : _GEN_3907; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3909 = 8'h45 == io_state_in_7 ? 8'h8a : _GEN_3908; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3910 = 8'h46 == io_state_in_7 ? 8'h8c : _GEN_3909; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3911 = 8'h47 == io_state_in_7 ? 8'h8e : _GEN_3910; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3912 = 8'h48 == io_state_in_7 ? 8'h90 : _GEN_3911; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3913 = 8'h49 == io_state_in_7 ? 8'h92 : _GEN_3912; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3914 = 8'h4a == io_state_in_7 ? 8'h94 : _GEN_3913; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3915 = 8'h4b == io_state_in_7 ? 8'h96 : _GEN_3914; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3916 = 8'h4c == io_state_in_7 ? 8'h98 : _GEN_3915; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3917 = 8'h4d == io_state_in_7 ? 8'h9a : _GEN_3916; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3918 = 8'h4e == io_state_in_7 ? 8'h9c : _GEN_3917; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3919 = 8'h4f == io_state_in_7 ? 8'h9e : _GEN_3918; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3920 = 8'h50 == io_state_in_7 ? 8'ha0 : _GEN_3919; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3921 = 8'h51 == io_state_in_7 ? 8'ha2 : _GEN_3920; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3922 = 8'h52 == io_state_in_7 ? 8'ha4 : _GEN_3921; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3923 = 8'h53 == io_state_in_7 ? 8'ha6 : _GEN_3922; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3924 = 8'h54 == io_state_in_7 ? 8'ha8 : _GEN_3923; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3925 = 8'h55 == io_state_in_7 ? 8'haa : _GEN_3924; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3926 = 8'h56 == io_state_in_7 ? 8'hac : _GEN_3925; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3927 = 8'h57 == io_state_in_7 ? 8'hae : _GEN_3926; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3928 = 8'h58 == io_state_in_7 ? 8'hb0 : _GEN_3927; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3929 = 8'h59 == io_state_in_7 ? 8'hb2 : _GEN_3928; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3930 = 8'h5a == io_state_in_7 ? 8'hb4 : _GEN_3929; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3931 = 8'h5b == io_state_in_7 ? 8'hb6 : _GEN_3930; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3932 = 8'h5c == io_state_in_7 ? 8'hb8 : _GEN_3931; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3933 = 8'h5d == io_state_in_7 ? 8'hba : _GEN_3932; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3934 = 8'h5e == io_state_in_7 ? 8'hbc : _GEN_3933; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3935 = 8'h5f == io_state_in_7 ? 8'hbe : _GEN_3934; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3936 = 8'h60 == io_state_in_7 ? 8'hc0 : _GEN_3935; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3937 = 8'h61 == io_state_in_7 ? 8'hc2 : _GEN_3936; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3938 = 8'h62 == io_state_in_7 ? 8'hc4 : _GEN_3937; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3939 = 8'h63 == io_state_in_7 ? 8'hc6 : _GEN_3938; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3940 = 8'h64 == io_state_in_7 ? 8'hc8 : _GEN_3939; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3941 = 8'h65 == io_state_in_7 ? 8'hca : _GEN_3940; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3942 = 8'h66 == io_state_in_7 ? 8'hcc : _GEN_3941; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3943 = 8'h67 == io_state_in_7 ? 8'hce : _GEN_3942; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3944 = 8'h68 == io_state_in_7 ? 8'hd0 : _GEN_3943; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3945 = 8'h69 == io_state_in_7 ? 8'hd2 : _GEN_3944; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3946 = 8'h6a == io_state_in_7 ? 8'hd4 : _GEN_3945; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3947 = 8'h6b == io_state_in_7 ? 8'hd6 : _GEN_3946; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3948 = 8'h6c == io_state_in_7 ? 8'hd8 : _GEN_3947; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3949 = 8'h6d == io_state_in_7 ? 8'hda : _GEN_3948; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3950 = 8'h6e == io_state_in_7 ? 8'hdc : _GEN_3949; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3951 = 8'h6f == io_state_in_7 ? 8'hde : _GEN_3950; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3952 = 8'h70 == io_state_in_7 ? 8'he0 : _GEN_3951; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3953 = 8'h71 == io_state_in_7 ? 8'he2 : _GEN_3952; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3954 = 8'h72 == io_state_in_7 ? 8'he4 : _GEN_3953; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3955 = 8'h73 == io_state_in_7 ? 8'he6 : _GEN_3954; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3956 = 8'h74 == io_state_in_7 ? 8'he8 : _GEN_3955; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3957 = 8'h75 == io_state_in_7 ? 8'hea : _GEN_3956; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3958 = 8'h76 == io_state_in_7 ? 8'hec : _GEN_3957; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3959 = 8'h77 == io_state_in_7 ? 8'hee : _GEN_3958; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3960 = 8'h78 == io_state_in_7 ? 8'hf0 : _GEN_3959; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3961 = 8'h79 == io_state_in_7 ? 8'hf2 : _GEN_3960; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3962 = 8'h7a == io_state_in_7 ? 8'hf4 : _GEN_3961; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3963 = 8'h7b == io_state_in_7 ? 8'hf6 : _GEN_3962; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3964 = 8'h7c == io_state_in_7 ? 8'hf8 : _GEN_3963; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3965 = 8'h7d == io_state_in_7 ? 8'hfa : _GEN_3964; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3966 = 8'h7e == io_state_in_7 ? 8'hfc : _GEN_3965; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3967 = 8'h7f == io_state_in_7 ? 8'hfe : _GEN_3966; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3968 = 8'h80 == io_state_in_7 ? 8'h1b : _GEN_3967; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3969 = 8'h81 == io_state_in_7 ? 8'h19 : _GEN_3968; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3970 = 8'h82 == io_state_in_7 ? 8'h1f : _GEN_3969; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3971 = 8'h83 == io_state_in_7 ? 8'h1d : _GEN_3970; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3972 = 8'h84 == io_state_in_7 ? 8'h13 : _GEN_3971; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3973 = 8'h85 == io_state_in_7 ? 8'h11 : _GEN_3972; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3974 = 8'h86 == io_state_in_7 ? 8'h17 : _GEN_3973; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3975 = 8'h87 == io_state_in_7 ? 8'h15 : _GEN_3974; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3976 = 8'h88 == io_state_in_7 ? 8'hb : _GEN_3975; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3977 = 8'h89 == io_state_in_7 ? 8'h9 : _GEN_3976; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3978 = 8'h8a == io_state_in_7 ? 8'hf : _GEN_3977; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3979 = 8'h8b == io_state_in_7 ? 8'hd : _GEN_3978; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3980 = 8'h8c == io_state_in_7 ? 8'h3 : _GEN_3979; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3981 = 8'h8d == io_state_in_7 ? 8'h1 : _GEN_3980; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3982 = 8'h8e == io_state_in_7 ? 8'h7 : _GEN_3981; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3983 = 8'h8f == io_state_in_7 ? 8'h5 : _GEN_3982; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3984 = 8'h90 == io_state_in_7 ? 8'h3b : _GEN_3983; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3985 = 8'h91 == io_state_in_7 ? 8'h39 : _GEN_3984; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3986 = 8'h92 == io_state_in_7 ? 8'h3f : _GEN_3985; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3987 = 8'h93 == io_state_in_7 ? 8'h3d : _GEN_3986; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3988 = 8'h94 == io_state_in_7 ? 8'h33 : _GEN_3987; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3989 = 8'h95 == io_state_in_7 ? 8'h31 : _GEN_3988; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3990 = 8'h96 == io_state_in_7 ? 8'h37 : _GEN_3989; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3991 = 8'h97 == io_state_in_7 ? 8'h35 : _GEN_3990; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3992 = 8'h98 == io_state_in_7 ? 8'h2b : _GEN_3991; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3993 = 8'h99 == io_state_in_7 ? 8'h29 : _GEN_3992; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3994 = 8'h9a == io_state_in_7 ? 8'h2f : _GEN_3993; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3995 = 8'h9b == io_state_in_7 ? 8'h2d : _GEN_3994; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3996 = 8'h9c == io_state_in_7 ? 8'h23 : _GEN_3995; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3997 = 8'h9d == io_state_in_7 ? 8'h21 : _GEN_3996; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3998 = 8'h9e == io_state_in_7 ? 8'h27 : _GEN_3997; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_3999 = 8'h9f == io_state_in_7 ? 8'h25 : _GEN_3998; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4000 = 8'ha0 == io_state_in_7 ? 8'h5b : _GEN_3999; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4001 = 8'ha1 == io_state_in_7 ? 8'h59 : _GEN_4000; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4002 = 8'ha2 == io_state_in_7 ? 8'h5f : _GEN_4001; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4003 = 8'ha3 == io_state_in_7 ? 8'h5d : _GEN_4002; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4004 = 8'ha4 == io_state_in_7 ? 8'h53 : _GEN_4003; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4005 = 8'ha5 == io_state_in_7 ? 8'h51 : _GEN_4004; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4006 = 8'ha6 == io_state_in_7 ? 8'h57 : _GEN_4005; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4007 = 8'ha7 == io_state_in_7 ? 8'h55 : _GEN_4006; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4008 = 8'ha8 == io_state_in_7 ? 8'h4b : _GEN_4007; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4009 = 8'ha9 == io_state_in_7 ? 8'h49 : _GEN_4008; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4010 = 8'haa == io_state_in_7 ? 8'h4f : _GEN_4009; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4011 = 8'hab == io_state_in_7 ? 8'h4d : _GEN_4010; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4012 = 8'hac == io_state_in_7 ? 8'h43 : _GEN_4011; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4013 = 8'had == io_state_in_7 ? 8'h41 : _GEN_4012; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4014 = 8'hae == io_state_in_7 ? 8'h47 : _GEN_4013; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4015 = 8'haf == io_state_in_7 ? 8'h45 : _GEN_4014; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4016 = 8'hb0 == io_state_in_7 ? 8'h7b : _GEN_4015; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4017 = 8'hb1 == io_state_in_7 ? 8'h79 : _GEN_4016; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4018 = 8'hb2 == io_state_in_7 ? 8'h7f : _GEN_4017; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4019 = 8'hb3 == io_state_in_7 ? 8'h7d : _GEN_4018; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4020 = 8'hb4 == io_state_in_7 ? 8'h73 : _GEN_4019; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4021 = 8'hb5 == io_state_in_7 ? 8'h71 : _GEN_4020; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4022 = 8'hb6 == io_state_in_7 ? 8'h77 : _GEN_4021; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4023 = 8'hb7 == io_state_in_7 ? 8'h75 : _GEN_4022; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4024 = 8'hb8 == io_state_in_7 ? 8'h6b : _GEN_4023; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4025 = 8'hb9 == io_state_in_7 ? 8'h69 : _GEN_4024; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4026 = 8'hba == io_state_in_7 ? 8'h6f : _GEN_4025; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4027 = 8'hbb == io_state_in_7 ? 8'h6d : _GEN_4026; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4028 = 8'hbc == io_state_in_7 ? 8'h63 : _GEN_4027; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4029 = 8'hbd == io_state_in_7 ? 8'h61 : _GEN_4028; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4030 = 8'hbe == io_state_in_7 ? 8'h67 : _GEN_4029; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4031 = 8'hbf == io_state_in_7 ? 8'h65 : _GEN_4030; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4032 = 8'hc0 == io_state_in_7 ? 8'h9b : _GEN_4031; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4033 = 8'hc1 == io_state_in_7 ? 8'h99 : _GEN_4032; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4034 = 8'hc2 == io_state_in_7 ? 8'h9f : _GEN_4033; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4035 = 8'hc3 == io_state_in_7 ? 8'h9d : _GEN_4034; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4036 = 8'hc4 == io_state_in_7 ? 8'h93 : _GEN_4035; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4037 = 8'hc5 == io_state_in_7 ? 8'h91 : _GEN_4036; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4038 = 8'hc6 == io_state_in_7 ? 8'h97 : _GEN_4037; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4039 = 8'hc7 == io_state_in_7 ? 8'h95 : _GEN_4038; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4040 = 8'hc8 == io_state_in_7 ? 8'h8b : _GEN_4039; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4041 = 8'hc9 == io_state_in_7 ? 8'h89 : _GEN_4040; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4042 = 8'hca == io_state_in_7 ? 8'h8f : _GEN_4041; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4043 = 8'hcb == io_state_in_7 ? 8'h8d : _GEN_4042; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4044 = 8'hcc == io_state_in_7 ? 8'h83 : _GEN_4043; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4045 = 8'hcd == io_state_in_7 ? 8'h81 : _GEN_4044; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4046 = 8'hce == io_state_in_7 ? 8'h87 : _GEN_4045; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4047 = 8'hcf == io_state_in_7 ? 8'h85 : _GEN_4046; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4048 = 8'hd0 == io_state_in_7 ? 8'hbb : _GEN_4047; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4049 = 8'hd1 == io_state_in_7 ? 8'hb9 : _GEN_4048; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4050 = 8'hd2 == io_state_in_7 ? 8'hbf : _GEN_4049; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4051 = 8'hd3 == io_state_in_7 ? 8'hbd : _GEN_4050; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4052 = 8'hd4 == io_state_in_7 ? 8'hb3 : _GEN_4051; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4053 = 8'hd5 == io_state_in_7 ? 8'hb1 : _GEN_4052; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4054 = 8'hd6 == io_state_in_7 ? 8'hb7 : _GEN_4053; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4055 = 8'hd7 == io_state_in_7 ? 8'hb5 : _GEN_4054; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4056 = 8'hd8 == io_state_in_7 ? 8'hab : _GEN_4055; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4057 = 8'hd9 == io_state_in_7 ? 8'ha9 : _GEN_4056; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4058 = 8'hda == io_state_in_7 ? 8'haf : _GEN_4057; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4059 = 8'hdb == io_state_in_7 ? 8'had : _GEN_4058; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4060 = 8'hdc == io_state_in_7 ? 8'ha3 : _GEN_4059; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4061 = 8'hdd == io_state_in_7 ? 8'ha1 : _GEN_4060; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4062 = 8'hde == io_state_in_7 ? 8'ha7 : _GEN_4061; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4063 = 8'hdf == io_state_in_7 ? 8'ha5 : _GEN_4062; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4064 = 8'he0 == io_state_in_7 ? 8'hdb : _GEN_4063; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4065 = 8'he1 == io_state_in_7 ? 8'hd9 : _GEN_4064; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4066 = 8'he2 == io_state_in_7 ? 8'hdf : _GEN_4065; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4067 = 8'he3 == io_state_in_7 ? 8'hdd : _GEN_4066; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4068 = 8'he4 == io_state_in_7 ? 8'hd3 : _GEN_4067; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4069 = 8'he5 == io_state_in_7 ? 8'hd1 : _GEN_4068; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4070 = 8'he6 == io_state_in_7 ? 8'hd7 : _GEN_4069; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4071 = 8'he7 == io_state_in_7 ? 8'hd5 : _GEN_4070; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4072 = 8'he8 == io_state_in_7 ? 8'hcb : _GEN_4071; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4073 = 8'he9 == io_state_in_7 ? 8'hc9 : _GEN_4072; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4074 = 8'hea == io_state_in_7 ? 8'hcf : _GEN_4073; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4075 = 8'heb == io_state_in_7 ? 8'hcd : _GEN_4074; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4076 = 8'hec == io_state_in_7 ? 8'hc3 : _GEN_4075; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4077 = 8'hed == io_state_in_7 ? 8'hc1 : _GEN_4076; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4078 = 8'hee == io_state_in_7 ? 8'hc7 : _GEN_4077; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4079 = 8'hef == io_state_in_7 ? 8'hc5 : _GEN_4078; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4080 = 8'hf0 == io_state_in_7 ? 8'hfb : _GEN_4079; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4081 = 8'hf1 == io_state_in_7 ? 8'hf9 : _GEN_4080; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4082 = 8'hf2 == io_state_in_7 ? 8'hff : _GEN_4081; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4083 = 8'hf3 == io_state_in_7 ? 8'hfd : _GEN_4082; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4084 = 8'hf4 == io_state_in_7 ? 8'hf3 : _GEN_4083; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4085 = 8'hf5 == io_state_in_7 ? 8'hf1 : _GEN_4084; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4086 = 8'hf6 == io_state_in_7 ? 8'hf7 : _GEN_4085; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4087 = 8'hf7 == io_state_in_7 ? 8'hf5 : _GEN_4086; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4088 = 8'hf8 == io_state_in_7 ? 8'heb : _GEN_4087; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4089 = 8'hf9 == io_state_in_7 ? 8'he9 : _GEN_4088; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4090 = 8'hfa == io_state_in_7 ? 8'hef : _GEN_4089; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4091 = 8'hfb == io_state_in_7 ? 8'hed : _GEN_4090; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4092 = 8'hfc == io_state_in_7 ? 8'he3 : _GEN_4091; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4093 = 8'hfd == io_state_in_7 ? 8'he1 : _GEN_4092; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4094 = 8'hfe == io_state_in_7 ? 8'he7 : _GEN_4093; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4095 = 8'hff == io_state_in_7 ? 8'he5 : _GEN_4094; // @[MixColumns.scala 133:{75,75}]
  wire [7:0] _GEN_4097 = 8'h1 == io_state_in_8 ? 8'h2 : 8'h0; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4098 = 8'h2 == io_state_in_8 ? 8'h4 : _GEN_4097; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4099 = 8'h3 == io_state_in_8 ? 8'h6 : _GEN_4098; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4100 = 8'h4 == io_state_in_8 ? 8'h8 : _GEN_4099; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4101 = 8'h5 == io_state_in_8 ? 8'ha : _GEN_4100; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4102 = 8'h6 == io_state_in_8 ? 8'hc : _GEN_4101; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4103 = 8'h7 == io_state_in_8 ? 8'he : _GEN_4102; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4104 = 8'h8 == io_state_in_8 ? 8'h10 : _GEN_4103; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4105 = 8'h9 == io_state_in_8 ? 8'h12 : _GEN_4104; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4106 = 8'ha == io_state_in_8 ? 8'h14 : _GEN_4105; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4107 = 8'hb == io_state_in_8 ? 8'h16 : _GEN_4106; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4108 = 8'hc == io_state_in_8 ? 8'h18 : _GEN_4107; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4109 = 8'hd == io_state_in_8 ? 8'h1a : _GEN_4108; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4110 = 8'he == io_state_in_8 ? 8'h1c : _GEN_4109; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4111 = 8'hf == io_state_in_8 ? 8'h1e : _GEN_4110; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4112 = 8'h10 == io_state_in_8 ? 8'h20 : _GEN_4111; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4113 = 8'h11 == io_state_in_8 ? 8'h22 : _GEN_4112; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4114 = 8'h12 == io_state_in_8 ? 8'h24 : _GEN_4113; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4115 = 8'h13 == io_state_in_8 ? 8'h26 : _GEN_4114; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4116 = 8'h14 == io_state_in_8 ? 8'h28 : _GEN_4115; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4117 = 8'h15 == io_state_in_8 ? 8'h2a : _GEN_4116; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4118 = 8'h16 == io_state_in_8 ? 8'h2c : _GEN_4117; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4119 = 8'h17 == io_state_in_8 ? 8'h2e : _GEN_4118; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4120 = 8'h18 == io_state_in_8 ? 8'h30 : _GEN_4119; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4121 = 8'h19 == io_state_in_8 ? 8'h32 : _GEN_4120; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4122 = 8'h1a == io_state_in_8 ? 8'h34 : _GEN_4121; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4123 = 8'h1b == io_state_in_8 ? 8'h36 : _GEN_4122; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4124 = 8'h1c == io_state_in_8 ? 8'h38 : _GEN_4123; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4125 = 8'h1d == io_state_in_8 ? 8'h3a : _GEN_4124; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4126 = 8'h1e == io_state_in_8 ? 8'h3c : _GEN_4125; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4127 = 8'h1f == io_state_in_8 ? 8'h3e : _GEN_4126; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4128 = 8'h20 == io_state_in_8 ? 8'h40 : _GEN_4127; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4129 = 8'h21 == io_state_in_8 ? 8'h42 : _GEN_4128; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4130 = 8'h22 == io_state_in_8 ? 8'h44 : _GEN_4129; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4131 = 8'h23 == io_state_in_8 ? 8'h46 : _GEN_4130; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4132 = 8'h24 == io_state_in_8 ? 8'h48 : _GEN_4131; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4133 = 8'h25 == io_state_in_8 ? 8'h4a : _GEN_4132; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4134 = 8'h26 == io_state_in_8 ? 8'h4c : _GEN_4133; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4135 = 8'h27 == io_state_in_8 ? 8'h4e : _GEN_4134; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4136 = 8'h28 == io_state_in_8 ? 8'h50 : _GEN_4135; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4137 = 8'h29 == io_state_in_8 ? 8'h52 : _GEN_4136; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4138 = 8'h2a == io_state_in_8 ? 8'h54 : _GEN_4137; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4139 = 8'h2b == io_state_in_8 ? 8'h56 : _GEN_4138; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4140 = 8'h2c == io_state_in_8 ? 8'h58 : _GEN_4139; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4141 = 8'h2d == io_state_in_8 ? 8'h5a : _GEN_4140; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4142 = 8'h2e == io_state_in_8 ? 8'h5c : _GEN_4141; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4143 = 8'h2f == io_state_in_8 ? 8'h5e : _GEN_4142; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4144 = 8'h30 == io_state_in_8 ? 8'h60 : _GEN_4143; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4145 = 8'h31 == io_state_in_8 ? 8'h62 : _GEN_4144; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4146 = 8'h32 == io_state_in_8 ? 8'h64 : _GEN_4145; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4147 = 8'h33 == io_state_in_8 ? 8'h66 : _GEN_4146; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4148 = 8'h34 == io_state_in_8 ? 8'h68 : _GEN_4147; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4149 = 8'h35 == io_state_in_8 ? 8'h6a : _GEN_4148; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4150 = 8'h36 == io_state_in_8 ? 8'h6c : _GEN_4149; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4151 = 8'h37 == io_state_in_8 ? 8'h6e : _GEN_4150; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4152 = 8'h38 == io_state_in_8 ? 8'h70 : _GEN_4151; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4153 = 8'h39 == io_state_in_8 ? 8'h72 : _GEN_4152; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4154 = 8'h3a == io_state_in_8 ? 8'h74 : _GEN_4153; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4155 = 8'h3b == io_state_in_8 ? 8'h76 : _GEN_4154; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4156 = 8'h3c == io_state_in_8 ? 8'h78 : _GEN_4155; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4157 = 8'h3d == io_state_in_8 ? 8'h7a : _GEN_4156; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4158 = 8'h3e == io_state_in_8 ? 8'h7c : _GEN_4157; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4159 = 8'h3f == io_state_in_8 ? 8'h7e : _GEN_4158; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4160 = 8'h40 == io_state_in_8 ? 8'h80 : _GEN_4159; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4161 = 8'h41 == io_state_in_8 ? 8'h82 : _GEN_4160; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4162 = 8'h42 == io_state_in_8 ? 8'h84 : _GEN_4161; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4163 = 8'h43 == io_state_in_8 ? 8'h86 : _GEN_4162; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4164 = 8'h44 == io_state_in_8 ? 8'h88 : _GEN_4163; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4165 = 8'h45 == io_state_in_8 ? 8'h8a : _GEN_4164; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4166 = 8'h46 == io_state_in_8 ? 8'h8c : _GEN_4165; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4167 = 8'h47 == io_state_in_8 ? 8'h8e : _GEN_4166; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4168 = 8'h48 == io_state_in_8 ? 8'h90 : _GEN_4167; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4169 = 8'h49 == io_state_in_8 ? 8'h92 : _GEN_4168; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4170 = 8'h4a == io_state_in_8 ? 8'h94 : _GEN_4169; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4171 = 8'h4b == io_state_in_8 ? 8'h96 : _GEN_4170; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4172 = 8'h4c == io_state_in_8 ? 8'h98 : _GEN_4171; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4173 = 8'h4d == io_state_in_8 ? 8'h9a : _GEN_4172; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4174 = 8'h4e == io_state_in_8 ? 8'h9c : _GEN_4173; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4175 = 8'h4f == io_state_in_8 ? 8'h9e : _GEN_4174; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4176 = 8'h50 == io_state_in_8 ? 8'ha0 : _GEN_4175; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4177 = 8'h51 == io_state_in_8 ? 8'ha2 : _GEN_4176; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4178 = 8'h52 == io_state_in_8 ? 8'ha4 : _GEN_4177; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4179 = 8'h53 == io_state_in_8 ? 8'ha6 : _GEN_4178; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4180 = 8'h54 == io_state_in_8 ? 8'ha8 : _GEN_4179; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4181 = 8'h55 == io_state_in_8 ? 8'haa : _GEN_4180; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4182 = 8'h56 == io_state_in_8 ? 8'hac : _GEN_4181; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4183 = 8'h57 == io_state_in_8 ? 8'hae : _GEN_4182; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4184 = 8'h58 == io_state_in_8 ? 8'hb0 : _GEN_4183; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4185 = 8'h59 == io_state_in_8 ? 8'hb2 : _GEN_4184; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4186 = 8'h5a == io_state_in_8 ? 8'hb4 : _GEN_4185; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4187 = 8'h5b == io_state_in_8 ? 8'hb6 : _GEN_4186; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4188 = 8'h5c == io_state_in_8 ? 8'hb8 : _GEN_4187; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4189 = 8'h5d == io_state_in_8 ? 8'hba : _GEN_4188; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4190 = 8'h5e == io_state_in_8 ? 8'hbc : _GEN_4189; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4191 = 8'h5f == io_state_in_8 ? 8'hbe : _GEN_4190; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4192 = 8'h60 == io_state_in_8 ? 8'hc0 : _GEN_4191; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4193 = 8'h61 == io_state_in_8 ? 8'hc2 : _GEN_4192; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4194 = 8'h62 == io_state_in_8 ? 8'hc4 : _GEN_4193; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4195 = 8'h63 == io_state_in_8 ? 8'hc6 : _GEN_4194; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4196 = 8'h64 == io_state_in_8 ? 8'hc8 : _GEN_4195; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4197 = 8'h65 == io_state_in_8 ? 8'hca : _GEN_4196; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4198 = 8'h66 == io_state_in_8 ? 8'hcc : _GEN_4197; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4199 = 8'h67 == io_state_in_8 ? 8'hce : _GEN_4198; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4200 = 8'h68 == io_state_in_8 ? 8'hd0 : _GEN_4199; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4201 = 8'h69 == io_state_in_8 ? 8'hd2 : _GEN_4200; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4202 = 8'h6a == io_state_in_8 ? 8'hd4 : _GEN_4201; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4203 = 8'h6b == io_state_in_8 ? 8'hd6 : _GEN_4202; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4204 = 8'h6c == io_state_in_8 ? 8'hd8 : _GEN_4203; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4205 = 8'h6d == io_state_in_8 ? 8'hda : _GEN_4204; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4206 = 8'h6e == io_state_in_8 ? 8'hdc : _GEN_4205; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4207 = 8'h6f == io_state_in_8 ? 8'hde : _GEN_4206; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4208 = 8'h70 == io_state_in_8 ? 8'he0 : _GEN_4207; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4209 = 8'h71 == io_state_in_8 ? 8'he2 : _GEN_4208; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4210 = 8'h72 == io_state_in_8 ? 8'he4 : _GEN_4209; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4211 = 8'h73 == io_state_in_8 ? 8'he6 : _GEN_4210; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4212 = 8'h74 == io_state_in_8 ? 8'he8 : _GEN_4211; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4213 = 8'h75 == io_state_in_8 ? 8'hea : _GEN_4212; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4214 = 8'h76 == io_state_in_8 ? 8'hec : _GEN_4213; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4215 = 8'h77 == io_state_in_8 ? 8'hee : _GEN_4214; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4216 = 8'h78 == io_state_in_8 ? 8'hf0 : _GEN_4215; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4217 = 8'h79 == io_state_in_8 ? 8'hf2 : _GEN_4216; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4218 = 8'h7a == io_state_in_8 ? 8'hf4 : _GEN_4217; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4219 = 8'h7b == io_state_in_8 ? 8'hf6 : _GEN_4218; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4220 = 8'h7c == io_state_in_8 ? 8'hf8 : _GEN_4219; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4221 = 8'h7d == io_state_in_8 ? 8'hfa : _GEN_4220; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4222 = 8'h7e == io_state_in_8 ? 8'hfc : _GEN_4221; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4223 = 8'h7f == io_state_in_8 ? 8'hfe : _GEN_4222; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4224 = 8'h80 == io_state_in_8 ? 8'h1b : _GEN_4223; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4225 = 8'h81 == io_state_in_8 ? 8'h19 : _GEN_4224; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4226 = 8'h82 == io_state_in_8 ? 8'h1f : _GEN_4225; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4227 = 8'h83 == io_state_in_8 ? 8'h1d : _GEN_4226; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4228 = 8'h84 == io_state_in_8 ? 8'h13 : _GEN_4227; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4229 = 8'h85 == io_state_in_8 ? 8'h11 : _GEN_4228; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4230 = 8'h86 == io_state_in_8 ? 8'h17 : _GEN_4229; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4231 = 8'h87 == io_state_in_8 ? 8'h15 : _GEN_4230; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4232 = 8'h88 == io_state_in_8 ? 8'hb : _GEN_4231; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4233 = 8'h89 == io_state_in_8 ? 8'h9 : _GEN_4232; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4234 = 8'h8a == io_state_in_8 ? 8'hf : _GEN_4233; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4235 = 8'h8b == io_state_in_8 ? 8'hd : _GEN_4234; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4236 = 8'h8c == io_state_in_8 ? 8'h3 : _GEN_4235; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4237 = 8'h8d == io_state_in_8 ? 8'h1 : _GEN_4236; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4238 = 8'h8e == io_state_in_8 ? 8'h7 : _GEN_4237; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4239 = 8'h8f == io_state_in_8 ? 8'h5 : _GEN_4238; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4240 = 8'h90 == io_state_in_8 ? 8'h3b : _GEN_4239; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4241 = 8'h91 == io_state_in_8 ? 8'h39 : _GEN_4240; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4242 = 8'h92 == io_state_in_8 ? 8'h3f : _GEN_4241; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4243 = 8'h93 == io_state_in_8 ? 8'h3d : _GEN_4242; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4244 = 8'h94 == io_state_in_8 ? 8'h33 : _GEN_4243; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4245 = 8'h95 == io_state_in_8 ? 8'h31 : _GEN_4244; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4246 = 8'h96 == io_state_in_8 ? 8'h37 : _GEN_4245; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4247 = 8'h97 == io_state_in_8 ? 8'h35 : _GEN_4246; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4248 = 8'h98 == io_state_in_8 ? 8'h2b : _GEN_4247; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4249 = 8'h99 == io_state_in_8 ? 8'h29 : _GEN_4248; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4250 = 8'h9a == io_state_in_8 ? 8'h2f : _GEN_4249; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4251 = 8'h9b == io_state_in_8 ? 8'h2d : _GEN_4250; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4252 = 8'h9c == io_state_in_8 ? 8'h23 : _GEN_4251; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4253 = 8'h9d == io_state_in_8 ? 8'h21 : _GEN_4252; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4254 = 8'h9e == io_state_in_8 ? 8'h27 : _GEN_4253; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4255 = 8'h9f == io_state_in_8 ? 8'h25 : _GEN_4254; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4256 = 8'ha0 == io_state_in_8 ? 8'h5b : _GEN_4255; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4257 = 8'ha1 == io_state_in_8 ? 8'h59 : _GEN_4256; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4258 = 8'ha2 == io_state_in_8 ? 8'h5f : _GEN_4257; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4259 = 8'ha3 == io_state_in_8 ? 8'h5d : _GEN_4258; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4260 = 8'ha4 == io_state_in_8 ? 8'h53 : _GEN_4259; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4261 = 8'ha5 == io_state_in_8 ? 8'h51 : _GEN_4260; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4262 = 8'ha6 == io_state_in_8 ? 8'h57 : _GEN_4261; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4263 = 8'ha7 == io_state_in_8 ? 8'h55 : _GEN_4262; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4264 = 8'ha8 == io_state_in_8 ? 8'h4b : _GEN_4263; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4265 = 8'ha9 == io_state_in_8 ? 8'h49 : _GEN_4264; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4266 = 8'haa == io_state_in_8 ? 8'h4f : _GEN_4265; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4267 = 8'hab == io_state_in_8 ? 8'h4d : _GEN_4266; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4268 = 8'hac == io_state_in_8 ? 8'h43 : _GEN_4267; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4269 = 8'had == io_state_in_8 ? 8'h41 : _GEN_4268; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4270 = 8'hae == io_state_in_8 ? 8'h47 : _GEN_4269; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4271 = 8'haf == io_state_in_8 ? 8'h45 : _GEN_4270; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4272 = 8'hb0 == io_state_in_8 ? 8'h7b : _GEN_4271; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4273 = 8'hb1 == io_state_in_8 ? 8'h79 : _GEN_4272; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4274 = 8'hb2 == io_state_in_8 ? 8'h7f : _GEN_4273; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4275 = 8'hb3 == io_state_in_8 ? 8'h7d : _GEN_4274; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4276 = 8'hb4 == io_state_in_8 ? 8'h73 : _GEN_4275; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4277 = 8'hb5 == io_state_in_8 ? 8'h71 : _GEN_4276; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4278 = 8'hb6 == io_state_in_8 ? 8'h77 : _GEN_4277; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4279 = 8'hb7 == io_state_in_8 ? 8'h75 : _GEN_4278; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4280 = 8'hb8 == io_state_in_8 ? 8'h6b : _GEN_4279; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4281 = 8'hb9 == io_state_in_8 ? 8'h69 : _GEN_4280; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4282 = 8'hba == io_state_in_8 ? 8'h6f : _GEN_4281; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4283 = 8'hbb == io_state_in_8 ? 8'h6d : _GEN_4282; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4284 = 8'hbc == io_state_in_8 ? 8'h63 : _GEN_4283; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4285 = 8'hbd == io_state_in_8 ? 8'h61 : _GEN_4284; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4286 = 8'hbe == io_state_in_8 ? 8'h67 : _GEN_4285; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4287 = 8'hbf == io_state_in_8 ? 8'h65 : _GEN_4286; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4288 = 8'hc0 == io_state_in_8 ? 8'h9b : _GEN_4287; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4289 = 8'hc1 == io_state_in_8 ? 8'h99 : _GEN_4288; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4290 = 8'hc2 == io_state_in_8 ? 8'h9f : _GEN_4289; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4291 = 8'hc3 == io_state_in_8 ? 8'h9d : _GEN_4290; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4292 = 8'hc4 == io_state_in_8 ? 8'h93 : _GEN_4291; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4293 = 8'hc5 == io_state_in_8 ? 8'h91 : _GEN_4292; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4294 = 8'hc6 == io_state_in_8 ? 8'h97 : _GEN_4293; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4295 = 8'hc7 == io_state_in_8 ? 8'h95 : _GEN_4294; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4296 = 8'hc8 == io_state_in_8 ? 8'h8b : _GEN_4295; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4297 = 8'hc9 == io_state_in_8 ? 8'h89 : _GEN_4296; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4298 = 8'hca == io_state_in_8 ? 8'h8f : _GEN_4297; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4299 = 8'hcb == io_state_in_8 ? 8'h8d : _GEN_4298; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4300 = 8'hcc == io_state_in_8 ? 8'h83 : _GEN_4299; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4301 = 8'hcd == io_state_in_8 ? 8'h81 : _GEN_4300; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4302 = 8'hce == io_state_in_8 ? 8'h87 : _GEN_4301; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4303 = 8'hcf == io_state_in_8 ? 8'h85 : _GEN_4302; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4304 = 8'hd0 == io_state_in_8 ? 8'hbb : _GEN_4303; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4305 = 8'hd1 == io_state_in_8 ? 8'hb9 : _GEN_4304; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4306 = 8'hd2 == io_state_in_8 ? 8'hbf : _GEN_4305; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4307 = 8'hd3 == io_state_in_8 ? 8'hbd : _GEN_4306; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4308 = 8'hd4 == io_state_in_8 ? 8'hb3 : _GEN_4307; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4309 = 8'hd5 == io_state_in_8 ? 8'hb1 : _GEN_4308; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4310 = 8'hd6 == io_state_in_8 ? 8'hb7 : _GEN_4309; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4311 = 8'hd7 == io_state_in_8 ? 8'hb5 : _GEN_4310; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4312 = 8'hd8 == io_state_in_8 ? 8'hab : _GEN_4311; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4313 = 8'hd9 == io_state_in_8 ? 8'ha9 : _GEN_4312; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4314 = 8'hda == io_state_in_8 ? 8'haf : _GEN_4313; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4315 = 8'hdb == io_state_in_8 ? 8'had : _GEN_4314; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4316 = 8'hdc == io_state_in_8 ? 8'ha3 : _GEN_4315; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4317 = 8'hdd == io_state_in_8 ? 8'ha1 : _GEN_4316; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4318 = 8'hde == io_state_in_8 ? 8'ha7 : _GEN_4317; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4319 = 8'hdf == io_state_in_8 ? 8'ha5 : _GEN_4318; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4320 = 8'he0 == io_state_in_8 ? 8'hdb : _GEN_4319; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4321 = 8'he1 == io_state_in_8 ? 8'hd9 : _GEN_4320; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4322 = 8'he2 == io_state_in_8 ? 8'hdf : _GEN_4321; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4323 = 8'he3 == io_state_in_8 ? 8'hdd : _GEN_4322; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4324 = 8'he4 == io_state_in_8 ? 8'hd3 : _GEN_4323; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4325 = 8'he5 == io_state_in_8 ? 8'hd1 : _GEN_4324; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4326 = 8'he6 == io_state_in_8 ? 8'hd7 : _GEN_4325; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4327 = 8'he7 == io_state_in_8 ? 8'hd5 : _GEN_4326; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4328 = 8'he8 == io_state_in_8 ? 8'hcb : _GEN_4327; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4329 = 8'he9 == io_state_in_8 ? 8'hc9 : _GEN_4328; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4330 = 8'hea == io_state_in_8 ? 8'hcf : _GEN_4329; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4331 = 8'heb == io_state_in_8 ? 8'hcd : _GEN_4330; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4332 = 8'hec == io_state_in_8 ? 8'hc3 : _GEN_4331; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4333 = 8'hed == io_state_in_8 ? 8'hc1 : _GEN_4332; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4334 = 8'hee == io_state_in_8 ? 8'hc7 : _GEN_4333; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4335 = 8'hef == io_state_in_8 ? 8'hc5 : _GEN_4334; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4336 = 8'hf0 == io_state_in_8 ? 8'hfb : _GEN_4335; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4337 = 8'hf1 == io_state_in_8 ? 8'hf9 : _GEN_4336; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4338 = 8'hf2 == io_state_in_8 ? 8'hff : _GEN_4337; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4339 = 8'hf3 == io_state_in_8 ? 8'hfd : _GEN_4338; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4340 = 8'hf4 == io_state_in_8 ? 8'hf3 : _GEN_4339; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4341 = 8'hf5 == io_state_in_8 ? 8'hf1 : _GEN_4340; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4342 = 8'hf6 == io_state_in_8 ? 8'hf7 : _GEN_4341; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4343 = 8'hf7 == io_state_in_8 ? 8'hf5 : _GEN_4342; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4344 = 8'hf8 == io_state_in_8 ? 8'heb : _GEN_4343; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4345 = 8'hf9 == io_state_in_8 ? 8'he9 : _GEN_4344; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4346 = 8'hfa == io_state_in_8 ? 8'hef : _GEN_4345; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4347 = 8'hfb == io_state_in_8 ? 8'hed : _GEN_4346; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4348 = 8'hfc == io_state_in_8 ? 8'he3 : _GEN_4347; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4349 = 8'hfd == io_state_in_8 ? 8'he1 : _GEN_4348; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4350 = 8'hfe == io_state_in_8 ? 8'he7 : _GEN_4349; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4351 = 8'hff == io_state_in_8 ? 8'he5 : _GEN_4350; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4353 = 8'h1 == io_state_in_9 ? 8'h3 : 8'h0; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4354 = 8'h2 == io_state_in_9 ? 8'h6 : _GEN_4353; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4355 = 8'h3 == io_state_in_9 ? 8'h5 : _GEN_4354; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4356 = 8'h4 == io_state_in_9 ? 8'hc : _GEN_4355; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4357 = 8'h5 == io_state_in_9 ? 8'hf : _GEN_4356; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4358 = 8'h6 == io_state_in_9 ? 8'ha : _GEN_4357; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4359 = 8'h7 == io_state_in_9 ? 8'h9 : _GEN_4358; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4360 = 8'h8 == io_state_in_9 ? 8'h18 : _GEN_4359; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4361 = 8'h9 == io_state_in_9 ? 8'h1b : _GEN_4360; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4362 = 8'ha == io_state_in_9 ? 8'h1e : _GEN_4361; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4363 = 8'hb == io_state_in_9 ? 8'h1d : _GEN_4362; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4364 = 8'hc == io_state_in_9 ? 8'h14 : _GEN_4363; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4365 = 8'hd == io_state_in_9 ? 8'h17 : _GEN_4364; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4366 = 8'he == io_state_in_9 ? 8'h12 : _GEN_4365; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4367 = 8'hf == io_state_in_9 ? 8'h11 : _GEN_4366; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4368 = 8'h10 == io_state_in_9 ? 8'h30 : _GEN_4367; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4369 = 8'h11 == io_state_in_9 ? 8'h33 : _GEN_4368; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4370 = 8'h12 == io_state_in_9 ? 8'h36 : _GEN_4369; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4371 = 8'h13 == io_state_in_9 ? 8'h35 : _GEN_4370; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4372 = 8'h14 == io_state_in_9 ? 8'h3c : _GEN_4371; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4373 = 8'h15 == io_state_in_9 ? 8'h3f : _GEN_4372; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4374 = 8'h16 == io_state_in_9 ? 8'h3a : _GEN_4373; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4375 = 8'h17 == io_state_in_9 ? 8'h39 : _GEN_4374; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4376 = 8'h18 == io_state_in_9 ? 8'h28 : _GEN_4375; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4377 = 8'h19 == io_state_in_9 ? 8'h2b : _GEN_4376; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4378 = 8'h1a == io_state_in_9 ? 8'h2e : _GEN_4377; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4379 = 8'h1b == io_state_in_9 ? 8'h2d : _GEN_4378; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4380 = 8'h1c == io_state_in_9 ? 8'h24 : _GEN_4379; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4381 = 8'h1d == io_state_in_9 ? 8'h27 : _GEN_4380; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4382 = 8'h1e == io_state_in_9 ? 8'h22 : _GEN_4381; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4383 = 8'h1f == io_state_in_9 ? 8'h21 : _GEN_4382; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4384 = 8'h20 == io_state_in_9 ? 8'h60 : _GEN_4383; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4385 = 8'h21 == io_state_in_9 ? 8'h63 : _GEN_4384; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4386 = 8'h22 == io_state_in_9 ? 8'h66 : _GEN_4385; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4387 = 8'h23 == io_state_in_9 ? 8'h65 : _GEN_4386; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4388 = 8'h24 == io_state_in_9 ? 8'h6c : _GEN_4387; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4389 = 8'h25 == io_state_in_9 ? 8'h6f : _GEN_4388; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4390 = 8'h26 == io_state_in_9 ? 8'h6a : _GEN_4389; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4391 = 8'h27 == io_state_in_9 ? 8'h69 : _GEN_4390; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4392 = 8'h28 == io_state_in_9 ? 8'h78 : _GEN_4391; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4393 = 8'h29 == io_state_in_9 ? 8'h7b : _GEN_4392; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4394 = 8'h2a == io_state_in_9 ? 8'h7e : _GEN_4393; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4395 = 8'h2b == io_state_in_9 ? 8'h7d : _GEN_4394; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4396 = 8'h2c == io_state_in_9 ? 8'h74 : _GEN_4395; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4397 = 8'h2d == io_state_in_9 ? 8'h77 : _GEN_4396; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4398 = 8'h2e == io_state_in_9 ? 8'h72 : _GEN_4397; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4399 = 8'h2f == io_state_in_9 ? 8'h71 : _GEN_4398; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4400 = 8'h30 == io_state_in_9 ? 8'h50 : _GEN_4399; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4401 = 8'h31 == io_state_in_9 ? 8'h53 : _GEN_4400; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4402 = 8'h32 == io_state_in_9 ? 8'h56 : _GEN_4401; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4403 = 8'h33 == io_state_in_9 ? 8'h55 : _GEN_4402; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4404 = 8'h34 == io_state_in_9 ? 8'h5c : _GEN_4403; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4405 = 8'h35 == io_state_in_9 ? 8'h5f : _GEN_4404; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4406 = 8'h36 == io_state_in_9 ? 8'h5a : _GEN_4405; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4407 = 8'h37 == io_state_in_9 ? 8'h59 : _GEN_4406; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4408 = 8'h38 == io_state_in_9 ? 8'h48 : _GEN_4407; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4409 = 8'h39 == io_state_in_9 ? 8'h4b : _GEN_4408; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4410 = 8'h3a == io_state_in_9 ? 8'h4e : _GEN_4409; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4411 = 8'h3b == io_state_in_9 ? 8'h4d : _GEN_4410; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4412 = 8'h3c == io_state_in_9 ? 8'h44 : _GEN_4411; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4413 = 8'h3d == io_state_in_9 ? 8'h47 : _GEN_4412; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4414 = 8'h3e == io_state_in_9 ? 8'h42 : _GEN_4413; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4415 = 8'h3f == io_state_in_9 ? 8'h41 : _GEN_4414; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4416 = 8'h40 == io_state_in_9 ? 8'hc0 : _GEN_4415; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4417 = 8'h41 == io_state_in_9 ? 8'hc3 : _GEN_4416; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4418 = 8'h42 == io_state_in_9 ? 8'hc6 : _GEN_4417; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4419 = 8'h43 == io_state_in_9 ? 8'hc5 : _GEN_4418; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4420 = 8'h44 == io_state_in_9 ? 8'hcc : _GEN_4419; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4421 = 8'h45 == io_state_in_9 ? 8'hcf : _GEN_4420; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4422 = 8'h46 == io_state_in_9 ? 8'hca : _GEN_4421; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4423 = 8'h47 == io_state_in_9 ? 8'hc9 : _GEN_4422; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4424 = 8'h48 == io_state_in_9 ? 8'hd8 : _GEN_4423; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4425 = 8'h49 == io_state_in_9 ? 8'hdb : _GEN_4424; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4426 = 8'h4a == io_state_in_9 ? 8'hde : _GEN_4425; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4427 = 8'h4b == io_state_in_9 ? 8'hdd : _GEN_4426; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4428 = 8'h4c == io_state_in_9 ? 8'hd4 : _GEN_4427; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4429 = 8'h4d == io_state_in_9 ? 8'hd7 : _GEN_4428; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4430 = 8'h4e == io_state_in_9 ? 8'hd2 : _GEN_4429; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4431 = 8'h4f == io_state_in_9 ? 8'hd1 : _GEN_4430; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4432 = 8'h50 == io_state_in_9 ? 8'hf0 : _GEN_4431; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4433 = 8'h51 == io_state_in_9 ? 8'hf3 : _GEN_4432; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4434 = 8'h52 == io_state_in_9 ? 8'hf6 : _GEN_4433; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4435 = 8'h53 == io_state_in_9 ? 8'hf5 : _GEN_4434; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4436 = 8'h54 == io_state_in_9 ? 8'hfc : _GEN_4435; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4437 = 8'h55 == io_state_in_9 ? 8'hff : _GEN_4436; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4438 = 8'h56 == io_state_in_9 ? 8'hfa : _GEN_4437; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4439 = 8'h57 == io_state_in_9 ? 8'hf9 : _GEN_4438; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4440 = 8'h58 == io_state_in_9 ? 8'he8 : _GEN_4439; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4441 = 8'h59 == io_state_in_9 ? 8'heb : _GEN_4440; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4442 = 8'h5a == io_state_in_9 ? 8'hee : _GEN_4441; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4443 = 8'h5b == io_state_in_9 ? 8'hed : _GEN_4442; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4444 = 8'h5c == io_state_in_9 ? 8'he4 : _GEN_4443; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4445 = 8'h5d == io_state_in_9 ? 8'he7 : _GEN_4444; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4446 = 8'h5e == io_state_in_9 ? 8'he2 : _GEN_4445; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4447 = 8'h5f == io_state_in_9 ? 8'he1 : _GEN_4446; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4448 = 8'h60 == io_state_in_9 ? 8'ha0 : _GEN_4447; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4449 = 8'h61 == io_state_in_9 ? 8'ha3 : _GEN_4448; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4450 = 8'h62 == io_state_in_9 ? 8'ha6 : _GEN_4449; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4451 = 8'h63 == io_state_in_9 ? 8'ha5 : _GEN_4450; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4452 = 8'h64 == io_state_in_9 ? 8'hac : _GEN_4451; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4453 = 8'h65 == io_state_in_9 ? 8'haf : _GEN_4452; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4454 = 8'h66 == io_state_in_9 ? 8'haa : _GEN_4453; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4455 = 8'h67 == io_state_in_9 ? 8'ha9 : _GEN_4454; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4456 = 8'h68 == io_state_in_9 ? 8'hb8 : _GEN_4455; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4457 = 8'h69 == io_state_in_9 ? 8'hbb : _GEN_4456; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4458 = 8'h6a == io_state_in_9 ? 8'hbe : _GEN_4457; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4459 = 8'h6b == io_state_in_9 ? 8'hbd : _GEN_4458; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4460 = 8'h6c == io_state_in_9 ? 8'hb4 : _GEN_4459; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4461 = 8'h6d == io_state_in_9 ? 8'hb7 : _GEN_4460; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4462 = 8'h6e == io_state_in_9 ? 8'hb2 : _GEN_4461; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4463 = 8'h6f == io_state_in_9 ? 8'hb1 : _GEN_4462; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4464 = 8'h70 == io_state_in_9 ? 8'h90 : _GEN_4463; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4465 = 8'h71 == io_state_in_9 ? 8'h93 : _GEN_4464; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4466 = 8'h72 == io_state_in_9 ? 8'h96 : _GEN_4465; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4467 = 8'h73 == io_state_in_9 ? 8'h95 : _GEN_4466; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4468 = 8'h74 == io_state_in_9 ? 8'h9c : _GEN_4467; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4469 = 8'h75 == io_state_in_9 ? 8'h9f : _GEN_4468; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4470 = 8'h76 == io_state_in_9 ? 8'h9a : _GEN_4469; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4471 = 8'h77 == io_state_in_9 ? 8'h99 : _GEN_4470; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4472 = 8'h78 == io_state_in_9 ? 8'h88 : _GEN_4471; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4473 = 8'h79 == io_state_in_9 ? 8'h8b : _GEN_4472; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4474 = 8'h7a == io_state_in_9 ? 8'h8e : _GEN_4473; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4475 = 8'h7b == io_state_in_9 ? 8'h8d : _GEN_4474; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4476 = 8'h7c == io_state_in_9 ? 8'h84 : _GEN_4475; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4477 = 8'h7d == io_state_in_9 ? 8'h87 : _GEN_4476; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4478 = 8'h7e == io_state_in_9 ? 8'h82 : _GEN_4477; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4479 = 8'h7f == io_state_in_9 ? 8'h81 : _GEN_4478; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4480 = 8'h80 == io_state_in_9 ? 8'h9b : _GEN_4479; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4481 = 8'h81 == io_state_in_9 ? 8'h98 : _GEN_4480; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4482 = 8'h82 == io_state_in_9 ? 8'h9d : _GEN_4481; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4483 = 8'h83 == io_state_in_9 ? 8'h9e : _GEN_4482; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4484 = 8'h84 == io_state_in_9 ? 8'h97 : _GEN_4483; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4485 = 8'h85 == io_state_in_9 ? 8'h94 : _GEN_4484; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4486 = 8'h86 == io_state_in_9 ? 8'h91 : _GEN_4485; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4487 = 8'h87 == io_state_in_9 ? 8'h92 : _GEN_4486; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4488 = 8'h88 == io_state_in_9 ? 8'h83 : _GEN_4487; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4489 = 8'h89 == io_state_in_9 ? 8'h80 : _GEN_4488; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4490 = 8'h8a == io_state_in_9 ? 8'h85 : _GEN_4489; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4491 = 8'h8b == io_state_in_9 ? 8'h86 : _GEN_4490; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4492 = 8'h8c == io_state_in_9 ? 8'h8f : _GEN_4491; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4493 = 8'h8d == io_state_in_9 ? 8'h8c : _GEN_4492; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4494 = 8'h8e == io_state_in_9 ? 8'h89 : _GEN_4493; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4495 = 8'h8f == io_state_in_9 ? 8'h8a : _GEN_4494; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4496 = 8'h90 == io_state_in_9 ? 8'hab : _GEN_4495; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4497 = 8'h91 == io_state_in_9 ? 8'ha8 : _GEN_4496; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4498 = 8'h92 == io_state_in_9 ? 8'had : _GEN_4497; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4499 = 8'h93 == io_state_in_9 ? 8'hae : _GEN_4498; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4500 = 8'h94 == io_state_in_9 ? 8'ha7 : _GEN_4499; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4501 = 8'h95 == io_state_in_9 ? 8'ha4 : _GEN_4500; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4502 = 8'h96 == io_state_in_9 ? 8'ha1 : _GEN_4501; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4503 = 8'h97 == io_state_in_9 ? 8'ha2 : _GEN_4502; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4504 = 8'h98 == io_state_in_9 ? 8'hb3 : _GEN_4503; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4505 = 8'h99 == io_state_in_9 ? 8'hb0 : _GEN_4504; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4506 = 8'h9a == io_state_in_9 ? 8'hb5 : _GEN_4505; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4507 = 8'h9b == io_state_in_9 ? 8'hb6 : _GEN_4506; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4508 = 8'h9c == io_state_in_9 ? 8'hbf : _GEN_4507; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4509 = 8'h9d == io_state_in_9 ? 8'hbc : _GEN_4508; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4510 = 8'h9e == io_state_in_9 ? 8'hb9 : _GEN_4509; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4511 = 8'h9f == io_state_in_9 ? 8'hba : _GEN_4510; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4512 = 8'ha0 == io_state_in_9 ? 8'hfb : _GEN_4511; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4513 = 8'ha1 == io_state_in_9 ? 8'hf8 : _GEN_4512; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4514 = 8'ha2 == io_state_in_9 ? 8'hfd : _GEN_4513; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4515 = 8'ha3 == io_state_in_9 ? 8'hfe : _GEN_4514; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4516 = 8'ha4 == io_state_in_9 ? 8'hf7 : _GEN_4515; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4517 = 8'ha5 == io_state_in_9 ? 8'hf4 : _GEN_4516; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4518 = 8'ha6 == io_state_in_9 ? 8'hf1 : _GEN_4517; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4519 = 8'ha7 == io_state_in_9 ? 8'hf2 : _GEN_4518; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4520 = 8'ha8 == io_state_in_9 ? 8'he3 : _GEN_4519; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4521 = 8'ha9 == io_state_in_9 ? 8'he0 : _GEN_4520; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4522 = 8'haa == io_state_in_9 ? 8'he5 : _GEN_4521; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4523 = 8'hab == io_state_in_9 ? 8'he6 : _GEN_4522; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4524 = 8'hac == io_state_in_9 ? 8'hef : _GEN_4523; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4525 = 8'had == io_state_in_9 ? 8'hec : _GEN_4524; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4526 = 8'hae == io_state_in_9 ? 8'he9 : _GEN_4525; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4527 = 8'haf == io_state_in_9 ? 8'hea : _GEN_4526; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4528 = 8'hb0 == io_state_in_9 ? 8'hcb : _GEN_4527; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4529 = 8'hb1 == io_state_in_9 ? 8'hc8 : _GEN_4528; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4530 = 8'hb2 == io_state_in_9 ? 8'hcd : _GEN_4529; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4531 = 8'hb3 == io_state_in_9 ? 8'hce : _GEN_4530; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4532 = 8'hb4 == io_state_in_9 ? 8'hc7 : _GEN_4531; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4533 = 8'hb5 == io_state_in_9 ? 8'hc4 : _GEN_4532; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4534 = 8'hb6 == io_state_in_9 ? 8'hc1 : _GEN_4533; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4535 = 8'hb7 == io_state_in_9 ? 8'hc2 : _GEN_4534; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4536 = 8'hb8 == io_state_in_9 ? 8'hd3 : _GEN_4535; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4537 = 8'hb9 == io_state_in_9 ? 8'hd0 : _GEN_4536; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4538 = 8'hba == io_state_in_9 ? 8'hd5 : _GEN_4537; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4539 = 8'hbb == io_state_in_9 ? 8'hd6 : _GEN_4538; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4540 = 8'hbc == io_state_in_9 ? 8'hdf : _GEN_4539; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4541 = 8'hbd == io_state_in_9 ? 8'hdc : _GEN_4540; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4542 = 8'hbe == io_state_in_9 ? 8'hd9 : _GEN_4541; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4543 = 8'hbf == io_state_in_9 ? 8'hda : _GEN_4542; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4544 = 8'hc0 == io_state_in_9 ? 8'h5b : _GEN_4543; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4545 = 8'hc1 == io_state_in_9 ? 8'h58 : _GEN_4544; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4546 = 8'hc2 == io_state_in_9 ? 8'h5d : _GEN_4545; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4547 = 8'hc3 == io_state_in_9 ? 8'h5e : _GEN_4546; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4548 = 8'hc4 == io_state_in_9 ? 8'h57 : _GEN_4547; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4549 = 8'hc5 == io_state_in_9 ? 8'h54 : _GEN_4548; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4550 = 8'hc6 == io_state_in_9 ? 8'h51 : _GEN_4549; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4551 = 8'hc7 == io_state_in_9 ? 8'h52 : _GEN_4550; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4552 = 8'hc8 == io_state_in_9 ? 8'h43 : _GEN_4551; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4553 = 8'hc9 == io_state_in_9 ? 8'h40 : _GEN_4552; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4554 = 8'hca == io_state_in_9 ? 8'h45 : _GEN_4553; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4555 = 8'hcb == io_state_in_9 ? 8'h46 : _GEN_4554; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4556 = 8'hcc == io_state_in_9 ? 8'h4f : _GEN_4555; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4557 = 8'hcd == io_state_in_9 ? 8'h4c : _GEN_4556; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4558 = 8'hce == io_state_in_9 ? 8'h49 : _GEN_4557; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4559 = 8'hcf == io_state_in_9 ? 8'h4a : _GEN_4558; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4560 = 8'hd0 == io_state_in_9 ? 8'h6b : _GEN_4559; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4561 = 8'hd1 == io_state_in_9 ? 8'h68 : _GEN_4560; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4562 = 8'hd2 == io_state_in_9 ? 8'h6d : _GEN_4561; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4563 = 8'hd3 == io_state_in_9 ? 8'h6e : _GEN_4562; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4564 = 8'hd4 == io_state_in_9 ? 8'h67 : _GEN_4563; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4565 = 8'hd5 == io_state_in_9 ? 8'h64 : _GEN_4564; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4566 = 8'hd6 == io_state_in_9 ? 8'h61 : _GEN_4565; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4567 = 8'hd7 == io_state_in_9 ? 8'h62 : _GEN_4566; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4568 = 8'hd8 == io_state_in_9 ? 8'h73 : _GEN_4567; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4569 = 8'hd9 == io_state_in_9 ? 8'h70 : _GEN_4568; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4570 = 8'hda == io_state_in_9 ? 8'h75 : _GEN_4569; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4571 = 8'hdb == io_state_in_9 ? 8'h76 : _GEN_4570; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4572 = 8'hdc == io_state_in_9 ? 8'h7f : _GEN_4571; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4573 = 8'hdd == io_state_in_9 ? 8'h7c : _GEN_4572; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4574 = 8'hde == io_state_in_9 ? 8'h79 : _GEN_4573; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4575 = 8'hdf == io_state_in_9 ? 8'h7a : _GEN_4574; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4576 = 8'he0 == io_state_in_9 ? 8'h3b : _GEN_4575; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4577 = 8'he1 == io_state_in_9 ? 8'h38 : _GEN_4576; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4578 = 8'he2 == io_state_in_9 ? 8'h3d : _GEN_4577; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4579 = 8'he3 == io_state_in_9 ? 8'h3e : _GEN_4578; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4580 = 8'he4 == io_state_in_9 ? 8'h37 : _GEN_4579; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4581 = 8'he5 == io_state_in_9 ? 8'h34 : _GEN_4580; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4582 = 8'he6 == io_state_in_9 ? 8'h31 : _GEN_4581; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4583 = 8'he7 == io_state_in_9 ? 8'h32 : _GEN_4582; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4584 = 8'he8 == io_state_in_9 ? 8'h23 : _GEN_4583; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4585 = 8'he9 == io_state_in_9 ? 8'h20 : _GEN_4584; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4586 = 8'hea == io_state_in_9 ? 8'h25 : _GEN_4585; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4587 = 8'heb == io_state_in_9 ? 8'h26 : _GEN_4586; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4588 = 8'hec == io_state_in_9 ? 8'h2f : _GEN_4587; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4589 = 8'hed == io_state_in_9 ? 8'h2c : _GEN_4588; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4590 = 8'hee == io_state_in_9 ? 8'h29 : _GEN_4589; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4591 = 8'hef == io_state_in_9 ? 8'h2a : _GEN_4590; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4592 = 8'hf0 == io_state_in_9 ? 8'hb : _GEN_4591; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4593 = 8'hf1 == io_state_in_9 ? 8'h8 : _GEN_4592; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4594 = 8'hf2 == io_state_in_9 ? 8'hd : _GEN_4593; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4595 = 8'hf3 == io_state_in_9 ? 8'he : _GEN_4594; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4596 = 8'hf4 == io_state_in_9 ? 8'h7 : _GEN_4595; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4597 = 8'hf5 == io_state_in_9 ? 8'h4 : _GEN_4596; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4598 = 8'hf6 == io_state_in_9 ? 8'h1 : _GEN_4597; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4599 = 8'hf7 == io_state_in_9 ? 8'h2 : _GEN_4598; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4600 = 8'hf8 == io_state_in_9 ? 8'h13 : _GEN_4599; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4601 = 8'hf9 == io_state_in_9 ? 8'h10 : _GEN_4600; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4602 = 8'hfa == io_state_in_9 ? 8'h15 : _GEN_4601; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4603 = 8'hfb == io_state_in_9 ? 8'h16 : _GEN_4602; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4604 = 8'hfc == io_state_in_9 ? 8'h1f : _GEN_4603; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4605 = 8'hfd == io_state_in_9 ? 8'h1c : _GEN_4604; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4606 = 8'hfe == io_state_in_9 ? 8'h19 : _GEN_4605; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _GEN_4607 = 8'hff == io_state_in_9 ? 8'h1a : _GEN_4606; // @[MixColumns.scala 135:{41,41}]
  wire [7:0] _tmp_state_8_T = _GEN_4351 ^ _GEN_4607; // @[MixColumns.scala 135:41]
  wire [7:0] _tmp_state_8_T_1 = _tmp_state_8_T ^ io_state_in_10; // @[MixColumns.scala 135:65]
  wire [7:0] _GEN_4609 = 8'h1 == io_state_in_9 ? 8'h2 : 8'h0; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4610 = 8'h2 == io_state_in_9 ? 8'h4 : _GEN_4609; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4611 = 8'h3 == io_state_in_9 ? 8'h6 : _GEN_4610; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4612 = 8'h4 == io_state_in_9 ? 8'h8 : _GEN_4611; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4613 = 8'h5 == io_state_in_9 ? 8'ha : _GEN_4612; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4614 = 8'h6 == io_state_in_9 ? 8'hc : _GEN_4613; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4615 = 8'h7 == io_state_in_9 ? 8'he : _GEN_4614; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4616 = 8'h8 == io_state_in_9 ? 8'h10 : _GEN_4615; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4617 = 8'h9 == io_state_in_9 ? 8'h12 : _GEN_4616; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4618 = 8'ha == io_state_in_9 ? 8'h14 : _GEN_4617; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4619 = 8'hb == io_state_in_9 ? 8'h16 : _GEN_4618; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4620 = 8'hc == io_state_in_9 ? 8'h18 : _GEN_4619; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4621 = 8'hd == io_state_in_9 ? 8'h1a : _GEN_4620; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4622 = 8'he == io_state_in_9 ? 8'h1c : _GEN_4621; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4623 = 8'hf == io_state_in_9 ? 8'h1e : _GEN_4622; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4624 = 8'h10 == io_state_in_9 ? 8'h20 : _GEN_4623; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4625 = 8'h11 == io_state_in_9 ? 8'h22 : _GEN_4624; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4626 = 8'h12 == io_state_in_9 ? 8'h24 : _GEN_4625; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4627 = 8'h13 == io_state_in_9 ? 8'h26 : _GEN_4626; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4628 = 8'h14 == io_state_in_9 ? 8'h28 : _GEN_4627; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4629 = 8'h15 == io_state_in_9 ? 8'h2a : _GEN_4628; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4630 = 8'h16 == io_state_in_9 ? 8'h2c : _GEN_4629; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4631 = 8'h17 == io_state_in_9 ? 8'h2e : _GEN_4630; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4632 = 8'h18 == io_state_in_9 ? 8'h30 : _GEN_4631; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4633 = 8'h19 == io_state_in_9 ? 8'h32 : _GEN_4632; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4634 = 8'h1a == io_state_in_9 ? 8'h34 : _GEN_4633; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4635 = 8'h1b == io_state_in_9 ? 8'h36 : _GEN_4634; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4636 = 8'h1c == io_state_in_9 ? 8'h38 : _GEN_4635; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4637 = 8'h1d == io_state_in_9 ? 8'h3a : _GEN_4636; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4638 = 8'h1e == io_state_in_9 ? 8'h3c : _GEN_4637; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4639 = 8'h1f == io_state_in_9 ? 8'h3e : _GEN_4638; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4640 = 8'h20 == io_state_in_9 ? 8'h40 : _GEN_4639; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4641 = 8'h21 == io_state_in_9 ? 8'h42 : _GEN_4640; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4642 = 8'h22 == io_state_in_9 ? 8'h44 : _GEN_4641; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4643 = 8'h23 == io_state_in_9 ? 8'h46 : _GEN_4642; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4644 = 8'h24 == io_state_in_9 ? 8'h48 : _GEN_4643; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4645 = 8'h25 == io_state_in_9 ? 8'h4a : _GEN_4644; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4646 = 8'h26 == io_state_in_9 ? 8'h4c : _GEN_4645; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4647 = 8'h27 == io_state_in_9 ? 8'h4e : _GEN_4646; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4648 = 8'h28 == io_state_in_9 ? 8'h50 : _GEN_4647; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4649 = 8'h29 == io_state_in_9 ? 8'h52 : _GEN_4648; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4650 = 8'h2a == io_state_in_9 ? 8'h54 : _GEN_4649; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4651 = 8'h2b == io_state_in_9 ? 8'h56 : _GEN_4650; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4652 = 8'h2c == io_state_in_9 ? 8'h58 : _GEN_4651; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4653 = 8'h2d == io_state_in_9 ? 8'h5a : _GEN_4652; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4654 = 8'h2e == io_state_in_9 ? 8'h5c : _GEN_4653; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4655 = 8'h2f == io_state_in_9 ? 8'h5e : _GEN_4654; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4656 = 8'h30 == io_state_in_9 ? 8'h60 : _GEN_4655; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4657 = 8'h31 == io_state_in_9 ? 8'h62 : _GEN_4656; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4658 = 8'h32 == io_state_in_9 ? 8'h64 : _GEN_4657; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4659 = 8'h33 == io_state_in_9 ? 8'h66 : _GEN_4658; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4660 = 8'h34 == io_state_in_9 ? 8'h68 : _GEN_4659; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4661 = 8'h35 == io_state_in_9 ? 8'h6a : _GEN_4660; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4662 = 8'h36 == io_state_in_9 ? 8'h6c : _GEN_4661; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4663 = 8'h37 == io_state_in_9 ? 8'h6e : _GEN_4662; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4664 = 8'h38 == io_state_in_9 ? 8'h70 : _GEN_4663; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4665 = 8'h39 == io_state_in_9 ? 8'h72 : _GEN_4664; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4666 = 8'h3a == io_state_in_9 ? 8'h74 : _GEN_4665; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4667 = 8'h3b == io_state_in_9 ? 8'h76 : _GEN_4666; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4668 = 8'h3c == io_state_in_9 ? 8'h78 : _GEN_4667; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4669 = 8'h3d == io_state_in_9 ? 8'h7a : _GEN_4668; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4670 = 8'h3e == io_state_in_9 ? 8'h7c : _GEN_4669; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4671 = 8'h3f == io_state_in_9 ? 8'h7e : _GEN_4670; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4672 = 8'h40 == io_state_in_9 ? 8'h80 : _GEN_4671; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4673 = 8'h41 == io_state_in_9 ? 8'h82 : _GEN_4672; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4674 = 8'h42 == io_state_in_9 ? 8'h84 : _GEN_4673; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4675 = 8'h43 == io_state_in_9 ? 8'h86 : _GEN_4674; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4676 = 8'h44 == io_state_in_9 ? 8'h88 : _GEN_4675; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4677 = 8'h45 == io_state_in_9 ? 8'h8a : _GEN_4676; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4678 = 8'h46 == io_state_in_9 ? 8'h8c : _GEN_4677; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4679 = 8'h47 == io_state_in_9 ? 8'h8e : _GEN_4678; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4680 = 8'h48 == io_state_in_9 ? 8'h90 : _GEN_4679; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4681 = 8'h49 == io_state_in_9 ? 8'h92 : _GEN_4680; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4682 = 8'h4a == io_state_in_9 ? 8'h94 : _GEN_4681; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4683 = 8'h4b == io_state_in_9 ? 8'h96 : _GEN_4682; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4684 = 8'h4c == io_state_in_9 ? 8'h98 : _GEN_4683; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4685 = 8'h4d == io_state_in_9 ? 8'h9a : _GEN_4684; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4686 = 8'h4e == io_state_in_9 ? 8'h9c : _GEN_4685; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4687 = 8'h4f == io_state_in_9 ? 8'h9e : _GEN_4686; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4688 = 8'h50 == io_state_in_9 ? 8'ha0 : _GEN_4687; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4689 = 8'h51 == io_state_in_9 ? 8'ha2 : _GEN_4688; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4690 = 8'h52 == io_state_in_9 ? 8'ha4 : _GEN_4689; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4691 = 8'h53 == io_state_in_9 ? 8'ha6 : _GEN_4690; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4692 = 8'h54 == io_state_in_9 ? 8'ha8 : _GEN_4691; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4693 = 8'h55 == io_state_in_9 ? 8'haa : _GEN_4692; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4694 = 8'h56 == io_state_in_9 ? 8'hac : _GEN_4693; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4695 = 8'h57 == io_state_in_9 ? 8'hae : _GEN_4694; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4696 = 8'h58 == io_state_in_9 ? 8'hb0 : _GEN_4695; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4697 = 8'h59 == io_state_in_9 ? 8'hb2 : _GEN_4696; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4698 = 8'h5a == io_state_in_9 ? 8'hb4 : _GEN_4697; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4699 = 8'h5b == io_state_in_9 ? 8'hb6 : _GEN_4698; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4700 = 8'h5c == io_state_in_9 ? 8'hb8 : _GEN_4699; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4701 = 8'h5d == io_state_in_9 ? 8'hba : _GEN_4700; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4702 = 8'h5e == io_state_in_9 ? 8'hbc : _GEN_4701; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4703 = 8'h5f == io_state_in_9 ? 8'hbe : _GEN_4702; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4704 = 8'h60 == io_state_in_9 ? 8'hc0 : _GEN_4703; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4705 = 8'h61 == io_state_in_9 ? 8'hc2 : _GEN_4704; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4706 = 8'h62 == io_state_in_9 ? 8'hc4 : _GEN_4705; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4707 = 8'h63 == io_state_in_9 ? 8'hc6 : _GEN_4706; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4708 = 8'h64 == io_state_in_9 ? 8'hc8 : _GEN_4707; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4709 = 8'h65 == io_state_in_9 ? 8'hca : _GEN_4708; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4710 = 8'h66 == io_state_in_9 ? 8'hcc : _GEN_4709; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4711 = 8'h67 == io_state_in_9 ? 8'hce : _GEN_4710; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4712 = 8'h68 == io_state_in_9 ? 8'hd0 : _GEN_4711; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4713 = 8'h69 == io_state_in_9 ? 8'hd2 : _GEN_4712; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4714 = 8'h6a == io_state_in_9 ? 8'hd4 : _GEN_4713; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4715 = 8'h6b == io_state_in_9 ? 8'hd6 : _GEN_4714; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4716 = 8'h6c == io_state_in_9 ? 8'hd8 : _GEN_4715; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4717 = 8'h6d == io_state_in_9 ? 8'hda : _GEN_4716; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4718 = 8'h6e == io_state_in_9 ? 8'hdc : _GEN_4717; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4719 = 8'h6f == io_state_in_9 ? 8'hde : _GEN_4718; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4720 = 8'h70 == io_state_in_9 ? 8'he0 : _GEN_4719; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4721 = 8'h71 == io_state_in_9 ? 8'he2 : _GEN_4720; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4722 = 8'h72 == io_state_in_9 ? 8'he4 : _GEN_4721; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4723 = 8'h73 == io_state_in_9 ? 8'he6 : _GEN_4722; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4724 = 8'h74 == io_state_in_9 ? 8'he8 : _GEN_4723; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4725 = 8'h75 == io_state_in_9 ? 8'hea : _GEN_4724; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4726 = 8'h76 == io_state_in_9 ? 8'hec : _GEN_4725; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4727 = 8'h77 == io_state_in_9 ? 8'hee : _GEN_4726; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4728 = 8'h78 == io_state_in_9 ? 8'hf0 : _GEN_4727; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4729 = 8'h79 == io_state_in_9 ? 8'hf2 : _GEN_4728; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4730 = 8'h7a == io_state_in_9 ? 8'hf4 : _GEN_4729; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4731 = 8'h7b == io_state_in_9 ? 8'hf6 : _GEN_4730; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4732 = 8'h7c == io_state_in_9 ? 8'hf8 : _GEN_4731; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4733 = 8'h7d == io_state_in_9 ? 8'hfa : _GEN_4732; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4734 = 8'h7e == io_state_in_9 ? 8'hfc : _GEN_4733; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4735 = 8'h7f == io_state_in_9 ? 8'hfe : _GEN_4734; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4736 = 8'h80 == io_state_in_9 ? 8'h1b : _GEN_4735; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4737 = 8'h81 == io_state_in_9 ? 8'h19 : _GEN_4736; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4738 = 8'h82 == io_state_in_9 ? 8'h1f : _GEN_4737; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4739 = 8'h83 == io_state_in_9 ? 8'h1d : _GEN_4738; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4740 = 8'h84 == io_state_in_9 ? 8'h13 : _GEN_4739; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4741 = 8'h85 == io_state_in_9 ? 8'h11 : _GEN_4740; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4742 = 8'h86 == io_state_in_9 ? 8'h17 : _GEN_4741; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4743 = 8'h87 == io_state_in_9 ? 8'h15 : _GEN_4742; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4744 = 8'h88 == io_state_in_9 ? 8'hb : _GEN_4743; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4745 = 8'h89 == io_state_in_9 ? 8'h9 : _GEN_4744; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4746 = 8'h8a == io_state_in_9 ? 8'hf : _GEN_4745; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4747 = 8'h8b == io_state_in_9 ? 8'hd : _GEN_4746; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4748 = 8'h8c == io_state_in_9 ? 8'h3 : _GEN_4747; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4749 = 8'h8d == io_state_in_9 ? 8'h1 : _GEN_4748; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4750 = 8'h8e == io_state_in_9 ? 8'h7 : _GEN_4749; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4751 = 8'h8f == io_state_in_9 ? 8'h5 : _GEN_4750; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4752 = 8'h90 == io_state_in_9 ? 8'h3b : _GEN_4751; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4753 = 8'h91 == io_state_in_9 ? 8'h39 : _GEN_4752; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4754 = 8'h92 == io_state_in_9 ? 8'h3f : _GEN_4753; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4755 = 8'h93 == io_state_in_9 ? 8'h3d : _GEN_4754; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4756 = 8'h94 == io_state_in_9 ? 8'h33 : _GEN_4755; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4757 = 8'h95 == io_state_in_9 ? 8'h31 : _GEN_4756; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4758 = 8'h96 == io_state_in_9 ? 8'h37 : _GEN_4757; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4759 = 8'h97 == io_state_in_9 ? 8'h35 : _GEN_4758; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4760 = 8'h98 == io_state_in_9 ? 8'h2b : _GEN_4759; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4761 = 8'h99 == io_state_in_9 ? 8'h29 : _GEN_4760; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4762 = 8'h9a == io_state_in_9 ? 8'h2f : _GEN_4761; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4763 = 8'h9b == io_state_in_9 ? 8'h2d : _GEN_4762; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4764 = 8'h9c == io_state_in_9 ? 8'h23 : _GEN_4763; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4765 = 8'h9d == io_state_in_9 ? 8'h21 : _GEN_4764; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4766 = 8'h9e == io_state_in_9 ? 8'h27 : _GEN_4765; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4767 = 8'h9f == io_state_in_9 ? 8'h25 : _GEN_4766; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4768 = 8'ha0 == io_state_in_9 ? 8'h5b : _GEN_4767; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4769 = 8'ha1 == io_state_in_9 ? 8'h59 : _GEN_4768; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4770 = 8'ha2 == io_state_in_9 ? 8'h5f : _GEN_4769; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4771 = 8'ha3 == io_state_in_9 ? 8'h5d : _GEN_4770; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4772 = 8'ha4 == io_state_in_9 ? 8'h53 : _GEN_4771; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4773 = 8'ha5 == io_state_in_9 ? 8'h51 : _GEN_4772; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4774 = 8'ha6 == io_state_in_9 ? 8'h57 : _GEN_4773; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4775 = 8'ha7 == io_state_in_9 ? 8'h55 : _GEN_4774; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4776 = 8'ha8 == io_state_in_9 ? 8'h4b : _GEN_4775; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4777 = 8'ha9 == io_state_in_9 ? 8'h49 : _GEN_4776; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4778 = 8'haa == io_state_in_9 ? 8'h4f : _GEN_4777; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4779 = 8'hab == io_state_in_9 ? 8'h4d : _GEN_4778; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4780 = 8'hac == io_state_in_9 ? 8'h43 : _GEN_4779; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4781 = 8'had == io_state_in_9 ? 8'h41 : _GEN_4780; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4782 = 8'hae == io_state_in_9 ? 8'h47 : _GEN_4781; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4783 = 8'haf == io_state_in_9 ? 8'h45 : _GEN_4782; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4784 = 8'hb0 == io_state_in_9 ? 8'h7b : _GEN_4783; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4785 = 8'hb1 == io_state_in_9 ? 8'h79 : _GEN_4784; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4786 = 8'hb2 == io_state_in_9 ? 8'h7f : _GEN_4785; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4787 = 8'hb3 == io_state_in_9 ? 8'h7d : _GEN_4786; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4788 = 8'hb4 == io_state_in_9 ? 8'h73 : _GEN_4787; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4789 = 8'hb5 == io_state_in_9 ? 8'h71 : _GEN_4788; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4790 = 8'hb6 == io_state_in_9 ? 8'h77 : _GEN_4789; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4791 = 8'hb7 == io_state_in_9 ? 8'h75 : _GEN_4790; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4792 = 8'hb8 == io_state_in_9 ? 8'h6b : _GEN_4791; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4793 = 8'hb9 == io_state_in_9 ? 8'h69 : _GEN_4792; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4794 = 8'hba == io_state_in_9 ? 8'h6f : _GEN_4793; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4795 = 8'hbb == io_state_in_9 ? 8'h6d : _GEN_4794; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4796 = 8'hbc == io_state_in_9 ? 8'h63 : _GEN_4795; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4797 = 8'hbd == io_state_in_9 ? 8'h61 : _GEN_4796; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4798 = 8'hbe == io_state_in_9 ? 8'h67 : _GEN_4797; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4799 = 8'hbf == io_state_in_9 ? 8'h65 : _GEN_4798; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4800 = 8'hc0 == io_state_in_9 ? 8'h9b : _GEN_4799; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4801 = 8'hc1 == io_state_in_9 ? 8'h99 : _GEN_4800; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4802 = 8'hc2 == io_state_in_9 ? 8'h9f : _GEN_4801; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4803 = 8'hc3 == io_state_in_9 ? 8'h9d : _GEN_4802; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4804 = 8'hc4 == io_state_in_9 ? 8'h93 : _GEN_4803; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4805 = 8'hc5 == io_state_in_9 ? 8'h91 : _GEN_4804; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4806 = 8'hc6 == io_state_in_9 ? 8'h97 : _GEN_4805; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4807 = 8'hc7 == io_state_in_9 ? 8'h95 : _GEN_4806; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4808 = 8'hc8 == io_state_in_9 ? 8'h8b : _GEN_4807; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4809 = 8'hc9 == io_state_in_9 ? 8'h89 : _GEN_4808; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4810 = 8'hca == io_state_in_9 ? 8'h8f : _GEN_4809; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4811 = 8'hcb == io_state_in_9 ? 8'h8d : _GEN_4810; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4812 = 8'hcc == io_state_in_9 ? 8'h83 : _GEN_4811; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4813 = 8'hcd == io_state_in_9 ? 8'h81 : _GEN_4812; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4814 = 8'hce == io_state_in_9 ? 8'h87 : _GEN_4813; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4815 = 8'hcf == io_state_in_9 ? 8'h85 : _GEN_4814; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4816 = 8'hd0 == io_state_in_9 ? 8'hbb : _GEN_4815; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4817 = 8'hd1 == io_state_in_9 ? 8'hb9 : _GEN_4816; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4818 = 8'hd2 == io_state_in_9 ? 8'hbf : _GEN_4817; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4819 = 8'hd3 == io_state_in_9 ? 8'hbd : _GEN_4818; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4820 = 8'hd4 == io_state_in_9 ? 8'hb3 : _GEN_4819; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4821 = 8'hd5 == io_state_in_9 ? 8'hb1 : _GEN_4820; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4822 = 8'hd6 == io_state_in_9 ? 8'hb7 : _GEN_4821; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4823 = 8'hd7 == io_state_in_9 ? 8'hb5 : _GEN_4822; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4824 = 8'hd8 == io_state_in_9 ? 8'hab : _GEN_4823; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4825 = 8'hd9 == io_state_in_9 ? 8'ha9 : _GEN_4824; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4826 = 8'hda == io_state_in_9 ? 8'haf : _GEN_4825; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4827 = 8'hdb == io_state_in_9 ? 8'had : _GEN_4826; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4828 = 8'hdc == io_state_in_9 ? 8'ha3 : _GEN_4827; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4829 = 8'hdd == io_state_in_9 ? 8'ha1 : _GEN_4828; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4830 = 8'hde == io_state_in_9 ? 8'ha7 : _GEN_4829; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4831 = 8'hdf == io_state_in_9 ? 8'ha5 : _GEN_4830; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4832 = 8'he0 == io_state_in_9 ? 8'hdb : _GEN_4831; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4833 = 8'he1 == io_state_in_9 ? 8'hd9 : _GEN_4832; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4834 = 8'he2 == io_state_in_9 ? 8'hdf : _GEN_4833; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4835 = 8'he3 == io_state_in_9 ? 8'hdd : _GEN_4834; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4836 = 8'he4 == io_state_in_9 ? 8'hd3 : _GEN_4835; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4837 = 8'he5 == io_state_in_9 ? 8'hd1 : _GEN_4836; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4838 = 8'he6 == io_state_in_9 ? 8'hd7 : _GEN_4837; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4839 = 8'he7 == io_state_in_9 ? 8'hd5 : _GEN_4838; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4840 = 8'he8 == io_state_in_9 ? 8'hcb : _GEN_4839; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4841 = 8'he9 == io_state_in_9 ? 8'hc9 : _GEN_4840; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4842 = 8'hea == io_state_in_9 ? 8'hcf : _GEN_4841; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4843 = 8'heb == io_state_in_9 ? 8'hcd : _GEN_4842; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4844 = 8'hec == io_state_in_9 ? 8'hc3 : _GEN_4843; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4845 = 8'hed == io_state_in_9 ? 8'hc1 : _GEN_4844; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4846 = 8'hee == io_state_in_9 ? 8'hc7 : _GEN_4845; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4847 = 8'hef == io_state_in_9 ? 8'hc5 : _GEN_4846; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4848 = 8'hf0 == io_state_in_9 ? 8'hfb : _GEN_4847; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4849 = 8'hf1 == io_state_in_9 ? 8'hf9 : _GEN_4848; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4850 = 8'hf2 == io_state_in_9 ? 8'hff : _GEN_4849; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4851 = 8'hf3 == io_state_in_9 ? 8'hfd : _GEN_4850; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4852 = 8'hf4 == io_state_in_9 ? 8'hf3 : _GEN_4851; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4853 = 8'hf5 == io_state_in_9 ? 8'hf1 : _GEN_4852; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4854 = 8'hf6 == io_state_in_9 ? 8'hf7 : _GEN_4853; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4855 = 8'hf7 == io_state_in_9 ? 8'hf5 : _GEN_4854; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4856 = 8'hf8 == io_state_in_9 ? 8'heb : _GEN_4855; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4857 = 8'hf9 == io_state_in_9 ? 8'he9 : _GEN_4856; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4858 = 8'hfa == io_state_in_9 ? 8'hef : _GEN_4857; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4859 = 8'hfb == io_state_in_9 ? 8'hed : _GEN_4858; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4860 = 8'hfc == io_state_in_9 ? 8'he3 : _GEN_4859; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4861 = 8'hfd == io_state_in_9 ? 8'he1 : _GEN_4860; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4862 = 8'hfe == io_state_in_9 ? 8'he7 : _GEN_4861; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _GEN_4863 = 8'hff == io_state_in_9 ? 8'he5 : _GEN_4862; // @[MixColumns.scala 136:{34,34}]
  wire [7:0] _tmp_state_9_T = io_state_in_8 ^ _GEN_4863; // @[MixColumns.scala 136:34]
  wire [7:0] _GEN_4865 = 8'h1 == io_state_in_10 ? 8'h3 : 8'h0; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4866 = 8'h2 == io_state_in_10 ? 8'h6 : _GEN_4865; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4867 = 8'h3 == io_state_in_10 ? 8'h5 : _GEN_4866; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4868 = 8'h4 == io_state_in_10 ? 8'hc : _GEN_4867; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4869 = 8'h5 == io_state_in_10 ? 8'hf : _GEN_4868; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4870 = 8'h6 == io_state_in_10 ? 8'ha : _GEN_4869; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4871 = 8'h7 == io_state_in_10 ? 8'h9 : _GEN_4870; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4872 = 8'h8 == io_state_in_10 ? 8'h18 : _GEN_4871; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4873 = 8'h9 == io_state_in_10 ? 8'h1b : _GEN_4872; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4874 = 8'ha == io_state_in_10 ? 8'h1e : _GEN_4873; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4875 = 8'hb == io_state_in_10 ? 8'h1d : _GEN_4874; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4876 = 8'hc == io_state_in_10 ? 8'h14 : _GEN_4875; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4877 = 8'hd == io_state_in_10 ? 8'h17 : _GEN_4876; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4878 = 8'he == io_state_in_10 ? 8'h12 : _GEN_4877; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4879 = 8'hf == io_state_in_10 ? 8'h11 : _GEN_4878; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4880 = 8'h10 == io_state_in_10 ? 8'h30 : _GEN_4879; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4881 = 8'h11 == io_state_in_10 ? 8'h33 : _GEN_4880; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4882 = 8'h12 == io_state_in_10 ? 8'h36 : _GEN_4881; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4883 = 8'h13 == io_state_in_10 ? 8'h35 : _GEN_4882; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4884 = 8'h14 == io_state_in_10 ? 8'h3c : _GEN_4883; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4885 = 8'h15 == io_state_in_10 ? 8'h3f : _GEN_4884; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4886 = 8'h16 == io_state_in_10 ? 8'h3a : _GEN_4885; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4887 = 8'h17 == io_state_in_10 ? 8'h39 : _GEN_4886; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4888 = 8'h18 == io_state_in_10 ? 8'h28 : _GEN_4887; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4889 = 8'h19 == io_state_in_10 ? 8'h2b : _GEN_4888; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4890 = 8'h1a == io_state_in_10 ? 8'h2e : _GEN_4889; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4891 = 8'h1b == io_state_in_10 ? 8'h2d : _GEN_4890; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4892 = 8'h1c == io_state_in_10 ? 8'h24 : _GEN_4891; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4893 = 8'h1d == io_state_in_10 ? 8'h27 : _GEN_4892; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4894 = 8'h1e == io_state_in_10 ? 8'h22 : _GEN_4893; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4895 = 8'h1f == io_state_in_10 ? 8'h21 : _GEN_4894; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4896 = 8'h20 == io_state_in_10 ? 8'h60 : _GEN_4895; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4897 = 8'h21 == io_state_in_10 ? 8'h63 : _GEN_4896; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4898 = 8'h22 == io_state_in_10 ? 8'h66 : _GEN_4897; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4899 = 8'h23 == io_state_in_10 ? 8'h65 : _GEN_4898; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4900 = 8'h24 == io_state_in_10 ? 8'h6c : _GEN_4899; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4901 = 8'h25 == io_state_in_10 ? 8'h6f : _GEN_4900; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4902 = 8'h26 == io_state_in_10 ? 8'h6a : _GEN_4901; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4903 = 8'h27 == io_state_in_10 ? 8'h69 : _GEN_4902; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4904 = 8'h28 == io_state_in_10 ? 8'h78 : _GEN_4903; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4905 = 8'h29 == io_state_in_10 ? 8'h7b : _GEN_4904; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4906 = 8'h2a == io_state_in_10 ? 8'h7e : _GEN_4905; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4907 = 8'h2b == io_state_in_10 ? 8'h7d : _GEN_4906; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4908 = 8'h2c == io_state_in_10 ? 8'h74 : _GEN_4907; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4909 = 8'h2d == io_state_in_10 ? 8'h77 : _GEN_4908; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4910 = 8'h2e == io_state_in_10 ? 8'h72 : _GEN_4909; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4911 = 8'h2f == io_state_in_10 ? 8'h71 : _GEN_4910; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4912 = 8'h30 == io_state_in_10 ? 8'h50 : _GEN_4911; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4913 = 8'h31 == io_state_in_10 ? 8'h53 : _GEN_4912; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4914 = 8'h32 == io_state_in_10 ? 8'h56 : _GEN_4913; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4915 = 8'h33 == io_state_in_10 ? 8'h55 : _GEN_4914; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4916 = 8'h34 == io_state_in_10 ? 8'h5c : _GEN_4915; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4917 = 8'h35 == io_state_in_10 ? 8'h5f : _GEN_4916; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4918 = 8'h36 == io_state_in_10 ? 8'h5a : _GEN_4917; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4919 = 8'h37 == io_state_in_10 ? 8'h59 : _GEN_4918; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4920 = 8'h38 == io_state_in_10 ? 8'h48 : _GEN_4919; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4921 = 8'h39 == io_state_in_10 ? 8'h4b : _GEN_4920; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4922 = 8'h3a == io_state_in_10 ? 8'h4e : _GEN_4921; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4923 = 8'h3b == io_state_in_10 ? 8'h4d : _GEN_4922; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4924 = 8'h3c == io_state_in_10 ? 8'h44 : _GEN_4923; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4925 = 8'h3d == io_state_in_10 ? 8'h47 : _GEN_4924; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4926 = 8'h3e == io_state_in_10 ? 8'h42 : _GEN_4925; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4927 = 8'h3f == io_state_in_10 ? 8'h41 : _GEN_4926; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4928 = 8'h40 == io_state_in_10 ? 8'hc0 : _GEN_4927; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4929 = 8'h41 == io_state_in_10 ? 8'hc3 : _GEN_4928; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4930 = 8'h42 == io_state_in_10 ? 8'hc6 : _GEN_4929; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4931 = 8'h43 == io_state_in_10 ? 8'hc5 : _GEN_4930; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4932 = 8'h44 == io_state_in_10 ? 8'hcc : _GEN_4931; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4933 = 8'h45 == io_state_in_10 ? 8'hcf : _GEN_4932; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4934 = 8'h46 == io_state_in_10 ? 8'hca : _GEN_4933; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4935 = 8'h47 == io_state_in_10 ? 8'hc9 : _GEN_4934; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4936 = 8'h48 == io_state_in_10 ? 8'hd8 : _GEN_4935; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4937 = 8'h49 == io_state_in_10 ? 8'hdb : _GEN_4936; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4938 = 8'h4a == io_state_in_10 ? 8'hde : _GEN_4937; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4939 = 8'h4b == io_state_in_10 ? 8'hdd : _GEN_4938; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4940 = 8'h4c == io_state_in_10 ? 8'hd4 : _GEN_4939; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4941 = 8'h4d == io_state_in_10 ? 8'hd7 : _GEN_4940; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4942 = 8'h4e == io_state_in_10 ? 8'hd2 : _GEN_4941; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4943 = 8'h4f == io_state_in_10 ? 8'hd1 : _GEN_4942; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4944 = 8'h50 == io_state_in_10 ? 8'hf0 : _GEN_4943; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4945 = 8'h51 == io_state_in_10 ? 8'hf3 : _GEN_4944; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4946 = 8'h52 == io_state_in_10 ? 8'hf6 : _GEN_4945; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4947 = 8'h53 == io_state_in_10 ? 8'hf5 : _GEN_4946; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4948 = 8'h54 == io_state_in_10 ? 8'hfc : _GEN_4947; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4949 = 8'h55 == io_state_in_10 ? 8'hff : _GEN_4948; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4950 = 8'h56 == io_state_in_10 ? 8'hfa : _GEN_4949; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4951 = 8'h57 == io_state_in_10 ? 8'hf9 : _GEN_4950; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4952 = 8'h58 == io_state_in_10 ? 8'he8 : _GEN_4951; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4953 = 8'h59 == io_state_in_10 ? 8'heb : _GEN_4952; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4954 = 8'h5a == io_state_in_10 ? 8'hee : _GEN_4953; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4955 = 8'h5b == io_state_in_10 ? 8'hed : _GEN_4954; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4956 = 8'h5c == io_state_in_10 ? 8'he4 : _GEN_4955; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4957 = 8'h5d == io_state_in_10 ? 8'he7 : _GEN_4956; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4958 = 8'h5e == io_state_in_10 ? 8'he2 : _GEN_4957; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4959 = 8'h5f == io_state_in_10 ? 8'he1 : _GEN_4958; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4960 = 8'h60 == io_state_in_10 ? 8'ha0 : _GEN_4959; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4961 = 8'h61 == io_state_in_10 ? 8'ha3 : _GEN_4960; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4962 = 8'h62 == io_state_in_10 ? 8'ha6 : _GEN_4961; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4963 = 8'h63 == io_state_in_10 ? 8'ha5 : _GEN_4962; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4964 = 8'h64 == io_state_in_10 ? 8'hac : _GEN_4963; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4965 = 8'h65 == io_state_in_10 ? 8'haf : _GEN_4964; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4966 = 8'h66 == io_state_in_10 ? 8'haa : _GEN_4965; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4967 = 8'h67 == io_state_in_10 ? 8'ha9 : _GEN_4966; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4968 = 8'h68 == io_state_in_10 ? 8'hb8 : _GEN_4967; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4969 = 8'h69 == io_state_in_10 ? 8'hbb : _GEN_4968; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4970 = 8'h6a == io_state_in_10 ? 8'hbe : _GEN_4969; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4971 = 8'h6b == io_state_in_10 ? 8'hbd : _GEN_4970; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4972 = 8'h6c == io_state_in_10 ? 8'hb4 : _GEN_4971; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4973 = 8'h6d == io_state_in_10 ? 8'hb7 : _GEN_4972; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4974 = 8'h6e == io_state_in_10 ? 8'hb2 : _GEN_4973; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4975 = 8'h6f == io_state_in_10 ? 8'hb1 : _GEN_4974; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4976 = 8'h70 == io_state_in_10 ? 8'h90 : _GEN_4975; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4977 = 8'h71 == io_state_in_10 ? 8'h93 : _GEN_4976; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4978 = 8'h72 == io_state_in_10 ? 8'h96 : _GEN_4977; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4979 = 8'h73 == io_state_in_10 ? 8'h95 : _GEN_4978; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4980 = 8'h74 == io_state_in_10 ? 8'h9c : _GEN_4979; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4981 = 8'h75 == io_state_in_10 ? 8'h9f : _GEN_4980; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4982 = 8'h76 == io_state_in_10 ? 8'h9a : _GEN_4981; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4983 = 8'h77 == io_state_in_10 ? 8'h99 : _GEN_4982; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4984 = 8'h78 == io_state_in_10 ? 8'h88 : _GEN_4983; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4985 = 8'h79 == io_state_in_10 ? 8'h8b : _GEN_4984; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4986 = 8'h7a == io_state_in_10 ? 8'h8e : _GEN_4985; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4987 = 8'h7b == io_state_in_10 ? 8'h8d : _GEN_4986; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4988 = 8'h7c == io_state_in_10 ? 8'h84 : _GEN_4987; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4989 = 8'h7d == io_state_in_10 ? 8'h87 : _GEN_4988; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4990 = 8'h7e == io_state_in_10 ? 8'h82 : _GEN_4989; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4991 = 8'h7f == io_state_in_10 ? 8'h81 : _GEN_4990; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4992 = 8'h80 == io_state_in_10 ? 8'h9b : _GEN_4991; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4993 = 8'h81 == io_state_in_10 ? 8'h98 : _GEN_4992; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4994 = 8'h82 == io_state_in_10 ? 8'h9d : _GEN_4993; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4995 = 8'h83 == io_state_in_10 ? 8'h9e : _GEN_4994; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4996 = 8'h84 == io_state_in_10 ? 8'h97 : _GEN_4995; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4997 = 8'h85 == io_state_in_10 ? 8'h94 : _GEN_4996; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4998 = 8'h86 == io_state_in_10 ? 8'h91 : _GEN_4997; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_4999 = 8'h87 == io_state_in_10 ? 8'h92 : _GEN_4998; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5000 = 8'h88 == io_state_in_10 ? 8'h83 : _GEN_4999; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5001 = 8'h89 == io_state_in_10 ? 8'h80 : _GEN_5000; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5002 = 8'h8a == io_state_in_10 ? 8'h85 : _GEN_5001; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5003 = 8'h8b == io_state_in_10 ? 8'h86 : _GEN_5002; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5004 = 8'h8c == io_state_in_10 ? 8'h8f : _GEN_5003; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5005 = 8'h8d == io_state_in_10 ? 8'h8c : _GEN_5004; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5006 = 8'h8e == io_state_in_10 ? 8'h89 : _GEN_5005; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5007 = 8'h8f == io_state_in_10 ? 8'h8a : _GEN_5006; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5008 = 8'h90 == io_state_in_10 ? 8'hab : _GEN_5007; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5009 = 8'h91 == io_state_in_10 ? 8'ha8 : _GEN_5008; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5010 = 8'h92 == io_state_in_10 ? 8'had : _GEN_5009; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5011 = 8'h93 == io_state_in_10 ? 8'hae : _GEN_5010; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5012 = 8'h94 == io_state_in_10 ? 8'ha7 : _GEN_5011; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5013 = 8'h95 == io_state_in_10 ? 8'ha4 : _GEN_5012; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5014 = 8'h96 == io_state_in_10 ? 8'ha1 : _GEN_5013; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5015 = 8'h97 == io_state_in_10 ? 8'ha2 : _GEN_5014; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5016 = 8'h98 == io_state_in_10 ? 8'hb3 : _GEN_5015; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5017 = 8'h99 == io_state_in_10 ? 8'hb0 : _GEN_5016; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5018 = 8'h9a == io_state_in_10 ? 8'hb5 : _GEN_5017; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5019 = 8'h9b == io_state_in_10 ? 8'hb6 : _GEN_5018; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5020 = 8'h9c == io_state_in_10 ? 8'hbf : _GEN_5019; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5021 = 8'h9d == io_state_in_10 ? 8'hbc : _GEN_5020; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5022 = 8'h9e == io_state_in_10 ? 8'hb9 : _GEN_5021; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5023 = 8'h9f == io_state_in_10 ? 8'hba : _GEN_5022; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5024 = 8'ha0 == io_state_in_10 ? 8'hfb : _GEN_5023; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5025 = 8'ha1 == io_state_in_10 ? 8'hf8 : _GEN_5024; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5026 = 8'ha2 == io_state_in_10 ? 8'hfd : _GEN_5025; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5027 = 8'ha3 == io_state_in_10 ? 8'hfe : _GEN_5026; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5028 = 8'ha4 == io_state_in_10 ? 8'hf7 : _GEN_5027; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5029 = 8'ha5 == io_state_in_10 ? 8'hf4 : _GEN_5028; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5030 = 8'ha6 == io_state_in_10 ? 8'hf1 : _GEN_5029; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5031 = 8'ha7 == io_state_in_10 ? 8'hf2 : _GEN_5030; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5032 = 8'ha8 == io_state_in_10 ? 8'he3 : _GEN_5031; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5033 = 8'ha9 == io_state_in_10 ? 8'he0 : _GEN_5032; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5034 = 8'haa == io_state_in_10 ? 8'he5 : _GEN_5033; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5035 = 8'hab == io_state_in_10 ? 8'he6 : _GEN_5034; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5036 = 8'hac == io_state_in_10 ? 8'hef : _GEN_5035; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5037 = 8'had == io_state_in_10 ? 8'hec : _GEN_5036; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5038 = 8'hae == io_state_in_10 ? 8'he9 : _GEN_5037; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5039 = 8'haf == io_state_in_10 ? 8'hea : _GEN_5038; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5040 = 8'hb0 == io_state_in_10 ? 8'hcb : _GEN_5039; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5041 = 8'hb1 == io_state_in_10 ? 8'hc8 : _GEN_5040; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5042 = 8'hb2 == io_state_in_10 ? 8'hcd : _GEN_5041; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5043 = 8'hb3 == io_state_in_10 ? 8'hce : _GEN_5042; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5044 = 8'hb4 == io_state_in_10 ? 8'hc7 : _GEN_5043; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5045 = 8'hb5 == io_state_in_10 ? 8'hc4 : _GEN_5044; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5046 = 8'hb6 == io_state_in_10 ? 8'hc1 : _GEN_5045; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5047 = 8'hb7 == io_state_in_10 ? 8'hc2 : _GEN_5046; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5048 = 8'hb8 == io_state_in_10 ? 8'hd3 : _GEN_5047; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5049 = 8'hb9 == io_state_in_10 ? 8'hd0 : _GEN_5048; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5050 = 8'hba == io_state_in_10 ? 8'hd5 : _GEN_5049; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5051 = 8'hbb == io_state_in_10 ? 8'hd6 : _GEN_5050; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5052 = 8'hbc == io_state_in_10 ? 8'hdf : _GEN_5051; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5053 = 8'hbd == io_state_in_10 ? 8'hdc : _GEN_5052; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5054 = 8'hbe == io_state_in_10 ? 8'hd9 : _GEN_5053; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5055 = 8'hbf == io_state_in_10 ? 8'hda : _GEN_5054; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5056 = 8'hc0 == io_state_in_10 ? 8'h5b : _GEN_5055; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5057 = 8'hc1 == io_state_in_10 ? 8'h58 : _GEN_5056; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5058 = 8'hc2 == io_state_in_10 ? 8'h5d : _GEN_5057; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5059 = 8'hc3 == io_state_in_10 ? 8'h5e : _GEN_5058; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5060 = 8'hc4 == io_state_in_10 ? 8'h57 : _GEN_5059; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5061 = 8'hc5 == io_state_in_10 ? 8'h54 : _GEN_5060; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5062 = 8'hc6 == io_state_in_10 ? 8'h51 : _GEN_5061; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5063 = 8'hc7 == io_state_in_10 ? 8'h52 : _GEN_5062; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5064 = 8'hc8 == io_state_in_10 ? 8'h43 : _GEN_5063; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5065 = 8'hc9 == io_state_in_10 ? 8'h40 : _GEN_5064; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5066 = 8'hca == io_state_in_10 ? 8'h45 : _GEN_5065; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5067 = 8'hcb == io_state_in_10 ? 8'h46 : _GEN_5066; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5068 = 8'hcc == io_state_in_10 ? 8'h4f : _GEN_5067; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5069 = 8'hcd == io_state_in_10 ? 8'h4c : _GEN_5068; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5070 = 8'hce == io_state_in_10 ? 8'h49 : _GEN_5069; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5071 = 8'hcf == io_state_in_10 ? 8'h4a : _GEN_5070; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5072 = 8'hd0 == io_state_in_10 ? 8'h6b : _GEN_5071; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5073 = 8'hd1 == io_state_in_10 ? 8'h68 : _GEN_5072; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5074 = 8'hd2 == io_state_in_10 ? 8'h6d : _GEN_5073; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5075 = 8'hd3 == io_state_in_10 ? 8'h6e : _GEN_5074; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5076 = 8'hd4 == io_state_in_10 ? 8'h67 : _GEN_5075; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5077 = 8'hd5 == io_state_in_10 ? 8'h64 : _GEN_5076; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5078 = 8'hd6 == io_state_in_10 ? 8'h61 : _GEN_5077; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5079 = 8'hd7 == io_state_in_10 ? 8'h62 : _GEN_5078; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5080 = 8'hd8 == io_state_in_10 ? 8'h73 : _GEN_5079; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5081 = 8'hd9 == io_state_in_10 ? 8'h70 : _GEN_5080; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5082 = 8'hda == io_state_in_10 ? 8'h75 : _GEN_5081; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5083 = 8'hdb == io_state_in_10 ? 8'h76 : _GEN_5082; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5084 = 8'hdc == io_state_in_10 ? 8'h7f : _GEN_5083; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5085 = 8'hdd == io_state_in_10 ? 8'h7c : _GEN_5084; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5086 = 8'hde == io_state_in_10 ? 8'h79 : _GEN_5085; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5087 = 8'hdf == io_state_in_10 ? 8'h7a : _GEN_5086; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5088 = 8'he0 == io_state_in_10 ? 8'h3b : _GEN_5087; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5089 = 8'he1 == io_state_in_10 ? 8'h38 : _GEN_5088; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5090 = 8'he2 == io_state_in_10 ? 8'h3d : _GEN_5089; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5091 = 8'he3 == io_state_in_10 ? 8'h3e : _GEN_5090; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5092 = 8'he4 == io_state_in_10 ? 8'h37 : _GEN_5091; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5093 = 8'he5 == io_state_in_10 ? 8'h34 : _GEN_5092; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5094 = 8'he6 == io_state_in_10 ? 8'h31 : _GEN_5093; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5095 = 8'he7 == io_state_in_10 ? 8'h32 : _GEN_5094; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5096 = 8'he8 == io_state_in_10 ? 8'h23 : _GEN_5095; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5097 = 8'he9 == io_state_in_10 ? 8'h20 : _GEN_5096; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5098 = 8'hea == io_state_in_10 ? 8'h25 : _GEN_5097; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5099 = 8'heb == io_state_in_10 ? 8'h26 : _GEN_5098; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5100 = 8'hec == io_state_in_10 ? 8'h2f : _GEN_5099; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5101 = 8'hed == io_state_in_10 ? 8'h2c : _GEN_5100; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5102 = 8'hee == io_state_in_10 ? 8'h29 : _GEN_5101; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5103 = 8'hef == io_state_in_10 ? 8'h2a : _GEN_5102; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5104 = 8'hf0 == io_state_in_10 ? 8'hb : _GEN_5103; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5105 = 8'hf1 == io_state_in_10 ? 8'h8 : _GEN_5104; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5106 = 8'hf2 == io_state_in_10 ? 8'hd : _GEN_5105; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5107 = 8'hf3 == io_state_in_10 ? 8'he : _GEN_5106; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5108 = 8'hf4 == io_state_in_10 ? 8'h7 : _GEN_5107; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5109 = 8'hf5 == io_state_in_10 ? 8'h4 : _GEN_5108; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5110 = 8'hf6 == io_state_in_10 ? 8'h1 : _GEN_5109; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5111 = 8'hf7 == io_state_in_10 ? 8'h2 : _GEN_5110; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5112 = 8'hf8 == io_state_in_10 ? 8'h13 : _GEN_5111; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5113 = 8'hf9 == io_state_in_10 ? 8'h10 : _GEN_5112; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5114 = 8'hfa == io_state_in_10 ? 8'h15 : _GEN_5113; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5115 = 8'hfb == io_state_in_10 ? 8'h16 : _GEN_5114; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5116 = 8'hfc == io_state_in_10 ? 8'h1f : _GEN_5115; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5117 = 8'hfd == io_state_in_10 ? 8'h1c : _GEN_5116; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5118 = 8'hfe == io_state_in_10 ? 8'h19 : _GEN_5117; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _GEN_5119 = 8'hff == io_state_in_10 ? 8'h1a : _GEN_5118; // @[MixColumns.scala 136:{58,58}]
  wire [7:0] _tmp_state_9_T_1 = _tmp_state_9_T ^ _GEN_5119; // @[MixColumns.scala 136:58]
  wire [7:0] _tmp_state_10_T = io_state_in_8 ^ io_state_in_9; // @[MixColumns.scala 137:35]
  wire [7:0] _GEN_5121 = 8'h1 == io_state_in_10 ? 8'h2 : 8'h0; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5122 = 8'h2 == io_state_in_10 ? 8'h4 : _GEN_5121; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5123 = 8'h3 == io_state_in_10 ? 8'h6 : _GEN_5122; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5124 = 8'h4 == io_state_in_10 ? 8'h8 : _GEN_5123; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5125 = 8'h5 == io_state_in_10 ? 8'ha : _GEN_5124; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5126 = 8'h6 == io_state_in_10 ? 8'hc : _GEN_5125; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5127 = 8'h7 == io_state_in_10 ? 8'he : _GEN_5126; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5128 = 8'h8 == io_state_in_10 ? 8'h10 : _GEN_5127; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5129 = 8'h9 == io_state_in_10 ? 8'h12 : _GEN_5128; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5130 = 8'ha == io_state_in_10 ? 8'h14 : _GEN_5129; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5131 = 8'hb == io_state_in_10 ? 8'h16 : _GEN_5130; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5132 = 8'hc == io_state_in_10 ? 8'h18 : _GEN_5131; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5133 = 8'hd == io_state_in_10 ? 8'h1a : _GEN_5132; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5134 = 8'he == io_state_in_10 ? 8'h1c : _GEN_5133; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5135 = 8'hf == io_state_in_10 ? 8'h1e : _GEN_5134; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5136 = 8'h10 == io_state_in_10 ? 8'h20 : _GEN_5135; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5137 = 8'h11 == io_state_in_10 ? 8'h22 : _GEN_5136; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5138 = 8'h12 == io_state_in_10 ? 8'h24 : _GEN_5137; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5139 = 8'h13 == io_state_in_10 ? 8'h26 : _GEN_5138; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5140 = 8'h14 == io_state_in_10 ? 8'h28 : _GEN_5139; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5141 = 8'h15 == io_state_in_10 ? 8'h2a : _GEN_5140; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5142 = 8'h16 == io_state_in_10 ? 8'h2c : _GEN_5141; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5143 = 8'h17 == io_state_in_10 ? 8'h2e : _GEN_5142; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5144 = 8'h18 == io_state_in_10 ? 8'h30 : _GEN_5143; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5145 = 8'h19 == io_state_in_10 ? 8'h32 : _GEN_5144; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5146 = 8'h1a == io_state_in_10 ? 8'h34 : _GEN_5145; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5147 = 8'h1b == io_state_in_10 ? 8'h36 : _GEN_5146; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5148 = 8'h1c == io_state_in_10 ? 8'h38 : _GEN_5147; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5149 = 8'h1d == io_state_in_10 ? 8'h3a : _GEN_5148; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5150 = 8'h1e == io_state_in_10 ? 8'h3c : _GEN_5149; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5151 = 8'h1f == io_state_in_10 ? 8'h3e : _GEN_5150; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5152 = 8'h20 == io_state_in_10 ? 8'h40 : _GEN_5151; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5153 = 8'h21 == io_state_in_10 ? 8'h42 : _GEN_5152; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5154 = 8'h22 == io_state_in_10 ? 8'h44 : _GEN_5153; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5155 = 8'h23 == io_state_in_10 ? 8'h46 : _GEN_5154; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5156 = 8'h24 == io_state_in_10 ? 8'h48 : _GEN_5155; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5157 = 8'h25 == io_state_in_10 ? 8'h4a : _GEN_5156; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5158 = 8'h26 == io_state_in_10 ? 8'h4c : _GEN_5157; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5159 = 8'h27 == io_state_in_10 ? 8'h4e : _GEN_5158; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5160 = 8'h28 == io_state_in_10 ? 8'h50 : _GEN_5159; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5161 = 8'h29 == io_state_in_10 ? 8'h52 : _GEN_5160; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5162 = 8'h2a == io_state_in_10 ? 8'h54 : _GEN_5161; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5163 = 8'h2b == io_state_in_10 ? 8'h56 : _GEN_5162; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5164 = 8'h2c == io_state_in_10 ? 8'h58 : _GEN_5163; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5165 = 8'h2d == io_state_in_10 ? 8'h5a : _GEN_5164; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5166 = 8'h2e == io_state_in_10 ? 8'h5c : _GEN_5165; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5167 = 8'h2f == io_state_in_10 ? 8'h5e : _GEN_5166; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5168 = 8'h30 == io_state_in_10 ? 8'h60 : _GEN_5167; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5169 = 8'h31 == io_state_in_10 ? 8'h62 : _GEN_5168; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5170 = 8'h32 == io_state_in_10 ? 8'h64 : _GEN_5169; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5171 = 8'h33 == io_state_in_10 ? 8'h66 : _GEN_5170; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5172 = 8'h34 == io_state_in_10 ? 8'h68 : _GEN_5171; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5173 = 8'h35 == io_state_in_10 ? 8'h6a : _GEN_5172; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5174 = 8'h36 == io_state_in_10 ? 8'h6c : _GEN_5173; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5175 = 8'h37 == io_state_in_10 ? 8'h6e : _GEN_5174; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5176 = 8'h38 == io_state_in_10 ? 8'h70 : _GEN_5175; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5177 = 8'h39 == io_state_in_10 ? 8'h72 : _GEN_5176; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5178 = 8'h3a == io_state_in_10 ? 8'h74 : _GEN_5177; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5179 = 8'h3b == io_state_in_10 ? 8'h76 : _GEN_5178; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5180 = 8'h3c == io_state_in_10 ? 8'h78 : _GEN_5179; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5181 = 8'h3d == io_state_in_10 ? 8'h7a : _GEN_5180; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5182 = 8'h3e == io_state_in_10 ? 8'h7c : _GEN_5181; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5183 = 8'h3f == io_state_in_10 ? 8'h7e : _GEN_5182; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5184 = 8'h40 == io_state_in_10 ? 8'h80 : _GEN_5183; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5185 = 8'h41 == io_state_in_10 ? 8'h82 : _GEN_5184; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5186 = 8'h42 == io_state_in_10 ? 8'h84 : _GEN_5185; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5187 = 8'h43 == io_state_in_10 ? 8'h86 : _GEN_5186; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5188 = 8'h44 == io_state_in_10 ? 8'h88 : _GEN_5187; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5189 = 8'h45 == io_state_in_10 ? 8'h8a : _GEN_5188; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5190 = 8'h46 == io_state_in_10 ? 8'h8c : _GEN_5189; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5191 = 8'h47 == io_state_in_10 ? 8'h8e : _GEN_5190; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5192 = 8'h48 == io_state_in_10 ? 8'h90 : _GEN_5191; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5193 = 8'h49 == io_state_in_10 ? 8'h92 : _GEN_5192; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5194 = 8'h4a == io_state_in_10 ? 8'h94 : _GEN_5193; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5195 = 8'h4b == io_state_in_10 ? 8'h96 : _GEN_5194; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5196 = 8'h4c == io_state_in_10 ? 8'h98 : _GEN_5195; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5197 = 8'h4d == io_state_in_10 ? 8'h9a : _GEN_5196; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5198 = 8'h4e == io_state_in_10 ? 8'h9c : _GEN_5197; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5199 = 8'h4f == io_state_in_10 ? 8'h9e : _GEN_5198; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5200 = 8'h50 == io_state_in_10 ? 8'ha0 : _GEN_5199; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5201 = 8'h51 == io_state_in_10 ? 8'ha2 : _GEN_5200; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5202 = 8'h52 == io_state_in_10 ? 8'ha4 : _GEN_5201; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5203 = 8'h53 == io_state_in_10 ? 8'ha6 : _GEN_5202; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5204 = 8'h54 == io_state_in_10 ? 8'ha8 : _GEN_5203; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5205 = 8'h55 == io_state_in_10 ? 8'haa : _GEN_5204; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5206 = 8'h56 == io_state_in_10 ? 8'hac : _GEN_5205; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5207 = 8'h57 == io_state_in_10 ? 8'hae : _GEN_5206; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5208 = 8'h58 == io_state_in_10 ? 8'hb0 : _GEN_5207; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5209 = 8'h59 == io_state_in_10 ? 8'hb2 : _GEN_5208; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5210 = 8'h5a == io_state_in_10 ? 8'hb4 : _GEN_5209; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5211 = 8'h5b == io_state_in_10 ? 8'hb6 : _GEN_5210; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5212 = 8'h5c == io_state_in_10 ? 8'hb8 : _GEN_5211; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5213 = 8'h5d == io_state_in_10 ? 8'hba : _GEN_5212; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5214 = 8'h5e == io_state_in_10 ? 8'hbc : _GEN_5213; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5215 = 8'h5f == io_state_in_10 ? 8'hbe : _GEN_5214; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5216 = 8'h60 == io_state_in_10 ? 8'hc0 : _GEN_5215; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5217 = 8'h61 == io_state_in_10 ? 8'hc2 : _GEN_5216; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5218 = 8'h62 == io_state_in_10 ? 8'hc4 : _GEN_5217; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5219 = 8'h63 == io_state_in_10 ? 8'hc6 : _GEN_5218; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5220 = 8'h64 == io_state_in_10 ? 8'hc8 : _GEN_5219; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5221 = 8'h65 == io_state_in_10 ? 8'hca : _GEN_5220; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5222 = 8'h66 == io_state_in_10 ? 8'hcc : _GEN_5221; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5223 = 8'h67 == io_state_in_10 ? 8'hce : _GEN_5222; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5224 = 8'h68 == io_state_in_10 ? 8'hd0 : _GEN_5223; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5225 = 8'h69 == io_state_in_10 ? 8'hd2 : _GEN_5224; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5226 = 8'h6a == io_state_in_10 ? 8'hd4 : _GEN_5225; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5227 = 8'h6b == io_state_in_10 ? 8'hd6 : _GEN_5226; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5228 = 8'h6c == io_state_in_10 ? 8'hd8 : _GEN_5227; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5229 = 8'h6d == io_state_in_10 ? 8'hda : _GEN_5228; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5230 = 8'h6e == io_state_in_10 ? 8'hdc : _GEN_5229; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5231 = 8'h6f == io_state_in_10 ? 8'hde : _GEN_5230; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5232 = 8'h70 == io_state_in_10 ? 8'he0 : _GEN_5231; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5233 = 8'h71 == io_state_in_10 ? 8'he2 : _GEN_5232; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5234 = 8'h72 == io_state_in_10 ? 8'he4 : _GEN_5233; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5235 = 8'h73 == io_state_in_10 ? 8'he6 : _GEN_5234; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5236 = 8'h74 == io_state_in_10 ? 8'he8 : _GEN_5235; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5237 = 8'h75 == io_state_in_10 ? 8'hea : _GEN_5236; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5238 = 8'h76 == io_state_in_10 ? 8'hec : _GEN_5237; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5239 = 8'h77 == io_state_in_10 ? 8'hee : _GEN_5238; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5240 = 8'h78 == io_state_in_10 ? 8'hf0 : _GEN_5239; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5241 = 8'h79 == io_state_in_10 ? 8'hf2 : _GEN_5240; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5242 = 8'h7a == io_state_in_10 ? 8'hf4 : _GEN_5241; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5243 = 8'h7b == io_state_in_10 ? 8'hf6 : _GEN_5242; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5244 = 8'h7c == io_state_in_10 ? 8'hf8 : _GEN_5243; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5245 = 8'h7d == io_state_in_10 ? 8'hfa : _GEN_5244; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5246 = 8'h7e == io_state_in_10 ? 8'hfc : _GEN_5245; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5247 = 8'h7f == io_state_in_10 ? 8'hfe : _GEN_5246; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5248 = 8'h80 == io_state_in_10 ? 8'h1b : _GEN_5247; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5249 = 8'h81 == io_state_in_10 ? 8'h19 : _GEN_5248; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5250 = 8'h82 == io_state_in_10 ? 8'h1f : _GEN_5249; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5251 = 8'h83 == io_state_in_10 ? 8'h1d : _GEN_5250; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5252 = 8'h84 == io_state_in_10 ? 8'h13 : _GEN_5251; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5253 = 8'h85 == io_state_in_10 ? 8'h11 : _GEN_5252; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5254 = 8'h86 == io_state_in_10 ? 8'h17 : _GEN_5253; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5255 = 8'h87 == io_state_in_10 ? 8'h15 : _GEN_5254; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5256 = 8'h88 == io_state_in_10 ? 8'hb : _GEN_5255; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5257 = 8'h89 == io_state_in_10 ? 8'h9 : _GEN_5256; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5258 = 8'h8a == io_state_in_10 ? 8'hf : _GEN_5257; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5259 = 8'h8b == io_state_in_10 ? 8'hd : _GEN_5258; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5260 = 8'h8c == io_state_in_10 ? 8'h3 : _GEN_5259; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5261 = 8'h8d == io_state_in_10 ? 8'h1 : _GEN_5260; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5262 = 8'h8e == io_state_in_10 ? 8'h7 : _GEN_5261; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5263 = 8'h8f == io_state_in_10 ? 8'h5 : _GEN_5262; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5264 = 8'h90 == io_state_in_10 ? 8'h3b : _GEN_5263; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5265 = 8'h91 == io_state_in_10 ? 8'h39 : _GEN_5264; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5266 = 8'h92 == io_state_in_10 ? 8'h3f : _GEN_5265; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5267 = 8'h93 == io_state_in_10 ? 8'h3d : _GEN_5266; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5268 = 8'h94 == io_state_in_10 ? 8'h33 : _GEN_5267; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5269 = 8'h95 == io_state_in_10 ? 8'h31 : _GEN_5268; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5270 = 8'h96 == io_state_in_10 ? 8'h37 : _GEN_5269; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5271 = 8'h97 == io_state_in_10 ? 8'h35 : _GEN_5270; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5272 = 8'h98 == io_state_in_10 ? 8'h2b : _GEN_5271; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5273 = 8'h99 == io_state_in_10 ? 8'h29 : _GEN_5272; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5274 = 8'h9a == io_state_in_10 ? 8'h2f : _GEN_5273; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5275 = 8'h9b == io_state_in_10 ? 8'h2d : _GEN_5274; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5276 = 8'h9c == io_state_in_10 ? 8'h23 : _GEN_5275; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5277 = 8'h9d == io_state_in_10 ? 8'h21 : _GEN_5276; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5278 = 8'h9e == io_state_in_10 ? 8'h27 : _GEN_5277; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5279 = 8'h9f == io_state_in_10 ? 8'h25 : _GEN_5278; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5280 = 8'ha0 == io_state_in_10 ? 8'h5b : _GEN_5279; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5281 = 8'ha1 == io_state_in_10 ? 8'h59 : _GEN_5280; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5282 = 8'ha2 == io_state_in_10 ? 8'h5f : _GEN_5281; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5283 = 8'ha3 == io_state_in_10 ? 8'h5d : _GEN_5282; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5284 = 8'ha4 == io_state_in_10 ? 8'h53 : _GEN_5283; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5285 = 8'ha5 == io_state_in_10 ? 8'h51 : _GEN_5284; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5286 = 8'ha6 == io_state_in_10 ? 8'h57 : _GEN_5285; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5287 = 8'ha7 == io_state_in_10 ? 8'h55 : _GEN_5286; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5288 = 8'ha8 == io_state_in_10 ? 8'h4b : _GEN_5287; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5289 = 8'ha9 == io_state_in_10 ? 8'h49 : _GEN_5288; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5290 = 8'haa == io_state_in_10 ? 8'h4f : _GEN_5289; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5291 = 8'hab == io_state_in_10 ? 8'h4d : _GEN_5290; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5292 = 8'hac == io_state_in_10 ? 8'h43 : _GEN_5291; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5293 = 8'had == io_state_in_10 ? 8'h41 : _GEN_5292; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5294 = 8'hae == io_state_in_10 ? 8'h47 : _GEN_5293; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5295 = 8'haf == io_state_in_10 ? 8'h45 : _GEN_5294; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5296 = 8'hb0 == io_state_in_10 ? 8'h7b : _GEN_5295; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5297 = 8'hb1 == io_state_in_10 ? 8'h79 : _GEN_5296; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5298 = 8'hb2 == io_state_in_10 ? 8'h7f : _GEN_5297; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5299 = 8'hb3 == io_state_in_10 ? 8'h7d : _GEN_5298; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5300 = 8'hb4 == io_state_in_10 ? 8'h73 : _GEN_5299; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5301 = 8'hb5 == io_state_in_10 ? 8'h71 : _GEN_5300; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5302 = 8'hb6 == io_state_in_10 ? 8'h77 : _GEN_5301; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5303 = 8'hb7 == io_state_in_10 ? 8'h75 : _GEN_5302; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5304 = 8'hb8 == io_state_in_10 ? 8'h6b : _GEN_5303; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5305 = 8'hb9 == io_state_in_10 ? 8'h69 : _GEN_5304; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5306 = 8'hba == io_state_in_10 ? 8'h6f : _GEN_5305; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5307 = 8'hbb == io_state_in_10 ? 8'h6d : _GEN_5306; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5308 = 8'hbc == io_state_in_10 ? 8'h63 : _GEN_5307; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5309 = 8'hbd == io_state_in_10 ? 8'h61 : _GEN_5308; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5310 = 8'hbe == io_state_in_10 ? 8'h67 : _GEN_5309; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5311 = 8'hbf == io_state_in_10 ? 8'h65 : _GEN_5310; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5312 = 8'hc0 == io_state_in_10 ? 8'h9b : _GEN_5311; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5313 = 8'hc1 == io_state_in_10 ? 8'h99 : _GEN_5312; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5314 = 8'hc2 == io_state_in_10 ? 8'h9f : _GEN_5313; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5315 = 8'hc3 == io_state_in_10 ? 8'h9d : _GEN_5314; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5316 = 8'hc4 == io_state_in_10 ? 8'h93 : _GEN_5315; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5317 = 8'hc5 == io_state_in_10 ? 8'h91 : _GEN_5316; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5318 = 8'hc6 == io_state_in_10 ? 8'h97 : _GEN_5317; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5319 = 8'hc7 == io_state_in_10 ? 8'h95 : _GEN_5318; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5320 = 8'hc8 == io_state_in_10 ? 8'h8b : _GEN_5319; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5321 = 8'hc9 == io_state_in_10 ? 8'h89 : _GEN_5320; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5322 = 8'hca == io_state_in_10 ? 8'h8f : _GEN_5321; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5323 = 8'hcb == io_state_in_10 ? 8'h8d : _GEN_5322; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5324 = 8'hcc == io_state_in_10 ? 8'h83 : _GEN_5323; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5325 = 8'hcd == io_state_in_10 ? 8'h81 : _GEN_5324; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5326 = 8'hce == io_state_in_10 ? 8'h87 : _GEN_5325; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5327 = 8'hcf == io_state_in_10 ? 8'h85 : _GEN_5326; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5328 = 8'hd0 == io_state_in_10 ? 8'hbb : _GEN_5327; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5329 = 8'hd1 == io_state_in_10 ? 8'hb9 : _GEN_5328; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5330 = 8'hd2 == io_state_in_10 ? 8'hbf : _GEN_5329; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5331 = 8'hd3 == io_state_in_10 ? 8'hbd : _GEN_5330; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5332 = 8'hd4 == io_state_in_10 ? 8'hb3 : _GEN_5331; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5333 = 8'hd5 == io_state_in_10 ? 8'hb1 : _GEN_5332; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5334 = 8'hd6 == io_state_in_10 ? 8'hb7 : _GEN_5333; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5335 = 8'hd7 == io_state_in_10 ? 8'hb5 : _GEN_5334; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5336 = 8'hd8 == io_state_in_10 ? 8'hab : _GEN_5335; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5337 = 8'hd9 == io_state_in_10 ? 8'ha9 : _GEN_5336; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5338 = 8'hda == io_state_in_10 ? 8'haf : _GEN_5337; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5339 = 8'hdb == io_state_in_10 ? 8'had : _GEN_5338; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5340 = 8'hdc == io_state_in_10 ? 8'ha3 : _GEN_5339; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5341 = 8'hdd == io_state_in_10 ? 8'ha1 : _GEN_5340; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5342 = 8'hde == io_state_in_10 ? 8'ha7 : _GEN_5341; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5343 = 8'hdf == io_state_in_10 ? 8'ha5 : _GEN_5342; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5344 = 8'he0 == io_state_in_10 ? 8'hdb : _GEN_5343; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5345 = 8'he1 == io_state_in_10 ? 8'hd9 : _GEN_5344; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5346 = 8'he2 == io_state_in_10 ? 8'hdf : _GEN_5345; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5347 = 8'he3 == io_state_in_10 ? 8'hdd : _GEN_5346; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5348 = 8'he4 == io_state_in_10 ? 8'hd3 : _GEN_5347; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5349 = 8'he5 == io_state_in_10 ? 8'hd1 : _GEN_5348; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5350 = 8'he6 == io_state_in_10 ? 8'hd7 : _GEN_5349; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5351 = 8'he7 == io_state_in_10 ? 8'hd5 : _GEN_5350; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5352 = 8'he8 == io_state_in_10 ? 8'hcb : _GEN_5351; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5353 = 8'he9 == io_state_in_10 ? 8'hc9 : _GEN_5352; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5354 = 8'hea == io_state_in_10 ? 8'hcf : _GEN_5353; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5355 = 8'heb == io_state_in_10 ? 8'hcd : _GEN_5354; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5356 = 8'hec == io_state_in_10 ? 8'hc3 : _GEN_5355; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5357 = 8'hed == io_state_in_10 ? 8'hc1 : _GEN_5356; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5358 = 8'hee == io_state_in_10 ? 8'hc7 : _GEN_5357; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5359 = 8'hef == io_state_in_10 ? 8'hc5 : _GEN_5358; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5360 = 8'hf0 == io_state_in_10 ? 8'hfb : _GEN_5359; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5361 = 8'hf1 == io_state_in_10 ? 8'hf9 : _GEN_5360; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5362 = 8'hf2 == io_state_in_10 ? 8'hff : _GEN_5361; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5363 = 8'hf3 == io_state_in_10 ? 8'hfd : _GEN_5362; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5364 = 8'hf4 == io_state_in_10 ? 8'hf3 : _GEN_5363; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5365 = 8'hf5 == io_state_in_10 ? 8'hf1 : _GEN_5364; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5366 = 8'hf6 == io_state_in_10 ? 8'hf7 : _GEN_5365; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5367 = 8'hf7 == io_state_in_10 ? 8'hf5 : _GEN_5366; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5368 = 8'hf8 == io_state_in_10 ? 8'heb : _GEN_5367; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5369 = 8'hf9 == io_state_in_10 ? 8'he9 : _GEN_5368; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5370 = 8'hfa == io_state_in_10 ? 8'hef : _GEN_5369; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5371 = 8'hfb == io_state_in_10 ? 8'hed : _GEN_5370; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5372 = 8'hfc == io_state_in_10 ? 8'he3 : _GEN_5371; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5373 = 8'hfd == io_state_in_10 ? 8'he1 : _GEN_5372; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5374 = 8'hfe == io_state_in_10 ? 8'he7 : _GEN_5373; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _GEN_5375 = 8'hff == io_state_in_10 ? 8'he5 : _GEN_5374; // @[MixColumns.scala 137:{52,52}]
  wire [7:0] _tmp_state_10_T_1 = _tmp_state_10_T ^ _GEN_5375; // @[MixColumns.scala 137:52]
  wire [7:0] _GEN_5377 = 8'h1 == io_state_in_11 ? 8'h3 : 8'h0; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5378 = 8'h2 == io_state_in_11 ? 8'h6 : _GEN_5377; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5379 = 8'h3 == io_state_in_11 ? 8'h5 : _GEN_5378; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5380 = 8'h4 == io_state_in_11 ? 8'hc : _GEN_5379; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5381 = 8'h5 == io_state_in_11 ? 8'hf : _GEN_5380; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5382 = 8'h6 == io_state_in_11 ? 8'ha : _GEN_5381; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5383 = 8'h7 == io_state_in_11 ? 8'h9 : _GEN_5382; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5384 = 8'h8 == io_state_in_11 ? 8'h18 : _GEN_5383; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5385 = 8'h9 == io_state_in_11 ? 8'h1b : _GEN_5384; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5386 = 8'ha == io_state_in_11 ? 8'h1e : _GEN_5385; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5387 = 8'hb == io_state_in_11 ? 8'h1d : _GEN_5386; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5388 = 8'hc == io_state_in_11 ? 8'h14 : _GEN_5387; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5389 = 8'hd == io_state_in_11 ? 8'h17 : _GEN_5388; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5390 = 8'he == io_state_in_11 ? 8'h12 : _GEN_5389; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5391 = 8'hf == io_state_in_11 ? 8'h11 : _GEN_5390; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5392 = 8'h10 == io_state_in_11 ? 8'h30 : _GEN_5391; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5393 = 8'h11 == io_state_in_11 ? 8'h33 : _GEN_5392; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5394 = 8'h12 == io_state_in_11 ? 8'h36 : _GEN_5393; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5395 = 8'h13 == io_state_in_11 ? 8'h35 : _GEN_5394; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5396 = 8'h14 == io_state_in_11 ? 8'h3c : _GEN_5395; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5397 = 8'h15 == io_state_in_11 ? 8'h3f : _GEN_5396; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5398 = 8'h16 == io_state_in_11 ? 8'h3a : _GEN_5397; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5399 = 8'h17 == io_state_in_11 ? 8'h39 : _GEN_5398; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5400 = 8'h18 == io_state_in_11 ? 8'h28 : _GEN_5399; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5401 = 8'h19 == io_state_in_11 ? 8'h2b : _GEN_5400; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5402 = 8'h1a == io_state_in_11 ? 8'h2e : _GEN_5401; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5403 = 8'h1b == io_state_in_11 ? 8'h2d : _GEN_5402; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5404 = 8'h1c == io_state_in_11 ? 8'h24 : _GEN_5403; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5405 = 8'h1d == io_state_in_11 ? 8'h27 : _GEN_5404; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5406 = 8'h1e == io_state_in_11 ? 8'h22 : _GEN_5405; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5407 = 8'h1f == io_state_in_11 ? 8'h21 : _GEN_5406; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5408 = 8'h20 == io_state_in_11 ? 8'h60 : _GEN_5407; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5409 = 8'h21 == io_state_in_11 ? 8'h63 : _GEN_5408; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5410 = 8'h22 == io_state_in_11 ? 8'h66 : _GEN_5409; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5411 = 8'h23 == io_state_in_11 ? 8'h65 : _GEN_5410; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5412 = 8'h24 == io_state_in_11 ? 8'h6c : _GEN_5411; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5413 = 8'h25 == io_state_in_11 ? 8'h6f : _GEN_5412; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5414 = 8'h26 == io_state_in_11 ? 8'h6a : _GEN_5413; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5415 = 8'h27 == io_state_in_11 ? 8'h69 : _GEN_5414; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5416 = 8'h28 == io_state_in_11 ? 8'h78 : _GEN_5415; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5417 = 8'h29 == io_state_in_11 ? 8'h7b : _GEN_5416; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5418 = 8'h2a == io_state_in_11 ? 8'h7e : _GEN_5417; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5419 = 8'h2b == io_state_in_11 ? 8'h7d : _GEN_5418; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5420 = 8'h2c == io_state_in_11 ? 8'h74 : _GEN_5419; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5421 = 8'h2d == io_state_in_11 ? 8'h77 : _GEN_5420; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5422 = 8'h2e == io_state_in_11 ? 8'h72 : _GEN_5421; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5423 = 8'h2f == io_state_in_11 ? 8'h71 : _GEN_5422; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5424 = 8'h30 == io_state_in_11 ? 8'h50 : _GEN_5423; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5425 = 8'h31 == io_state_in_11 ? 8'h53 : _GEN_5424; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5426 = 8'h32 == io_state_in_11 ? 8'h56 : _GEN_5425; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5427 = 8'h33 == io_state_in_11 ? 8'h55 : _GEN_5426; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5428 = 8'h34 == io_state_in_11 ? 8'h5c : _GEN_5427; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5429 = 8'h35 == io_state_in_11 ? 8'h5f : _GEN_5428; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5430 = 8'h36 == io_state_in_11 ? 8'h5a : _GEN_5429; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5431 = 8'h37 == io_state_in_11 ? 8'h59 : _GEN_5430; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5432 = 8'h38 == io_state_in_11 ? 8'h48 : _GEN_5431; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5433 = 8'h39 == io_state_in_11 ? 8'h4b : _GEN_5432; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5434 = 8'h3a == io_state_in_11 ? 8'h4e : _GEN_5433; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5435 = 8'h3b == io_state_in_11 ? 8'h4d : _GEN_5434; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5436 = 8'h3c == io_state_in_11 ? 8'h44 : _GEN_5435; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5437 = 8'h3d == io_state_in_11 ? 8'h47 : _GEN_5436; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5438 = 8'h3e == io_state_in_11 ? 8'h42 : _GEN_5437; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5439 = 8'h3f == io_state_in_11 ? 8'h41 : _GEN_5438; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5440 = 8'h40 == io_state_in_11 ? 8'hc0 : _GEN_5439; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5441 = 8'h41 == io_state_in_11 ? 8'hc3 : _GEN_5440; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5442 = 8'h42 == io_state_in_11 ? 8'hc6 : _GEN_5441; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5443 = 8'h43 == io_state_in_11 ? 8'hc5 : _GEN_5442; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5444 = 8'h44 == io_state_in_11 ? 8'hcc : _GEN_5443; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5445 = 8'h45 == io_state_in_11 ? 8'hcf : _GEN_5444; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5446 = 8'h46 == io_state_in_11 ? 8'hca : _GEN_5445; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5447 = 8'h47 == io_state_in_11 ? 8'hc9 : _GEN_5446; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5448 = 8'h48 == io_state_in_11 ? 8'hd8 : _GEN_5447; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5449 = 8'h49 == io_state_in_11 ? 8'hdb : _GEN_5448; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5450 = 8'h4a == io_state_in_11 ? 8'hde : _GEN_5449; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5451 = 8'h4b == io_state_in_11 ? 8'hdd : _GEN_5450; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5452 = 8'h4c == io_state_in_11 ? 8'hd4 : _GEN_5451; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5453 = 8'h4d == io_state_in_11 ? 8'hd7 : _GEN_5452; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5454 = 8'h4e == io_state_in_11 ? 8'hd2 : _GEN_5453; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5455 = 8'h4f == io_state_in_11 ? 8'hd1 : _GEN_5454; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5456 = 8'h50 == io_state_in_11 ? 8'hf0 : _GEN_5455; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5457 = 8'h51 == io_state_in_11 ? 8'hf3 : _GEN_5456; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5458 = 8'h52 == io_state_in_11 ? 8'hf6 : _GEN_5457; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5459 = 8'h53 == io_state_in_11 ? 8'hf5 : _GEN_5458; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5460 = 8'h54 == io_state_in_11 ? 8'hfc : _GEN_5459; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5461 = 8'h55 == io_state_in_11 ? 8'hff : _GEN_5460; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5462 = 8'h56 == io_state_in_11 ? 8'hfa : _GEN_5461; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5463 = 8'h57 == io_state_in_11 ? 8'hf9 : _GEN_5462; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5464 = 8'h58 == io_state_in_11 ? 8'he8 : _GEN_5463; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5465 = 8'h59 == io_state_in_11 ? 8'heb : _GEN_5464; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5466 = 8'h5a == io_state_in_11 ? 8'hee : _GEN_5465; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5467 = 8'h5b == io_state_in_11 ? 8'hed : _GEN_5466; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5468 = 8'h5c == io_state_in_11 ? 8'he4 : _GEN_5467; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5469 = 8'h5d == io_state_in_11 ? 8'he7 : _GEN_5468; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5470 = 8'h5e == io_state_in_11 ? 8'he2 : _GEN_5469; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5471 = 8'h5f == io_state_in_11 ? 8'he1 : _GEN_5470; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5472 = 8'h60 == io_state_in_11 ? 8'ha0 : _GEN_5471; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5473 = 8'h61 == io_state_in_11 ? 8'ha3 : _GEN_5472; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5474 = 8'h62 == io_state_in_11 ? 8'ha6 : _GEN_5473; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5475 = 8'h63 == io_state_in_11 ? 8'ha5 : _GEN_5474; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5476 = 8'h64 == io_state_in_11 ? 8'hac : _GEN_5475; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5477 = 8'h65 == io_state_in_11 ? 8'haf : _GEN_5476; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5478 = 8'h66 == io_state_in_11 ? 8'haa : _GEN_5477; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5479 = 8'h67 == io_state_in_11 ? 8'ha9 : _GEN_5478; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5480 = 8'h68 == io_state_in_11 ? 8'hb8 : _GEN_5479; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5481 = 8'h69 == io_state_in_11 ? 8'hbb : _GEN_5480; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5482 = 8'h6a == io_state_in_11 ? 8'hbe : _GEN_5481; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5483 = 8'h6b == io_state_in_11 ? 8'hbd : _GEN_5482; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5484 = 8'h6c == io_state_in_11 ? 8'hb4 : _GEN_5483; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5485 = 8'h6d == io_state_in_11 ? 8'hb7 : _GEN_5484; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5486 = 8'h6e == io_state_in_11 ? 8'hb2 : _GEN_5485; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5487 = 8'h6f == io_state_in_11 ? 8'hb1 : _GEN_5486; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5488 = 8'h70 == io_state_in_11 ? 8'h90 : _GEN_5487; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5489 = 8'h71 == io_state_in_11 ? 8'h93 : _GEN_5488; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5490 = 8'h72 == io_state_in_11 ? 8'h96 : _GEN_5489; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5491 = 8'h73 == io_state_in_11 ? 8'h95 : _GEN_5490; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5492 = 8'h74 == io_state_in_11 ? 8'h9c : _GEN_5491; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5493 = 8'h75 == io_state_in_11 ? 8'h9f : _GEN_5492; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5494 = 8'h76 == io_state_in_11 ? 8'h9a : _GEN_5493; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5495 = 8'h77 == io_state_in_11 ? 8'h99 : _GEN_5494; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5496 = 8'h78 == io_state_in_11 ? 8'h88 : _GEN_5495; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5497 = 8'h79 == io_state_in_11 ? 8'h8b : _GEN_5496; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5498 = 8'h7a == io_state_in_11 ? 8'h8e : _GEN_5497; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5499 = 8'h7b == io_state_in_11 ? 8'h8d : _GEN_5498; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5500 = 8'h7c == io_state_in_11 ? 8'h84 : _GEN_5499; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5501 = 8'h7d == io_state_in_11 ? 8'h87 : _GEN_5500; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5502 = 8'h7e == io_state_in_11 ? 8'h82 : _GEN_5501; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5503 = 8'h7f == io_state_in_11 ? 8'h81 : _GEN_5502; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5504 = 8'h80 == io_state_in_11 ? 8'h9b : _GEN_5503; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5505 = 8'h81 == io_state_in_11 ? 8'h98 : _GEN_5504; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5506 = 8'h82 == io_state_in_11 ? 8'h9d : _GEN_5505; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5507 = 8'h83 == io_state_in_11 ? 8'h9e : _GEN_5506; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5508 = 8'h84 == io_state_in_11 ? 8'h97 : _GEN_5507; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5509 = 8'h85 == io_state_in_11 ? 8'h94 : _GEN_5508; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5510 = 8'h86 == io_state_in_11 ? 8'h91 : _GEN_5509; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5511 = 8'h87 == io_state_in_11 ? 8'h92 : _GEN_5510; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5512 = 8'h88 == io_state_in_11 ? 8'h83 : _GEN_5511; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5513 = 8'h89 == io_state_in_11 ? 8'h80 : _GEN_5512; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5514 = 8'h8a == io_state_in_11 ? 8'h85 : _GEN_5513; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5515 = 8'h8b == io_state_in_11 ? 8'h86 : _GEN_5514; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5516 = 8'h8c == io_state_in_11 ? 8'h8f : _GEN_5515; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5517 = 8'h8d == io_state_in_11 ? 8'h8c : _GEN_5516; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5518 = 8'h8e == io_state_in_11 ? 8'h89 : _GEN_5517; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5519 = 8'h8f == io_state_in_11 ? 8'h8a : _GEN_5518; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5520 = 8'h90 == io_state_in_11 ? 8'hab : _GEN_5519; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5521 = 8'h91 == io_state_in_11 ? 8'ha8 : _GEN_5520; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5522 = 8'h92 == io_state_in_11 ? 8'had : _GEN_5521; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5523 = 8'h93 == io_state_in_11 ? 8'hae : _GEN_5522; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5524 = 8'h94 == io_state_in_11 ? 8'ha7 : _GEN_5523; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5525 = 8'h95 == io_state_in_11 ? 8'ha4 : _GEN_5524; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5526 = 8'h96 == io_state_in_11 ? 8'ha1 : _GEN_5525; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5527 = 8'h97 == io_state_in_11 ? 8'ha2 : _GEN_5526; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5528 = 8'h98 == io_state_in_11 ? 8'hb3 : _GEN_5527; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5529 = 8'h99 == io_state_in_11 ? 8'hb0 : _GEN_5528; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5530 = 8'h9a == io_state_in_11 ? 8'hb5 : _GEN_5529; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5531 = 8'h9b == io_state_in_11 ? 8'hb6 : _GEN_5530; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5532 = 8'h9c == io_state_in_11 ? 8'hbf : _GEN_5531; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5533 = 8'h9d == io_state_in_11 ? 8'hbc : _GEN_5532; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5534 = 8'h9e == io_state_in_11 ? 8'hb9 : _GEN_5533; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5535 = 8'h9f == io_state_in_11 ? 8'hba : _GEN_5534; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5536 = 8'ha0 == io_state_in_11 ? 8'hfb : _GEN_5535; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5537 = 8'ha1 == io_state_in_11 ? 8'hf8 : _GEN_5536; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5538 = 8'ha2 == io_state_in_11 ? 8'hfd : _GEN_5537; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5539 = 8'ha3 == io_state_in_11 ? 8'hfe : _GEN_5538; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5540 = 8'ha4 == io_state_in_11 ? 8'hf7 : _GEN_5539; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5541 = 8'ha5 == io_state_in_11 ? 8'hf4 : _GEN_5540; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5542 = 8'ha6 == io_state_in_11 ? 8'hf1 : _GEN_5541; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5543 = 8'ha7 == io_state_in_11 ? 8'hf2 : _GEN_5542; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5544 = 8'ha8 == io_state_in_11 ? 8'he3 : _GEN_5543; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5545 = 8'ha9 == io_state_in_11 ? 8'he0 : _GEN_5544; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5546 = 8'haa == io_state_in_11 ? 8'he5 : _GEN_5545; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5547 = 8'hab == io_state_in_11 ? 8'he6 : _GEN_5546; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5548 = 8'hac == io_state_in_11 ? 8'hef : _GEN_5547; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5549 = 8'had == io_state_in_11 ? 8'hec : _GEN_5548; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5550 = 8'hae == io_state_in_11 ? 8'he9 : _GEN_5549; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5551 = 8'haf == io_state_in_11 ? 8'hea : _GEN_5550; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5552 = 8'hb0 == io_state_in_11 ? 8'hcb : _GEN_5551; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5553 = 8'hb1 == io_state_in_11 ? 8'hc8 : _GEN_5552; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5554 = 8'hb2 == io_state_in_11 ? 8'hcd : _GEN_5553; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5555 = 8'hb3 == io_state_in_11 ? 8'hce : _GEN_5554; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5556 = 8'hb4 == io_state_in_11 ? 8'hc7 : _GEN_5555; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5557 = 8'hb5 == io_state_in_11 ? 8'hc4 : _GEN_5556; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5558 = 8'hb6 == io_state_in_11 ? 8'hc1 : _GEN_5557; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5559 = 8'hb7 == io_state_in_11 ? 8'hc2 : _GEN_5558; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5560 = 8'hb8 == io_state_in_11 ? 8'hd3 : _GEN_5559; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5561 = 8'hb9 == io_state_in_11 ? 8'hd0 : _GEN_5560; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5562 = 8'hba == io_state_in_11 ? 8'hd5 : _GEN_5561; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5563 = 8'hbb == io_state_in_11 ? 8'hd6 : _GEN_5562; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5564 = 8'hbc == io_state_in_11 ? 8'hdf : _GEN_5563; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5565 = 8'hbd == io_state_in_11 ? 8'hdc : _GEN_5564; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5566 = 8'hbe == io_state_in_11 ? 8'hd9 : _GEN_5565; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5567 = 8'hbf == io_state_in_11 ? 8'hda : _GEN_5566; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5568 = 8'hc0 == io_state_in_11 ? 8'h5b : _GEN_5567; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5569 = 8'hc1 == io_state_in_11 ? 8'h58 : _GEN_5568; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5570 = 8'hc2 == io_state_in_11 ? 8'h5d : _GEN_5569; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5571 = 8'hc3 == io_state_in_11 ? 8'h5e : _GEN_5570; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5572 = 8'hc4 == io_state_in_11 ? 8'h57 : _GEN_5571; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5573 = 8'hc5 == io_state_in_11 ? 8'h54 : _GEN_5572; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5574 = 8'hc6 == io_state_in_11 ? 8'h51 : _GEN_5573; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5575 = 8'hc7 == io_state_in_11 ? 8'h52 : _GEN_5574; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5576 = 8'hc8 == io_state_in_11 ? 8'h43 : _GEN_5575; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5577 = 8'hc9 == io_state_in_11 ? 8'h40 : _GEN_5576; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5578 = 8'hca == io_state_in_11 ? 8'h45 : _GEN_5577; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5579 = 8'hcb == io_state_in_11 ? 8'h46 : _GEN_5578; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5580 = 8'hcc == io_state_in_11 ? 8'h4f : _GEN_5579; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5581 = 8'hcd == io_state_in_11 ? 8'h4c : _GEN_5580; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5582 = 8'hce == io_state_in_11 ? 8'h49 : _GEN_5581; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5583 = 8'hcf == io_state_in_11 ? 8'h4a : _GEN_5582; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5584 = 8'hd0 == io_state_in_11 ? 8'h6b : _GEN_5583; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5585 = 8'hd1 == io_state_in_11 ? 8'h68 : _GEN_5584; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5586 = 8'hd2 == io_state_in_11 ? 8'h6d : _GEN_5585; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5587 = 8'hd3 == io_state_in_11 ? 8'h6e : _GEN_5586; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5588 = 8'hd4 == io_state_in_11 ? 8'h67 : _GEN_5587; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5589 = 8'hd5 == io_state_in_11 ? 8'h64 : _GEN_5588; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5590 = 8'hd6 == io_state_in_11 ? 8'h61 : _GEN_5589; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5591 = 8'hd7 == io_state_in_11 ? 8'h62 : _GEN_5590; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5592 = 8'hd8 == io_state_in_11 ? 8'h73 : _GEN_5591; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5593 = 8'hd9 == io_state_in_11 ? 8'h70 : _GEN_5592; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5594 = 8'hda == io_state_in_11 ? 8'h75 : _GEN_5593; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5595 = 8'hdb == io_state_in_11 ? 8'h76 : _GEN_5594; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5596 = 8'hdc == io_state_in_11 ? 8'h7f : _GEN_5595; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5597 = 8'hdd == io_state_in_11 ? 8'h7c : _GEN_5596; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5598 = 8'hde == io_state_in_11 ? 8'h79 : _GEN_5597; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5599 = 8'hdf == io_state_in_11 ? 8'h7a : _GEN_5598; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5600 = 8'he0 == io_state_in_11 ? 8'h3b : _GEN_5599; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5601 = 8'he1 == io_state_in_11 ? 8'h38 : _GEN_5600; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5602 = 8'he2 == io_state_in_11 ? 8'h3d : _GEN_5601; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5603 = 8'he3 == io_state_in_11 ? 8'h3e : _GEN_5602; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5604 = 8'he4 == io_state_in_11 ? 8'h37 : _GEN_5603; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5605 = 8'he5 == io_state_in_11 ? 8'h34 : _GEN_5604; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5606 = 8'he6 == io_state_in_11 ? 8'h31 : _GEN_5605; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5607 = 8'he7 == io_state_in_11 ? 8'h32 : _GEN_5606; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5608 = 8'he8 == io_state_in_11 ? 8'h23 : _GEN_5607; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5609 = 8'he9 == io_state_in_11 ? 8'h20 : _GEN_5608; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5610 = 8'hea == io_state_in_11 ? 8'h25 : _GEN_5609; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5611 = 8'heb == io_state_in_11 ? 8'h26 : _GEN_5610; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5612 = 8'hec == io_state_in_11 ? 8'h2f : _GEN_5611; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5613 = 8'hed == io_state_in_11 ? 8'h2c : _GEN_5612; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5614 = 8'hee == io_state_in_11 ? 8'h29 : _GEN_5613; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5615 = 8'hef == io_state_in_11 ? 8'h2a : _GEN_5614; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5616 = 8'hf0 == io_state_in_11 ? 8'hb : _GEN_5615; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5617 = 8'hf1 == io_state_in_11 ? 8'h8 : _GEN_5616; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5618 = 8'hf2 == io_state_in_11 ? 8'hd : _GEN_5617; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5619 = 8'hf3 == io_state_in_11 ? 8'he : _GEN_5618; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5620 = 8'hf4 == io_state_in_11 ? 8'h7 : _GEN_5619; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5621 = 8'hf5 == io_state_in_11 ? 8'h4 : _GEN_5620; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5622 = 8'hf6 == io_state_in_11 ? 8'h1 : _GEN_5621; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5623 = 8'hf7 == io_state_in_11 ? 8'h2 : _GEN_5622; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5624 = 8'hf8 == io_state_in_11 ? 8'h13 : _GEN_5623; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5625 = 8'hf9 == io_state_in_11 ? 8'h10 : _GEN_5624; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5626 = 8'hfa == io_state_in_11 ? 8'h15 : _GEN_5625; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5627 = 8'hfb == io_state_in_11 ? 8'h16 : _GEN_5626; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5628 = 8'hfc == io_state_in_11 ? 8'h1f : _GEN_5627; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5629 = 8'hfd == io_state_in_11 ? 8'h1c : _GEN_5628; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5630 = 8'hfe == io_state_in_11 ? 8'h19 : _GEN_5629; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5631 = 8'hff == io_state_in_11 ? 8'h1a : _GEN_5630; // @[MixColumns.scala 137:{77,77}]
  wire [7:0] _GEN_5633 = 8'h1 == io_state_in_8 ? 8'h3 : 8'h0; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5634 = 8'h2 == io_state_in_8 ? 8'h6 : _GEN_5633; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5635 = 8'h3 == io_state_in_8 ? 8'h5 : _GEN_5634; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5636 = 8'h4 == io_state_in_8 ? 8'hc : _GEN_5635; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5637 = 8'h5 == io_state_in_8 ? 8'hf : _GEN_5636; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5638 = 8'h6 == io_state_in_8 ? 8'ha : _GEN_5637; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5639 = 8'h7 == io_state_in_8 ? 8'h9 : _GEN_5638; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5640 = 8'h8 == io_state_in_8 ? 8'h18 : _GEN_5639; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5641 = 8'h9 == io_state_in_8 ? 8'h1b : _GEN_5640; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5642 = 8'ha == io_state_in_8 ? 8'h1e : _GEN_5641; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5643 = 8'hb == io_state_in_8 ? 8'h1d : _GEN_5642; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5644 = 8'hc == io_state_in_8 ? 8'h14 : _GEN_5643; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5645 = 8'hd == io_state_in_8 ? 8'h17 : _GEN_5644; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5646 = 8'he == io_state_in_8 ? 8'h12 : _GEN_5645; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5647 = 8'hf == io_state_in_8 ? 8'h11 : _GEN_5646; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5648 = 8'h10 == io_state_in_8 ? 8'h30 : _GEN_5647; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5649 = 8'h11 == io_state_in_8 ? 8'h33 : _GEN_5648; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5650 = 8'h12 == io_state_in_8 ? 8'h36 : _GEN_5649; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5651 = 8'h13 == io_state_in_8 ? 8'h35 : _GEN_5650; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5652 = 8'h14 == io_state_in_8 ? 8'h3c : _GEN_5651; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5653 = 8'h15 == io_state_in_8 ? 8'h3f : _GEN_5652; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5654 = 8'h16 == io_state_in_8 ? 8'h3a : _GEN_5653; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5655 = 8'h17 == io_state_in_8 ? 8'h39 : _GEN_5654; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5656 = 8'h18 == io_state_in_8 ? 8'h28 : _GEN_5655; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5657 = 8'h19 == io_state_in_8 ? 8'h2b : _GEN_5656; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5658 = 8'h1a == io_state_in_8 ? 8'h2e : _GEN_5657; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5659 = 8'h1b == io_state_in_8 ? 8'h2d : _GEN_5658; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5660 = 8'h1c == io_state_in_8 ? 8'h24 : _GEN_5659; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5661 = 8'h1d == io_state_in_8 ? 8'h27 : _GEN_5660; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5662 = 8'h1e == io_state_in_8 ? 8'h22 : _GEN_5661; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5663 = 8'h1f == io_state_in_8 ? 8'h21 : _GEN_5662; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5664 = 8'h20 == io_state_in_8 ? 8'h60 : _GEN_5663; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5665 = 8'h21 == io_state_in_8 ? 8'h63 : _GEN_5664; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5666 = 8'h22 == io_state_in_8 ? 8'h66 : _GEN_5665; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5667 = 8'h23 == io_state_in_8 ? 8'h65 : _GEN_5666; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5668 = 8'h24 == io_state_in_8 ? 8'h6c : _GEN_5667; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5669 = 8'h25 == io_state_in_8 ? 8'h6f : _GEN_5668; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5670 = 8'h26 == io_state_in_8 ? 8'h6a : _GEN_5669; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5671 = 8'h27 == io_state_in_8 ? 8'h69 : _GEN_5670; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5672 = 8'h28 == io_state_in_8 ? 8'h78 : _GEN_5671; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5673 = 8'h29 == io_state_in_8 ? 8'h7b : _GEN_5672; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5674 = 8'h2a == io_state_in_8 ? 8'h7e : _GEN_5673; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5675 = 8'h2b == io_state_in_8 ? 8'h7d : _GEN_5674; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5676 = 8'h2c == io_state_in_8 ? 8'h74 : _GEN_5675; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5677 = 8'h2d == io_state_in_8 ? 8'h77 : _GEN_5676; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5678 = 8'h2e == io_state_in_8 ? 8'h72 : _GEN_5677; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5679 = 8'h2f == io_state_in_8 ? 8'h71 : _GEN_5678; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5680 = 8'h30 == io_state_in_8 ? 8'h50 : _GEN_5679; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5681 = 8'h31 == io_state_in_8 ? 8'h53 : _GEN_5680; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5682 = 8'h32 == io_state_in_8 ? 8'h56 : _GEN_5681; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5683 = 8'h33 == io_state_in_8 ? 8'h55 : _GEN_5682; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5684 = 8'h34 == io_state_in_8 ? 8'h5c : _GEN_5683; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5685 = 8'h35 == io_state_in_8 ? 8'h5f : _GEN_5684; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5686 = 8'h36 == io_state_in_8 ? 8'h5a : _GEN_5685; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5687 = 8'h37 == io_state_in_8 ? 8'h59 : _GEN_5686; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5688 = 8'h38 == io_state_in_8 ? 8'h48 : _GEN_5687; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5689 = 8'h39 == io_state_in_8 ? 8'h4b : _GEN_5688; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5690 = 8'h3a == io_state_in_8 ? 8'h4e : _GEN_5689; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5691 = 8'h3b == io_state_in_8 ? 8'h4d : _GEN_5690; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5692 = 8'h3c == io_state_in_8 ? 8'h44 : _GEN_5691; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5693 = 8'h3d == io_state_in_8 ? 8'h47 : _GEN_5692; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5694 = 8'h3e == io_state_in_8 ? 8'h42 : _GEN_5693; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5695 = 8'h3f == io_state_in_8 ? 8'h41 : _GEN_5694; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5696 = 8'h40 == io_state_in_8 ? 8'hc0 : _GEN_5695; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5697 = 8'h41 == io_state_in_8 ? 8'hc3 : _GEN_5696; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5698 = 8'h42 == io_state_in_8 ? 8'hc6 : _GEN_5697; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5699 = 8'h43 == io_state_in_8 ? 8'hc5 : _GEN_5698; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5700 = 8'h44 == io_state_in_8 ? 8'hcc : _GEN_5699; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5701 = 8'h45 == io_state_in_8 ? 8'hcf : _GEN_5700; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5702 = 8'h46 == io_state_in_8 ? 8'hca : _GEN_5701; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5703 = 8'h47 == io_state_in_8 ? 8'hc9 : _GEN_5702; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5704 = 8'h48 == io_state_in_8 ? 8'hd8 : _GEN_5703; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5705 = 8'h49 == io_state_in_8 ? 8'hdb : _GEN_5704; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5706 = 8'h4a == io_state_in_8 ? 8'hde : _GEN_5705; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5707 = 8'h4b == io_state_in_8 ? 8'hdd : _GEN_5706; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5708 = 8'h4c == io_state_in_8 ? 8'hd4 : _GEN_5707; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5709 = 8'h4d == io_state_in_8 ? 8'hd7 : _GEN_5708; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5710 = 8'h4e == io_state_in_8 ? 8'hd2 : _GEN_5709; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5711 = 8'h4f == io_state_in_8 ? 8'hd1 : _GEN_5710; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5712 = 8'h50 == io_state_in_8 ? 8'hf0 : _GEN_5711; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5713 = 8'h51 == io_state_in_8 ? 8'hf3 : _GEN_5712; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5714 = 8'h52 == io_state_in_8 ? 8'hf6 : _GEN_5713; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5715 = 8'h53 == io_state_in_8 ? 8'hf5 : _GEN_5714; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5716 = 8'h54 == io_state_in_8 ? 8'hfc : _GEN_5715; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5717 = 8'h55 == io_state_in_8 ? 8'hff : _GEN_5716; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5718 = 8'h56 == io_state_in_8 ? 8'hfa : _GEN_5717; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5719 = 8'h57 == io_state_in_8 ? 8'hf9 : _GEN_5718; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5720 = 8'h58 == io_state_in_8 ? 8'he8 : _GEN_5719; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5721 = 8'h59 == io_state_in_8 ? 8'heb : _GEN_5720; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5722 = 8'h5a == io_state_in_8 ? 8'hee : _GEN_5721; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5723 = 8'h5b == io_state_in_8 ? 8'hed : _GEN_5722; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5724 = 8'h5c == io_state_in_8 ? 8'he4 : _GEN_5723; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5725 = 8'h5d == io_state_in_8 ? 8'he7 : _GEN_5724; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5726 = 8'h5e == io_state_in_8 ? 8'he2 : _GEN_5725; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5727 = 8'h5f == io_state_in_8 ? 8'he1 : _GEN_5726; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5728 = 8'h60 == io_state_in_8 ? 8'ha0 : _GEN_5727; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5729 = 8'h61 == io_state_in_8 ? 8'ha3 : _GEN_5728; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5730 = 8'h62 == io_state_in_8 ? 8'ha6 : _GEN_5729; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5731 = 8'h63 == io_state_in_8 ? 8'ha5 : _GEN_5730; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5732 = 8'h64 == io_state_in_8 ? 8'hac : _GEN_5731; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5733 = 8'h65 == io_state_in_8 ? 8'haf : _GEN_5732; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5734 = 8'h66 == io_state_in_8 ? 8'haa : _GEN_5733; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5735 = 8'h67 == io_state_in_8 ? 8'ha9 : _GEN_5734; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5736 = 8'h68 == io_state_in_8 ? 8'hb8 : _GEN_5735; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5737 = 8'h69 == io_state_in_8 ? 8'hbb : _GEN_5736; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5738 = 8'h6a == io_state_in_8 ? 8'hbe : _GEN_5737; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5739 = 8'h6b == io_state_in_8 ? 8'hbd : _GEN_5738; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5740 = 8'h6c == io_state_in_8 ? 8'hb4 : _GEN_5739; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5741 = 8'h6d == io_state_in_8 ? 8'hb7 : _GEN_5740; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5742 = 8'h6e == io_state_in_8 ? 8'hb2 : _GEN_5741; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5743 = 8'h6f == io_state_in_8 ? 8'hb1 : _GEN_5742; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5744 = 8'h70 == io_state_in_8 ? 8'h90 : _GEN_5743; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5745 = 8'h71 == io_state_in_8 ? 8'h93 : _GEN_5744; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5746 = 8'h72 == io_state_in_8 ? 8'h96 : _GEN_5745; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5747 = 8'h73 == io_state_in_8 ? 8'h95 : _GEN_5746; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5748 = 8'h74 == io_state_in_8 ? 8'h9c : _GEN_5747; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5749 = 8'h75 == io_state_in_8 ? 8'h9f : _GEN_5748; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5750 = 8'h76 == io_state_in_8 ? 8'h9a : _GEN_5749; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5751 = 8'h77 == io_state_in_8 ? 8'h99 : _GEN_5750; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5752 = 8'h78 == io_state_in_8 ? 8'h88 : _GEN_5751; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5753 = 8'h79 == io_state_in_8 ? 8'h8b : _GEN_5752; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5754 = 8'h7a == io_state_in_8 ? 8'h8e : _GEN_5753; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5755 = 8'h7b == io_state_in_8 ? 8'h8d : _GEN_5754; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5756 = 8'h7c == io_state_in_8 ? 8'h84 : _GEN_5755; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5757 = 8'h7d == io_state_in_8 ? 8'h87 : _GEN_5756; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5758 = 8'h7e == io_state_in_8 ? 8'h82 : _GEN_5757; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5759 = 8'h7f == io_state_in_8 ? 8'h81 : _GEN_5758; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5760 = 8'h80 == io_state_in_8 ? 8'h9b : _GEN_5759; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5761 = 8'h81 == io_state_in_8 ? 8'h98 : _GEN_5760; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5762 = 8'h82 == io_state_in_8 ? 8'h9d : _GEN_5761; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5763 = 8'h83 == io_state_in_8 ? 8'h9e : _GEN_5762; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5764 = 8'h84 == io_state_in_8 ? 8'h97 : _GEN_5763; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5765 = 8'h85 == io_state_in_8 ? 8'h94 : _GEN_5764; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5766 = 8'h86 == io_state_in_8 ? 8'h91 : _GEN_5765; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5767 = 8'h87 == io_state_in_8 ? 8'h92 : _GEN_5766; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5768 = 8'h88 == io_state_in_8 ? 8'h83 : _GEN_5767; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5769 = 8'h89 == io_state_in_8 ? 8'h80 : _GEN_5768; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5770 = 8'h8a == io_state_in_8 ? 8'h85 : _GEN_5769; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5771 = 8'h8b == io_state_in_8 ? 8'h86 : _GEN_5770; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5772 = 8'h8c == io_state_in_8 ? 8'h8f : _GEN_5771; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5773 = 8'h8d == io_state_in_8 ? 8'h8c : _GEN_5772; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5774 = 8'h8e == io_state_in_8 ? 8'h89 : _GEN_5773; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5775 = 8'h8f == io_state_in_8 ? 8'h8a : _GEN_5774; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5776 = 8'h90 == io_state_in_8 ? 8'hab : _GEN_5775; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5777 = 8'h91 == io_state_in_8 ? 8'ha8 : _GEN_5776; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5778 = 8'h92 == io_state_in_8 ? 8'had : _GEN_5777; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5779 = 8'h93 == io_state_in_8 ? 8'hae : _GEN_5778; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5780 = 8'h94 == io_state_in_8 ? 8'ha7 : _GEN_5779; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5781 = 8'h95 == io_state_in_8 ? 8'ha4 : _GEN_5780; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5782 = 8'h96 == io_state_in_8 ? 8'ha1 : _GEN_5781; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5783 = 8'h97 == io_state_in_8 ? 8'ha2 : _GEN_5782; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5784 = 8'h98 == io_state_in_8 ? 8'hb3 : _GEN_5783; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5785 = 8'h99 == io_state_in_8 ? 8'hb0 : _GEN_5784; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5786 = 8'h9a == io_state_in_8 ? 8'hb5 : _GEN_5785; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5787 = 8'h9b == io_state_in_8 ? 8'hb6 : _GEN_5786; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5788 = 8'h9c == io_state_in_8 ? 8'hbf : _GEN_5787; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5789 = 8'h9d == io_state_in_8 ? 8'hbc : _GEN_5788; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5790 = 8'h9e == io_state_in_8 ? 8'hb9 : _GEN_5789; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5791 = 8'h9f == io_state_in_8 ? 8'hba : _GEN_5790; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5792 = 8'ha0 == io_state_in_8 ? 8'hfb : _GEN_5791; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5793 = 8'ha1 == io_state_in_8 ? 8'hf8 : _GEN_5792; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5794 = 8'ha2 == io_state_in_8 ? 8'hfd : _GEN_5793; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5795 = 8'ha3 == io_state_in_8 ? 8'hfe : _GEN_5794; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5796 = 8'ha4 == io_state_in_8 ? 8'hf7 : _GEN_5795; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5797 = 8'ha5 == io_state_in_8 ? 8'hf4 : _GEN_5796; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5798 = 8'ha6 == io_state_in_8 ? 8'hf1 : _GEN_5797; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5799 = 8'ha7 == io_state_in_8 ? 8'hf2 : _GEN_5798; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5800 = 8'ha8 == io_state_in_8 ? 8'he3 : _GEN_5799; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5801 = 8'ha9 == io_state_in_8 ? 8'he0 : _GEN_5800; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5802 = 8'haa == io_state_in_8 ? 8'he5 : _GEN_5801; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5803 = 8'hab == io_state_in_8 ? 8'he6 : _GEN_5802; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5804 = 8'hac == io_state_in_8 ? 8'hef : _GEN_5803; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5805 = 8'had == io_state_in_8 ? 8'hec : _GEN_5804; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5806 = 8'hae == io_state_in_8 ? 8'he9 : _GEN_5805; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5807 = 8'haf == io_state_in_8 ? 8'hea : _GEN_5806; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5808 = 8'hb0 == io_state_in_8 ? 8'hcb : _GEN_5807; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5809 = 8'hb1 == io_state_in_8 ? 8'hc8 : _GEN_5808; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5810 = 8'hb2 == io_state_in_8 ? 8'hcd : _GEN_5809; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5811 = 8'hb3 == io_state_in_8 ? 8'hce : _GEN_5810; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5812 = 8'hb4 == io_state_in_8 ? 8'hc7 : _GEN_5811; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5813 = 8'hb5 == io_state_in_8 ? 8'hc4 : _GEN_5812; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5814 = 8'hb6 == io_state_in_8 ? 8'hc1 : _GEN_5813; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5815 = 8'hb7 == io_state_in_8 ? 8'hc2 : _GEN_5814; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5816 = 8'hb8 == io_state_in_8 ? 8'hd3 : _GEN_5815; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5817 = 8'hb9 == io_state_in_8 ? 8'hd0 : _GEN_5816; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5818 = 8'hba == io_state_in_8 ? 8'hd5 : _GEN_5817; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5819 = 8'hbb == io_state_in_8 ? 8'hd6 : _GEN_5818; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5820 = 8'hbc == io_state_in_8 ? 8'hdf : _GEN_5819; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5821 = 8'hbd == io_state_in_8 ? 8'hdc : _GEN_5820; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5822 = 8'hbe == io_state_in_8 ? 8'hd9 : _GEN_5821; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5823 = 8'hbf == io_state_in_8 ? 8'hda : _GEN_5822; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5824 = 8'hc0 == io_state_in_8 ? 8'h5b : _GEN_5823; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5825 = 8'hc1 == io_state_in_8 ? 8'h58 : _GEN_5824; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5826 = 8'hc2 == io_state_in_8 ? 8'h5d : _GEN_5825; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5827 = 8'hc3 == io_state_in_8 ? 8'h5e : _GEN_5826; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5828 = 8'hc4 == io_state_in_8 ? 8'h57 : _GEN_5827; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5829 = 8'hc5 == io_state_in_8 ? 8'h54 : _GEN_5828; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5830 = 8'hc6 == io_state_in_8 ? 8'h51 : _GEN_5829; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5831 = 8'hc7 == io_state_in_8 ? 8'h52 : _GEN_5830; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5832 = 8'hc8 == io_state_in_8 ? 8'h43 : _GEN_5831; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5833 = 8'hc9 == io_state_in_8 ? 8'h40 : _GEN_5832; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5834 = 8'hca == io_state_in_8 ? 8'h45 : _GEN_5833; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5835 = 8'hcb == io_state_in_8 ? 8'h46 : _GEN_5834; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5836 = 8'hcc == io_state_in_8 ? 8'h4f : _GEN_5835; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5837 = 8'hcd == io_state_in_8 ? 8'h4c : _GEN_5836; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5838 = 8'hce == io_state_in_8 ? 8'h49 : _GEN_5837; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5839 = 8'hcf == io_state_in_8 ? 8'h4a : _GEN_5838; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5840 = 8'hd0 == io_state_in_8 ? 8'h6b : _GEN_5839; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5841 = 8'hd1 == io_state_in_8 ? 8'h68 : _GEN_5840; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5842 = 8'hd2 == io_state_in_8 ? 8'h6d : _GEN_5841; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5843 = 8'hd3 == io_state_in_8 ? 8'h6e : _GEN_5842; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5844 = 8'hd4 == io_state_in_8 ? 8'h67 : _GEN_5843; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5845 = 8'hd5 == io_state_in_8 ? 8'h64 : _GEN_5844; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5846 = 8'hd6 == io_state_in_8 ? 8'h61 : _GEN_5845; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5847 = 8'hd7 == io_state_in_8 ? 8'h62 : _GEN_5846; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5848 = 8'hd8 == io_state_in_8 ? 8'h73 : _GEN_5847; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5849 = 8'hd9 == io_state_in_8 ? 8'h70 : _GEN_5848; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5850 = 8'hda == io_state_in_8 ? 8'h75 : _GEN_5849; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5851 = 8'hdb == io_state_in_8 ? 8'h76 : _GEN_5850; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5852 = 8'hdc == io_state_in_8 ? 8'h7f : _GEN_5851; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5853 = 8'hdd == io_state_in_8 ? 8'h7c : _GEN_5852; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5854 = 8'hde == io_state_in_8 ? 8'h79 : _GEN_5853; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5855 = 8'hdf == io_state_in_8 ? 8'h7a : _GEN_5854; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5856 = 8'he0 == io_state_in_8 ? 8'h3b : _GEN_5855; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5857 = 8'he1 == io_state_in_8 ? 8'h38 : _GEN_5856; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5858 = 8'he2 == io_state_in_8 ? 8'h3d : _GEN_5857; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5859 = 8'he3 == io_state_in_8 ? 8'h3e : _GEN_5858; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5860 = 8'he4 == io_state_in_8 ? 8'h37 : _GEN_5859; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5861 = 8'he5 == io_state_in_8 ? 8'h34 : _GEN_5860; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5862 = 8'he6 == io_state_in_8 ? 8'h31 : _GEN_5861; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5863 = 8'he7 == io_state_in_8 ? 8'h32 : _GEN_5862; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5864 = 8'he8 == io_state_in_8 ? 8'h23 : _GEN_5863; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5865 = 8'he9 == io_state_in_8 ? 8'h20 : _GEN_5864; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5866 = 8'hea == io_state_in_8 ? 8'h25 : _GEN_5865; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5867 = 8'heb == io_state_in_8 ? 8'h26 : _GEN_5866; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5868 = 8'hec == io_state_in_8 ? 8'h2f : _GEN_5867; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5869 = 8'hed == io_state_in_8 ? 8'h2c : _GEN_5868; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5870 = 8'hee == io_state_in_8 ? 8'h29 : _GEN_5869; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5871 = 8'hef == io_state_in_8 ? 8'h2a : _GEN_5870; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5872 = 8'hf0 == io_state_in_8 ? 8'hb : _GEN_5871; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5873 = 8'hf1 == io_state_in_8 ? 8'h8 : _GEN_5872; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5874 = 8'hf2 == io_state_in_8 ? 8'hd : _GEN_5873; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5875 = 8'hf3 == io_state_in_8 ? 8'he : _GEN_5874; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5876 = 8'hf4 == io_state_in_8 ? 8'h7 : _GEN_5875; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5877 = 8'hf5 == io_state_in_8 ? 8'h4 : _GEN_5876; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5878 = 8'hf6 == io_state_in_8 ? 8'h1 : _GEN_5877; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5879 = 8'hf7 == io_state_in_8 ? 8'h2 : _GEN_5878; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5880 = 8'hf8 == io_state_in_8 ? 8'h13 : _GEN_5879; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5881 = 8'hf9 == io_state_in_8 ? 8'h10 : _GEN_5880; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5882 = 8'hfa == io_state_in_8 ? 8'h15 : _GEN_5881; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5883 = 8'hfb == io_state_in_8 ? 8'h16 : _GEN_5882; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5884 = 8'hfc == io_state_in_8 ? 8'h1f : _GEN_5883; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5885 = 8'hfd == io_state_in_8 ? 8'h1c : _GEN_5884; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5886 = 8'hfe == io_state_in_8 ? 8'h19 : _GEN_5885; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _GEN_5887 = 8'hff == io_state_in_8 ? 8'h1a : _GEN_5886; // @[MixColumns.scala 138:{42,42}]
  wire [7:0] _tmp_state_11_T = _GEN_5887 ^ io_state_in_9; // @[MixColumns.scala 138:42]
  wire [7:0] _tmp_state_11_T_1 = _tmp_state_11_T ^ io_state_in_10; // @[MixColumns.scala 138:59]
  wire [7:0] _GEN_5889 = 8'h1 == io_state_in_11 ? 8'h2 : 8'h0; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5890 = 8'h2 == io_state_in_11 ? 8'h4 : _GEN_5889; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5891 = 8'h3 == io_state_in_11 ? 8'h6 : _GEN_5890; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5892 = 8'h4 == io_state_in_11 ? 8'h8 : _GEN_5891; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5893 = 8'h5 == io_state_in_11 ? 8'ha : _GEN_5892; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5894 = 8'h6 == io_state_in_11 ? 8'hc : _GEN_5893; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5895 = 8'h7 == io_state_in_11 ? 8'he : _GEN_5894; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5896 = 8'h8 == io_state_in_11 ? 8'h10 : _GEN_5895; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5897 = 8'h9 == io_state_in_11 ? 8'h12 : _GEN_5896; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5898 = 8'ha == io_state_in_11 ? 8'h14 : _GEN_5897; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5899 = 8'hb == io_state_in_11 ? 8'h16 : _GEN_5898; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5900 = 8'hc == io_state_in_11 ? 8'h18 : _GEN_5899; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5901 = 8'hd == io_state_in_11 ? 8'h1a : _GEN_5900; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5902 = 8'he == io_state_in_11 ? 8'h1c : _GEN_5901; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5903 = 8'hf == io_state_in_11 ? 8'h1e : _GEN_5902; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5904 = 8'h10 == io_state_in_11 ? 8'h20 : _GEN_5903; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5905 = 8'h11 == io_state_in_11 ? 8'h22 : _GEN_5904; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5906 = 8'h12 == io_state_in_11 ? 8'h24 : _GEN_5905; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5907 = 8'h13 == io_state_in_11 ? 8'h26 : _GEN_5906; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5908 = 8'h14 == io_state_in_11 ? 8'h28 : _GEN_5907; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5909 = 8'h15 == io_state_in_11 ? 8'h2a : _GEN_5908; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5910 = 8'h16 == io_state_in_11 ? 8'h2c : _GEN_5909; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5911 = 8'h17 == io_state_in_11 ? 8'h2e : _GEN_5910; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5912 = 8'h18 == io_state_in_11 ? 8'h30 : _GEN_5911; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5913 = 8'h19 == io_state_in_11 ? 8'h32 : _GEN_5912; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5914 = 8'h1a == io_state_in_11 ? 8'h34 : _GEN_5913; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5915 = 8'h1b == io_state_in_11 ? 8'h36 : _GEN_5914; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5916 = 8'h1c == io_state_in_11 ? 8'h38 : _GEN_5915; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5917 = 8'h1d == io_state_in_11 ? 8'h3a : _GEN_5916; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5918 = 8'h1e == io_state_in_11 ? 8'h3c : _GEN_5917; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5919 = 8'h1f == io_state_in_11 ? 8'h3e : _GEN_5918; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5920 = 8'h20 == io_state_in_11 ? 8'h40 : _GEN_5919; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5921 = 8'h21 == io_state_in_11 ? 8'h42 : _GEN_5920; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5922 = 8'h22 == io_state_in_11 ? 8'h44 : _GEN_5921; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5923 = 8'h23 == io_state_in_11 ? 8'h46 : _GEN_5922; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5924 = 8'h24 == io_state_in_11 ? 8'h48 : _GEN_5923; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5925 = 8'h25 == io_state_in_11 ? 8'h4a : _GEN_5924; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5926 = 8'h26 == io_state_in_11 ? 8'h4c : _GEN_5925; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5927 = 8'h27 == io_state_in_11 ? 8'h4e : _GEN_5926; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5928 = 8'h28 == io_state_in_11 ? 8'h50 : _GEN_5927; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5929 = 8'h29 == io_state_in_11 ? 8'h52 : _GEN_5928; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5930 = 8'h2a == io_state_in_11 ? 8'h54 : _GEN_5929; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5931 = 8'h2b == io_state_in_11 ? 8'h56 : _GEN_5930; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5932 = 8'h2c == io_state_in_11 ? 8'h58 : _GEN_5931; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5933 = 8'h2d == io_state_in_11 ? 8'h5a : _GEN_5932; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5934 = 8'h2e == io_state_in_11 ? 8'h5c : _GEN_5933; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5935 = 8'h2f == io_state_in_11 ? 8'h5e : _GEN_5934; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5936 = 8'h30 == io_state_in_11 ? 8'h60 : _GEN_5935; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5937 = 8'h31 == io_state_in_11 ? 8'h62 : _GEN_5936; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5938 = 8'h32 == io_state_in_11 ? 8'h64 : _GEN_5937; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5939 = 8'h33 == io_state_in_11 ? 8'h66 : _GEN_5938; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5940 = 8'h34 == io_state_in_11 ? 8'h68 : _GEN_5939; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5941 = 8'h35 == io_state_in_11 ? 8'h6a : _GEN_5940; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5942 = 8'h36 == io_state_in_11 ? 8'h6c : _GEN_5941; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5943 = 8'h37 == io_state_in_11 ? 8'h6e : _GEN_5942; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5944 = 8'h38 == io_state_in_11 ? 8'h70 : _GEN_5943; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5945 = 8'h39 == io_state_in_11 ? 8'h72 : _GEN_5944; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5946 = 8'h3a == io_state_in_11 ? 8'h74 : _GEN_5945; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5947 = 8'h3b == io_state_in_11 ? 8'h76 : _GEN_5946; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5948 = 8'h3c == io_state_in_11 ? 8'h78 : _GEN_5947; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5949 = 8'h3d == io_state_in_11 ? 8'h7a : _GEN_5948; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5950 = 8'h3e == io_state_in_11 ? 8'h7c : _GEN_5949; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5951 = 8'h3f == io_state_in_11 ? 8'h7e : _GEN_5950; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5952 = 8'h40 == io_state_in_11 ? 8'h80 : _GEN_5951; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5953 = 8'h41 == io_state_in_11 ? 8'h82 : _GEN_5952; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5954 = 8'h42 == io_state_in_11 ? 8'h84 : _GEN_5953; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5955 = 8'h43 == io_state_in_11 ? 8'h86 : _GEN_5954; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5956 = 8'h44 == io_state_in_11 ? 8'h88 : _GEN_5955; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5957 = 8'h45 == io_state_in_11 ? 8'h8a : _GEN_5956; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5958 = 8'h46 == io_state_in_11 ? 8'h8c : _GEN_5957; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5959 = 8'h47 == io_state_in_11 ? 8'h8e : _GEN_5958; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5960 = 8'h48 == io_state_in_11 ? 8'h90 : _GEN_5959; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5961 = 8'h49 == io_state_in_11 ? 8'h92 : _GEN_5960; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5962 = 8'h4a == io_state_in_11 ? 8'h94 : _GEN_5961; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5963 = 8'h4b == io_state_in_11 ? 8'h96 : _GEN_5962; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5964 = 8'h4c == io_state_in_11 ? 8'h98 : _GEN_5963; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5965 = 8'h4d == io_state_in_11 ? 8'h9a : _GEN_5964; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5966 = 8'h4e == io_state_in_11 ? 8'h9c : _GEN_5965; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5967 = 8'h4f == io_state_in_11 ? 8'h9e : _GEN_5966; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5968 = 8'h50 == io_state_in_11 ? 8'ha0 : _GEN_5967; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5969 = 8'h51 == io_state_in_11 ? 8'ha2 : _GEN_5968; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5970 = 8'h52 == io_state_in_11 ? 8'ha4 : _GEN_5969; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5971 = 8'h53 == io_state_in_11 ? 8'ha6 : _GEN_5970; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5972 = 8'h54 == io_state_in_11 ? 8'ha8 : _GEN_5971; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5973 = 8'h55 == io_state_in_11 ? 8'haa : _GEN_5972; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5974 = 8'h56 == io_state_in_11 ? 8'hac : _GEN_5973; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5975 = 8'h57 == io_state_in_11 ? 8'hae : _GEN_5974; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5976 = 8'h58 == io_state_in_11 ? 8'hb0 : _GEN_5975; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5977 = 8'h59 == io_state_in_11 ? 8'hb2 : _GEN_5976; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5978 = 8'h5a == io_state_in_11 ? 8'hb4 : _GEN_5977; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5979 = 8'h5b == io_state_in_11 ? 8'hb6 : _GEN_5978; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5980 = 8'h5c == io_state_in_11 ? 8'hb8 : _GEN_5979; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5981 = 8'h5d == io_state_in_11 ? 8'hba : _GEN_5980; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5982 = 8'h5e == io_state_in_11 ? 8'hbc : _GEN_5981; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5983 = 8'h5f == io_state_in_11 ? 8'hbe : _GEN_5982; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5984 = 8'h60 == io_state_in_11 ? 8'hc0 : _GEN_5983; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5985 = 8'h61 == io_state_in_11 ? 8'hc2 : _GEN_5984; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5986 = 8'h62 == io_state_in_11 ? 8'hc4 : _GEN_5985; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5987 = 8'h63 == io_state_in_11 ? 8'hc6 : _GEN_5986; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5988 = 8'h64 == io_state_in_11 ? 8'hc8 : _GEN_5987; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5989 = 8'h65 == io_state_in_11 ? 8'hca : _GEN_5988; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5990 = 8'h66 == io_state_in_11 ? 8'hcc : _GEN_5989; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5991 = 8'h67 == io_state_in_11 ? 8'hce : _GEN_5990; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5992 = 8'h68 == io_state_in_11 ? 8'hd0 : _GEN_5991; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5993 = 8'h69 == io_state_in_11 ? 8'hd2 : _GEN_5992; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5994 = 8'h6a == io_state_in_11 ? 8'hd4 : _GEN_5993; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5995 = 8'h6b == io_state_in_11 ? 8'hd6 : _GEN_5994; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5996 = 8'h6c == io_state_in_11 ? 8'hd8 : _GEN_5995; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5997 = 8'h6d == io_state_in_11 ? 8'hda : _GEN_5996; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5998 = 8'h6e == io_state_in_11 ? 8'hdc : _GEN_5997; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_5999 = 8'h6f == io_state_in_11 ? 8'hde : _GEN_5998; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6000 = 8'h70 == io_state_in_11 ? 8'he0 : _GEN_5999; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6001 = 8'h71 == io_state_in_11 ? 8'he2 : _GEN_6000; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6002 = 8'h72 == io_state_in_11 ? 8'he4 : _GEN_6001; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6003 = 8'h73 == io_state_in_11 ? 8'he6 : _GEN_6002; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6004 = 8'h74 == io_state_in_11 ? 8'he8 : _GEN_6003; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6005 = 8'h75 == io_state_in_11 ? 8'hea : _GEN_6004; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6006 = 8'h76 == io_state_in_11 ? 8'hec : _GEN_6005; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6007 = 8'h77 == io_state_in_11 ? 8'hee : _GEN_6006; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6008 = 8'h78 == io_state_in_11 ? 8'hf0 : _GEN_6007; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6009 = 8'h79 == io_state_in_11 ? 8'hf2 : _GEN_6008; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6010 = 8'h7a == io_state_in_11 ? 8'hf4 : _GEN_6009; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6011 = 8'h7b == io_state_in_11 ? 8'hf6 : _GEN_6010; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6012 = 8'h7c == io_state_in_11 ? 8'hf8 : _GEN_6011; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6013 = 8'h7d == io_state_in_11 ? 8'hfa : _GEN_6012; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6014 = 8'h7e == io_state_in_11 ? 8'hfc : _GEN_6013; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6015 = 8'h7f == io_state_in_11 ? 8'hfe : _GEN_6014; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6016 = 8'h80 == io_state_in_11 ? 8'h1b : _GEN_6015; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6017 = 8'h81 == io_state_in_11 ? 8'h19 : _GEN_6016; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6018 = 8'h82 == io_state_in_11 ? 8'h1f : _GEN_6017; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6019 = 8'h83 == io_state_in_11 ? 8'h1d : _GEN_6018; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6020 = 8'h84 == io_state_in_11 ? 8'h13 : _GEN_6019; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6021 = 8'h85 == io_state_in_11 ? 8'h11 : _GEN_6020; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6022 = 8'h86 == io_state_in_11 ? 8'h17 : _GEN_6021; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6023 = 8'h87 == io_state_in_11 ? 8'h15 : _GEN_6022; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6024 = 8'h88 == io_state_in_11 ? 8'hb : _GEN_6023; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6025 = 8'h89 == io_state_in_11 ? 8'h9 : _GEN_6024; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6026 = 8'h8a == io_state_in_11 ? 8'hf : _GEN_6025; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6027 = 8'h8b == io_state_in_11 ? 8'hd : _GEN_6026; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6028 = 8'h8c == io_state_in_11 ? 8'h3 : _GEN_6027; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6029 = 8'h8d == io_state_in_11 ? 8'h1 : _GEN_6028; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6030 = 8'h8e == io_state_in_11 ? 8'h7 : _GEN_6029; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6031 = 8'h8f == io_state_in_11 ? 8'h5 : _GEN_6030; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6032 = 8'h90 == io_state_in_11 ? 8'h3b : _GEN_6031; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6033 = 8'h91 == io_state_in_11 ? 8'h39 : _GEN_6032; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6034 = 8'h92 == io_state_in_11 ? 8'h3f : _GEN_6033; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6035 = 8'h93 == io_state_in_11 ? 8'h3d : _GEN_6034; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6036 = 8'h94 == io_state_in_11 ? 8'h33 : _GEN_6035; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6037 = 8'h95 == io_state_in_11 ? 8'h31 : _GEN_6036; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6038 = 8'h96 == io_state_in_11 ? 8'h37 : _GEN_6037; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6039 = 8'h97 == io_state_in_11 ? 8'h35 : _GEN_6038; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6040 = 8'h98 == io_state_in_11 ? 8'h2b : _GEN_6039; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6041 = 8'h99 == io_state_in_11 ? 8'h29 : _GEN_6040; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6042 = 8'h9a == io_state_in_11 ? 8'h2f : _GEN_6041; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6043 = 8'h9b == io_state_in_11 ? 8'h2d : _GEN_6042; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6044 = 8'h9c == io_state_in_11 ? 8'h23 : _GEN_6043; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6045 = 8'h9d == io_state_in_11 ? 8'h21 : _GEN_6044; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6046 = 8'h9e == io_state_in_11 ? 8'h27 : _GEN_6045; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6047 = 8'h9f == io_state_in_11 ? 8'h25 : _GEN_6046; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6048 = 8'ha0 == io_state_in_11 ? 8'h5b : _GEN_6047; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6049 = 8'ha1 == io_state_in_11 ? 8'h59 : _GEN_6048; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6050 = 8'ha2 == io_state_in_11 ? 8'h5f : _GEN_6049; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6051 = 8'ha3 == io_state_in_11 ? 8'h5d : _GEN_6050; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6052 = 8'ha4 == io_state_in_11 ? 8'h53 : _GEN_6051; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6053 = 8'ha5 == io_state_in_11 ? 8'h51 : _GEN_6052; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6054 = 8'ha6 == io_state_in_11 ? 8'h57 : _GEN_6053; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6055 = 8'ha7 == io_state_in_11 ? 8'h55 : _GEN_6054; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6056 = 8'ha8 == io_state_in_11 ? 8'h4b : _GEN_6055; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6057 = 8'ha9 == io_state_in_11 ? 8'h49 : _GEN_6056; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6058 = 8'haa == io_state_in_11 ? 8'h4f : _GEN_6057; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6059 = 8'hab == io_state_in_11 ? 8'h4d : _GEN_6058; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6060 = 8'hac == io_state_in_11 ? 8'h43 : _GEN_6059; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6061 = 8'had == io_state_in_11 ? 8'h41 : _GEN_6060; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6062 = 8'hae == io_state_in_11 ? 8'h47 : _GEN_6061; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6063 = 8'haf == io_state_in_11 ? 8'h45 : _GEN_6062; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6064 = 8'hb0 == io_state_in_11 ? 8'h7b : _GEN_6063; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6065 = 8'hb1 == io_state_in_11 ? 8'h79 : _GEN_6064; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6066 = 8'hb2 == io_state_in_11 ? 8'h7f : _GEN_6065; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6067 = 8'hb3 == io_state_in_11 ? 8'h7d : _GEN_6066; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6068 = 8'hb4 == io_state_in_11 ? 8'h73 : _GEN_6067; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6069 = 8'hb5 == io_state_in_11 ? 8'h71 : _GEN_6068; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6070 = 8'hb6 == io_state_in_11 ? 8'h77 : _GEN_6069; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6071 = 8'hb7 == io_state_in_11 ? 8'h75 : _GEN_6070; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6072 = 8'hb8 == io_state_in_11 ? 8'h6b : _GEN_6071; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6073 = 8'hb9 == io_state_in_11 ? 8'h69 : _GEN_6072; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6074 = 8'hba == io_state_in_11 ? 8'h6f : _GEN_6073; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6075 = 8'hbb == io_state_in_11 ? 8'h6d : _GEN_6074; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6076 = 8'hbc == io_state_in_11 ? 8'h63 : _GEN_6075; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6077 = 8'hbd == io_state_in_11 ? 8'h61 : _GEN_6076; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6078 = 8'hbe == io_state_in_11 ? 8'h67 : _GEN_6077; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6079 = 8'hbf == io_state_in_11 ? 8'h65 : _GEN_6078; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6080 = 8'hc0 == io_state_in_11 ? 8'h9b : _GEN_6079; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6081 = 8'hc1 == io_state_in_11 ? 8'h99 : _GEN_6080; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6082 = 8'hc2 == io_state_in_11 ? 8'h9f : _GEN_6081; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6083 = 8'hc3 == io_state_in_11 ? 8'h9d : _GEN_6082; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6084 = 8'hc4 == io_state_in_11 ? 8'h93 : _GEN_6083; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6085 = 8'hc5 == io_state_in_11 ? 8'h91 : _GEN_6084; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6086 = 8'hc6 == io_state_in_11 ? 8'h97 : _GEN_6085; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6087 = 8'hc7 == io_state_in_11 ? 8'h95 : _GEN_6086; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6088 = 8'hc8 == io_state_in_11 ? 8'h8b : _GEN_6087; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6089 = 8'hc9 == io_state_in_11 ? 8'h89 : _GEN_6088; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6090 = 8'hca == io_state_in_11 ? 8'h8f : _GEN_6089; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6091 = 8'hcb == io_state_in_11 ? 8'h8d : _GEN_6090; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6092 = 8'hcc == io_state_in_11 ? 8'h83 : _GEN_6091; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6093 = 8'hcd == io_state_in_11 ? 8'h81 : _GEN_6092; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6094 = 8'hce == io_state_in_11 ? 8'h87 : _GEN_6093; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6095 = 8'hcf == io_state_in_11 ? 8'h85 : _GEN_6094; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6096 = 8'hd0 == io_state_in_11 ? 8'hbb : _GEN_6095; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6097 = 8'hd1 == io_state_in_11 ? 8'hb9 : _GEN_6096; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6098 = 8'hd2 == io_state_in_11 ? 8'hbf : _GEN_6097; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6099 = 8'hd3 == io_state_in_11 ? 8'hbd : _GEN_6098; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6100 = 8'hd4 == io_state_in_11 ? 8'hb3 : _GEN_6099; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6101 = 8'hd5 == io_state_in_11 ? 8'hb1 : _GEN_6100; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6102 = 8'hd6 == io_state_in_11 ? 8'hb7 : _GEN_6101; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6103 = 8'hd7 == io_state_in_11 ? 8'hb5 : _GEN_6102; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6104 = 8'hd8 == io_state_in_11 ? 8'hab : _GEN_6103; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6105 = 8'hd9 == io_state_in_11 ? 8'ha9 : _GEN_6104; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6106 = 8'hda == io_state_in_11 ? 8'haf : _GEN_6105; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6107 = 8'hdb == io_state_in_11 ? 8'had : _GEN_6106; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6108 = 8'hdc == io_state_in_11 ? 8'ha3 : _GEN_6107; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6109 = 8'hdd == io_state_in_11 ? 8'ha1 : _GEN_6108; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6110 = 8'hde == io_state_in_11 ? 8'ha7 : _GEN_6109; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6111 = 8'hdf == io_state_in_11 ? 8'ha5 : _GEN_6110; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6112 = 8'he0 == io_state_in_11 ? 8'hdb : _GEN_6111; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6113 = 8'he1 == io_state_in_11 ? 8'hd9 : _GEN_6112; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6114 = 8'he2 == io_state_in_11 ? 8'hdf : _GEN_6113; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6115 = 8'he3 == io_state_in_11 ? 8'hdd : _GEN_6114; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6116 = 8'he4 == io_state_in_11 ? 8'hd3 : _GEN_6115; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6117 = 8'he5 == io_state_in_11 ? 8'hd1 : _GEN_6116; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6118 = 8'he6 == io_state_in_11 ? 8'hd7 : _GEN_6117; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6119 = 8'he7 == io_state_in_11 ? 8'hd5 : _GEN_6118; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6120 = 8'he8 == io_state_in_11 ? 8'hcb : _GEN_6119; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6121 = 8'he9 == io_state_in_11 ? 8'hc9 : _GEN_6120; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6122 = 8'hea == io_state_in_11 ? 8'hcf : _GEN_6121; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6123 = 8'heb == io_state_in_11 ? 8'hcd : _GEN_6122; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6124 = 8'hec == io_state_in_11 ? 8'hc3 : _GEN_6123; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6125 = 8'hed == io_state_in_11 ? 8'hc1 : _GEN_6124; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6126 = 8'hee == io_state_in_11 ? 8'hc7 : _GEN_6125; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6127 = 8'hef == io_state_in_11 ? 8'hc5 : _GEN_6126; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6128 = 8'hf0 == io_state_in_11 ? 8'hfb : _GEN_6127; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6129 = 8'hf1 == io_state_in_11 ? 8'hf9 : _GEN_6128; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6130 = 8'hf2 == io_state_in_11 ? 8'hff : _GEN_6129; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6131 = 8'hf3 == io_state_in_11 ? 8'hfd : _GEN_6130; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6132 = 8'hf4 == io_state_in_11 ? 8'hf3 : _GEN_6131; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6133 = 8'hf5 == io_state_in_11 ? 8'hf1 : _GEN_6132; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6134 = 8'hf6 == io_state_in_11 ? 8'hf7 : _GEN_6133; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6135 = 8'hf7 == io_state_in_11 ? 8'hf5 : _GEN_6134; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6136 = 8'hf8 == io_state_in_11 ? 8'heb : _GEN_6135; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6137 = 8'hf9 == io_state_in_11 ? 8'he9 : _GEN_6136; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6138 = 8'hfa == io_state_in_11 ? 8'hef : _GEN_6137; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6139 = 8'hfb == io_state_in_11 ? 8'hed : _GEN_6138; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6140 = 8'hfc == io_state_in_11 ? 8'he3 : _GEN_6139; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6141 = 8'hfd == io_state_in_11 ? 8'he1 : _GEN_6140; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6142 = 8'hfe == io_state_in_11 ? 8'he7 : _GEN_6141; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6143 = 8'hff == io_state_in_11 ? 8'he5 : _GEN_6142; // @[MixColumns.scala 138:{77,77}]
  wire [7:0] _GEN_6145 = 8'h1 == io_state_in_12 ? 8'h2 : 8'h0; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6146 = 8'h2 == io_state_in_12 ? 8'h4 : _GEN_6145; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6147 = 8'h3 == io_state_in_12 ? 8'h6 : _GEN_6146; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6148 = 8'h4 == io_state_in_12 ? 8'h8 : _GEN_6147; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6149 = 8'h5 == io_state_in_12 ? 8'ha : _GEN_6148; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6150 = 8'h6 == io_state_in_12 ? 8'hc : _GEN_6149; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6151 = 8'h7 == io_state_in_12 ? 8'he : _GEN_6150; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6152 = 8'h8 == io_state_in_12 ? 8'h10 : _GEN_6151; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6153 = 8'h9 == io_state_in_12 ? 8'h12 : _GEN_6152; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6154 = 8'ha == io_state_in_12 ? 8'h14 : _GEN_6153; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6155 = 8'hb == io_state_in_12 ? 8'h16 : _GEN_6154; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6156 = 8'hc == io_state_in_12 ? 8'h18 : _GEN_6155; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6157 = 8'hd == io_state_in_12 ? 8'h1a : _GEN_6156; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6158 = 8'he == io_state_in_12 ? 8'h1c : _GEN_6157; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6159 = 8'hf == io_state_in_12 ? 8'h1e : _GEN_6158; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6160 = 8'h10 == io_state_in_12 ? 8'h20 : _GEN_6159; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6161 = 8'h11 == io_state_in_12 ? 8'h22 : _GEN_6160; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6162 = 8'h12 == io_state_in_12 ? 8'h24 : _GEN_6161; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6163 = 8'h13 == io_state_in_12 ? 8'h26 : _GEN_6162; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6164 = 8'h14 == io_state_in_12 ? 8'h28 : _GEN_6163; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6165 = 8'h15 == io_state_in_12 ? 8'h2a : _GEN_6164; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6166 = 8'h16 == io_state_in_12 ? 8'h2c : _GEN_6165; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6167 = 8'h17 == io_state_in_12 ? 8'h2e : _GEN_6166; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6168 = 8'h18 == io_state_in_12 ? 8'h30 : _GEN_6167; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6169 = 8'h19 == io_state_in_12 ? 8'h32 : _GEN_6168; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6170 = 8'h1a == io_state_in_12 ? 8'h34 : _GEN_6169; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6171 = 8'h1b == io_state_in_12 ? 8'h36 : _GEN_6170; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6172 = 8'h1c == io_state_in_12 ? 8'h38 : _GEN_6171; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6173 = 8'h1d == io_state_in_12 ? 8'h3a : _GEN_6172; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6174 = 8'h1e == io_state_in_12 ? 8'h3c : _GEN_6173; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6175 = 8'h1f == io_state_in_12 ? 8'h3e : _GEN_6174; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6176 = 8'h20 == io_state_in_12 ? 8'h40 : _GEN_6175; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6177 = 8'h21 == io_state_in_12 ? 8'h42 : _GEN_6176; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6178 = 8'h22 == io_state_in_12 ? 8'h44 : _GEN_6177; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6179 = 8'h23 == io_state_in_12 ? 8'h46 : _GEN_6178; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6180 = 8'h24 == io_state_in_12 ? 8'h48 : _GEN_6179; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6181 = 8'h25 == io_state_in_12 ? 8'h4a : _GEN_6180; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6182 = 8'h26 == io_state_in_12 ? 8'h4c : _GEN_6181; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6183 = 8'h27 == io_state_in_12 ? 8'h4e : _GEN_6182; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6184 = 8'h28 == io_state_in_12 ? 8'h50 : _GEN_6183; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6185 = 8'h29 == io_state_in_12 ? 8'h52 : _GEN_6184; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6186 = 8'h2a == io_state_in_12 ? 8'h54 : _GEN_6185; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6187 = 8'h2b == io_state_in_12 ? 8'h56 : _GEN_6186; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6188 = 8'h2c == io_state_in_12 ? 8'h58 : _GEN_6187; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6189 = 8'h2d == io_state_in_12 ? 8'h5a : _GEN_6188; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6190 = 8'h2e == io_state_in_12 ? 8'h5c : _GEN_6189; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6191 = 8'h2f == io_state_in_12 ? 8'h5e : _GEN_6190; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6192 = 8'h30 == io_state_in_12 ? 8'h60 : _GEN_6191; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6193 = 8'h31 == io_state_in_12 ? 8'h62 : _GEN_6192; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6194 = 8'h32 == io_state_in_12 ? 8'h64 : _GEN_6193; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6195 = 8'h33 == io_state_in_12 ? 8'h66 : _GEN_6194; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6196 = 8'h34 == io_state_in_12 ? 8'h68 : _GEN_6195; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6197 = 8'h35 == io_state_in_12 ? 8'h6a : _GEN_6196; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6198 = 8'h36 == io_state_in_12 ? 8'h6c : _GEN_6197; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6199 = 8'h37 == io_state_in_12 ? 8'h6e : _GEN_6198; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6200 = 8'h38 == io_state_in_12 ? 8'h70 : _GEN_6199; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6201 = 8'h39 == io_state_in_12 ? 8'h72 : _GEN_6200; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6202 = 8'h3a == io_state_in_12 ? 8'h74 : _GEN_6201; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6203 = 8'h3b == io_state_in_12 ? 8'h76 : _GEN_6202; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6204 = 8'h3c == io_state_in_12 ? 8'h78 : _GEN_6203; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6205 = 8'h3d == io_state_in_12 ? 8'h7a : _GEN_6204; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6206 = 8'h3e == io_state_in_12 ? 8'h7c : _GEN_6205; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6207 = 8'h3f == io_state_in_12 ? 8'h7e : _GEN_6206; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6208 = 8'h40 == io_state_in_12 ? 8'h80 : _GEN_6207; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6209 = 8'h41 == io_state_in_12 ? 8'h82 : _GEN_6208; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6210 = 8'h42 == io_state_in_12 ? 8'h84 : _GEN_6209; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6211 = 8'h43 == io_state_in_12 ? 8'h86 : _GEN_6210; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6212 = 8'h44 == io_state_in_12 ? 8'h88 : _GEN_6211; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6213 = 8'h45 == io_state_in_12 ? 8'h8a : _GEN_6212; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6214 = 8'h46 == io_state_in_12 ? 8'h8c : _GEN_6213; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6215 = 8'h47 == io_state_in_12 ? 8'h8e : _GEN_6214; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6216 = 8'h48 == io_state_in_12 ? 8'h90 : _GEN_6215; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6217 = 8'h49 == io_state_in_12 ? 8'h92 : _GEN_6216; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6218 = 8'h4a == io_state_in_12 ? 8'h94 : _GEN_6217; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6219 = 8'h4b == io_state_in_12 ? 8'h96 : _GEN_6218; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6220 = 8'h4c == io_state_in_12 ? 8'h98 : _GEN_6219; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6221 = 8'h4d == io_state_in_12 ? 8'h9a : _GEN_6220; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6222 = 8'h4e == io_state_in_12 ? 8'h9c : _GEN_6221; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6223 = 8'h4f == io_state_in_12 ? 8'h9e : _GEN_6222; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6224 = 8'h50 == io_state_in_12 ? 8'ha0 : _GEN_6223; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6225 = 8'h51 == io_state_in_12 ? 8'ha2 : _GEN_6224; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6226 = 8'h52 == io_state_in_12 ? 8'ha4 : _GEN_6225; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6227 = 8'h53 == io_state_in_12 ? 8'ha6 : _GEN_6226; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6228 = 8'h54 == io_state_in_12 ? 8'ha8 : _GEN_6227; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6229 = 8'h55 == io_state_in_12 ? 8'haa : _GEN_6228; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6230 = 8'h56 == io_state_in_12 ? 8'hac : _GEN_6229; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6231 = 8'h57 == io_state_in_12 ? 8'hae : _GEN_6230; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6232 = 8'h58 == io_state_in_12 ? 8'hb0 : _GEN_6231; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6233 = 8'h59 == io_state_in_12 ? 8'hb2 : _GEN_6232; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6234 = 8'h5a == io_state_in_12 ? 8'hb4 : _GEN_6233; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6235 = 8'h5b == io_state_in_12 ? 8'hb6 : _GEN_6234; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6236 = 8'h5c == io_state_in_12 ? 8'hb8 : _GEN_6235; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6237 = 8'h5d == io_state_in_12 ? 8'hba : _GEN_6236; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6238 = 8'h5e == io_state_in_12 ? 8'hbc : _GEN_6237; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6239 = 8'h5f == io_state_in_12 ? 8'hbe : _GEN_6238; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6240 = 8'h60 == io_state_in_12 ? 8'hc0 : _GEN_6239; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6241 = 8'h61 == io_state_in_12 ? 8'hc2 : _GEN_6240; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6242 = 8'h62 == io_state_in_12 ? 8'hc4 : _GEN_6241; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6243 = 8'h63 == io_state_in_12 ? 8'hc6 : _GEN_6242; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6244 = 8'h64 == io_state_in_12 ? 8'hc8 : _GEN_6243; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6245 = 8'h65 == io_state_in_12 ? 8'hca : _GEN_6244; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6246 = 8'h66 == io_state_in_12 ? 8'hcc : _GEN_6245; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6247 = 8'h67 == io_state_in_12 ? 8'hce : _GEN_6246; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6248 = 8'h68 == io_state_in_12 ? 8'hd0 : _GEN_6247; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6249 = 8'h69 == io_state_in_12 ? 8'hd2 : _GEN_6248; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6250 = 8'h6a == io_state_in_12 ? 8'hd4 : _GEN_6249; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6251 = 8'h6b == io_state_in_12 ? 8'hd6 : _GEN_6250; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6252 = 8'h6c == io_state_in_12 ? 8'hd8 : _GEN_6251; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6253 = 8'h6d == io_state_in_12 ? 8'hda : _GEN_6252; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6254 = 8'h6e == io_state_in_12 ? 8'hdc : _GEN_6253; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6255 = 8'h6f == io_state_in_12 ? 8'hde : _GEN_6254; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6256 = 8'h70 == io_state_in_12 ? 8'he0 : _GEN_6255; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6257 = 8'h71 == io_state_in_12 ? 8'he2 : _GEN_6256; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6258 = 8'h72 == io_state_in_12 ? 8'he4 : _GEN_6257; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6259 = 8'h73 == io_state_in_12 ? 8'he6 : _GEN_6258; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6260 = 8'h74 == io_state_in_12 ? 8'he8 : _GEN_6259; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6261 = 8'h75 == io_state_in_12 ? 8'hea : _GEN_6260; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6262 = 8'h76 == io_state_in_12 ? 8'hec : _GEN_6261; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6263 = 8'h77 == io_state_in_12 ? 8'hee : _GEN_6262; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6264 = 8'h78 == io_state_in_12 ? 8'hf0 : _GEN_6263; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6265 = 8'h79 == io_state_in_12 ? 8'hf2 : _GEN_6264; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6266 = 8'h7a == io_state_in_12 ? 8'hf4 : _GEN_6265; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6267 = 8'h7b == io_state_in_12 ? 8'hf6 : _GEN_6266; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6268 = 8'h7c == io_state_in_12 ? 8'hf8 : _GEN_6267; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6269 = 8'h7d == io_state_in_12 ? 8'hfa : _GEN_6268; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6270 = 8'h7e == io_state_in_12 ? 8'hfc : _GEN_6269; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6271 = 8'h7f == io_state_in_12 ? 8'hfe : _GEN_6270; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6272 = 8'h80 == io_state_in_12 ? 8'h1b : _GEN_6271; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6273 = 8'h81 == io_state_in_12 ? 8'h19 : _GEN_6272; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6274 = 8'h82 == io_state_in_12 ? 8'h1f : _GEN_6273; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6275 = 8'h83 == io_state_in_12 ? 8'h1d : _GEN_6274; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6276 = 8'h84 == io_state_in_12 ? 8'h13 : _GEN_6275; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6277 = 8'h85 == io_state_in_12 ? 8'h11 : _GEN_6276; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6278 = 8'h86 == io_state_in_12 ? 8'h17 : _GEN_6277; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6279 = 8'h87 == io_state_in_12 ? 8'h15 : _GEN_6278; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6280 = 8'h88 == io_state_in_12 ? 8'hb : _GEN_6279; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6281 = 8'h89 == io_state_in_12 ? 8'h9 : _GEN_6280; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6282 = 8'h8a == io_state_in_12 ? 8'hf : _GEN_6281; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6283 = 8'h8b == io_state_in_12 ? 8'hd : _GEN_6282; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6284 = 8'h8c == io_state_in_12 ? 8'h3 : _GEN_6283; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6285 = 8'h8d == io_state_in_12 ? 8'h1 : _GEN_6284; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6286 = 8'h8e == io_state_in_12 ? 8'h7 : _GEN_6285; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6287 = 8'h8f == io_state_in_12 ? 8'h5 : _GEN_6286; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6288 = 8'h90 == io_state_in_12 ? 8'h3b : _GEN_6287; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6289 = 8'h91 == io_state_in_12 ? 8'h39 : _GEN_6288; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6290 = 8'h92 == io_state_in_12 ? 8'h3f : _GEN_6289; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6291 = 8'h93 == io_state_in_12 ? 8'h3d : _GEN_6290; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6292 = 8'h94 == io_state_in_12 ? 8'h33 : _GEN_6291; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6293 = 8'h95 == io_state_in_12 ? 8'h31 : _GEN_6292; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6294 = 8'h96 == io_state_in_12 ? 8'h37 : _GEN_6293; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6295 = 8'h97 == io_state_in_12 ? 8'h35 : _GEN_6294; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6296 = 8'h98 == io_state_in_12 ? 8'h2b : _GEN_6295; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6297 = 8'h99 == io_state_in_12 ? 8'h29 : _GEN_6296; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6298 = 8'h9a == io_state_in_12 ? 8'h2f : _GEN_6297; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6299 = 8'h9b == io_state_in_12 ? 8'h2d : _GEN_6298; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6300 = 8'h9c == io_state_in_12 ? 8'h23 : _GEN_6299; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6301 = 8'h9d == io_state_in_12 ? 8'h21 : _GEN_6300; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6302 = 8'h9e == io_state_in_12 ? 8'h27 : _GEN_6301; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6303 = 8'h9f == io_state_in_12 ? 8'h25 : _GEN_6302; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6304 = 8'ha0 == io_state_in_12 ? 8'h5b : _GEN_6303; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6305 = 8'ha1 == io_state_in_12 ? 8'h59 : _GEN_6304; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6306 = 8'ha2 == io_state_in_12 ? 8'h5f : _GEN_6305; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6307 = 8'ha3 == io_state_in_12 ? 8'h5d : _GEN_6306; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6308 = 8'ha4 == io_state_in_12 ? 8'h53 : _GEN_6307; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6309 = 8'ha5 == io_state_in_12 ? 8'h51 : _GEN_6308; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6310 = 8'ha6 == io_state_in_12 ? 8'h57 : _GEN_6309; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6311 = 8'ha7 == io_state_in_12 ? 8'h55 : _GEN_6310; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6312 = 8'ha8 == io_state_in_12 ? 8'h4b : _GEN_6311; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6313 = 8'ha9 == io_state_in_12 ? 8'h49 : _GEN_6312; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6314 = 8'haa == io_state_in_12 ? 8'h4f : _GEN_6313; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6315 = 8'hab == io_state_in_12 ? 8'h4d : _GEN_6314; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6316 = 8'hac == io_state_in_12 ? 8'h43 : _GEN_6315; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6317 = 8'had == io_state_in_12 ? 8'h41 : _GEN_6316; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6318 = 8'hae == io_state_in_12 ? 8'h47 : _GEN_6317; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6319 = 8'haf == io_state_in_12 ? 8'h45 : _GEN_6318; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6320 = 8'hb0 == io_state_in_12 ? 8'h7b : _GEN_6319; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6321 = 8'hb1 == io_state_in_12 ? 8'h79 : _GEN_6320; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6322 = 8'hb2 == io_state_in_12 ? 8'h7f : _GEN_6321; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6323 = 8'hb3 == io_state_in_12 ? 8'h7d : _GEN_6322; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6324 = 8'hb4 == io_state_in_12 ? 8'h73 : _GEN_6323; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6325 = 8'hb5 == io_state_in_12 ? 8'h71 : _GEN_6324; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6326 = 8'hb6 == io_state_in_12 ? 8'h77 : _GEN_6325; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6327 = 8'hb7 == io_state_in_12 ? 8'h75 : _GEN_6326; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6328 = 8'hb8 == io_state_in_12 ? 8'h6b : _GEN_6327; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6329 = 8'hb9 == io_state_in_12 ? 8'h69 : _GEN_6328; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6330 = 8'hba == io_state_in_12 ? 8'h6f : _GEN_6329; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6331 = 8'hbb == io_state_in_12 ? 8'h6d : _GEN_6330; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6332 = 8'hbc == io_state_in_12 ? 8'h63 : _GEN_6331; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6333 = 8'hbd == io_state_in_12 ? 8'h61 : _GEN_6332; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6334 = 8'hbe == io_state_in_12 ? 8'h67 : _GEN_6333; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6335 = 8'hbf == io_state_in_12 ? 8'h65 : _GEN_6334; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6336 = 8'hc0 == io_state_in_12 ? 8'h9b : _GEN_6335; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6337 = 8'hc1 == io_state_in_12 ? 8'h99 : _GEN_6336; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6338 = 8'hc2 == io_state_in_12 ? 8'h9f : _GEN_6337; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6339 = 8'hc3 == io_state_in_12 ? 8'h9d : _GEN_6338; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6340 = 8'hc4 == io_state_in_12 ? 8'h93 : _GEN_6339; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6341 = 8'hc5 == io_state_in_12 ? 8'h91 : _GEN_6340; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6342 = 8'hc6 == io_state_in_12 ? 8'h97 : _GEN_6341; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6343 = 8'hc7 == io_state_in_12 ? 8'h95 : _GEN_6342; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6344 = 8'hc8 == io_state_in_12 ? 8'h8b : _GEN_6343; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6345 = 8'hc9 == io_state_in_12 ? 8'h89 : _GEN_6344; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6346 = 8'hca == io_state_in_12 ? 8'h8f : _GEN_6345; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6347 = 8'hcb == io_state_in_12 ? 8'h8d : _GEN_6346; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6348 = 8'hcc == io_state_in_12 ? 8'h83 : _GEN_6347; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6349 = 8'hcd == io_state_in_12 ? 8'h81 : _GEN_6348; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6350 = 8'hce == io_state_in_12 ? 8'h87 : _GEN_6349; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6351 = 8'hcf == io_state_in_12 ? 8'h85 : _GEN_6350; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6352 = 8'hd0 == io_state_in_12 ? 8'hbb : _GEN_6351; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6353 = 8'hd1 == io_state_in_12 ? 8'hb9 : _GEN_6352; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6354 = 8'hd2 == io_state_in_12 ? 8'hbf : _GEN_6353; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6355 = 8'hd3 == io_state_in_12 ? 8'hbd : _GEN_6354; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6356 = 8'hd4 == io_state_in_12 ? 8'hb3 : _GEN_6355; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6357 = 8'hd5 == io_state_in_12 ? 8'hb1 : _GEN_6356; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6358 = 8'hd6 == io_state_in_12 ? 8'hb7 : _GEN_6357; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6359 = 8'hd7 == io_state_in_12 ? 8'hb5 : _GEN_6358; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6360 = 8'hd8 == io_state_in_12 ? 8'hab : _GEN_6359; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6361 = 8'hd9 == io_state_in_12 ? 8'ha9 : _GEN_6360; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6362 = 8'hda == io_state_in_12 ? 8'haf : _GEN_6361; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6363 = 8'hdb == io_state_in_12 ? 8'had : _GEN_6362; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6364 = 8'hdc == io_state_in_12 ? 8'ha3 : _GEN_6363; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6365 = 8'hdd == io_state_in_12 ? 8'ha1 : _GEN_6364; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6366 = 8'hde == io_state_in_12 ? 8'ha7 : _GEN_6365; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6367 = 8'hdf == io_state_in_12 ? 8'ha5 : _GEN_6366; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6368 = 8'he0 == io_state_in_12 ? 8'hdb : _GEN_6367; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6369 = 8'he1 == io_state_in_12 ? 8'hd9 : _GEN_6368; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6370 = 8'he2 == io_state_in_12 ? 8'hdf : _GEN_6369; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6371 = 8'he3 == io_state_in_12 ? 8'hdd : _GEN_6370; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6372 = 8'he4 == io_state_in_12 ? 8'hd3 : _GEN_6371; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6373 = 8'he5 == io_state_in_12 ? 8'hd1 : _GEN_6372; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6374 = 8'he6 == io_state_in_12 ? 8'hd7 : _GEN_6373; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6375 = 8'he7 == io_state_in_12 ? 8'hd5 : _GEN_6374; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6376 = 8'he8 == io_state_in_12 ? 8'hcb : _GEN_6375; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6377 = 8'he9 == io_state_in_12 ? 8'hc9 : _GEN_6376; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6378 = 8'hea == io_state_in_12 ? 8'hcf : _GEN_6377; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6379 = 8'heb == io_state_in_12 ? 8'hcd : _GEN_6378; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6380 = 8'hec == io_state_in_12 ? 8'hc3 : _GEN_6379; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6381 = 8'hed == io_state_in_12 ? 8'hc1 : _GEN_6380; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6382 = 8'hee == io_state_in_12 ? 8'hc7 : _GEN_6381; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6383 = 8'hef == io_state_in_12 ? 8'hc5 : _GEN_6382; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6384 = 8'hf0 == io_state_in_12 ? 8'hfb : _GEN_6383; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6385 = 8'hf1 == io_state_in_12 ? 8'hf9 : _GEN_6384; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6386 = 8'hf2 == io_state_in_12 ? 8'hff : _GEN_6385; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6387 = 8'hf3 == io_state_in_12 ? 8'hfd : _GEN_6386; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6388 = 8'hf4 == io_state_in_12 ? 8'hf3 : _GEN_6387; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6389 = 8'hf5 == io_state_in_12 ? 8'hf1 : _GEN_6388; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6390 = 8'hf6 == io_state_in_12 ? 8'hf7 : _GEN_6389; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6391 = 8'hf7 == io_state_in_12 ? 8'hf5 : _GEN_6390; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6392 = 8'hf8 == io_state_in_12 ? 8'heb : _GEN_6391; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6393 = 8'hf9 == io_state_in_12 ? 8'he9 : _GEN_6392; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6394 = 8'hfa == io_state_in_12 ? 8'hef : _GEN_6393; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6395 = 8'hfb == io_state_in_12 ? 8'hed : _GEN_6394; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6396 = 8'hfc == io_state_in_12 ? 8'he3 : _GEN_6395; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6397 = 8'hfd == io_state_in_12 ? 8'he1 : _GEN_6396; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6398 = 8'hfe == io_state_in_12 ? 8'he7 : _GEN_6397; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6399 = 8'hff == io_state_in_12 ? 8'he5 : _GEN_6398; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6401 = 8'h1 == io_state_in_13 ? 8'h3 : 8'h0; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6402 = 8'h2 == io_state_in_13 ? 8'h6 : _GEN_6401; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6403 = 8'h3 == io_state_in_13 ? 8'h5 : _GEN_6402; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6404 = 8'h4 == io_state_in_13 ? 8'hc : _GEN_6403; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6405 = 8'h5 == io_state_in_13 ? 8'hf : _GEN_6404; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6406 = 8'h6 == io_state_in_13 ? 8'ha : _GEN_6405; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6407 = 8'h7 == io_state_in_13 ? 8'h9 : _GEN_6406; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6408 = 8'h8 == io_state_in_13 ? 8'h18 : _GEN_6407; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6409 = 8'h9 == io_state_in_13 ? 8'h1b : _GEN_6408; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6410 = 8'ha == io_state_in_13 ? 8'h1e : _GEN_6409; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6411 = 8'hb == io_state_in_13 ? 8'h1d : _GEN_6410; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6412 = 8'hc == io_state_in_13 ? 8'h14 : _GEN_6411; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6413 = 8'hd == io_state_in_13 ? 8'h17 : _GEN_6412; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6414 = 8'he == io_state_in_13 ? 8'h12 : _GEN_6413; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6415 = 8'hf == io_state_in_13 ? 8'h11 : _GEN_6414; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6416 = 8'h10 == io_state_in_13 ? 8'h30 : _GEN_6415; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6417 = 8'h11 == io_state_in_13 ? 8'h33 : _GEN_6416; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6418 = 8'h12 == io_state_in_13 ? 8'h36 : _GEN_6417; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6419 = 8'h13 == io_state_in_13 ? 8'h35 : _GEN_6418; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6420 = 8'h14 == io_state_in_13 ? 8'h3c : _GEN_6419; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6421 = 8'h15 == io_state_in_13 ? 8'h3f : _GEN_6420; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6422 = 8'h16 == io_state_in_13 ? 8'h3a : _GEN_6421; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6423 = 8'h17 == io_state_in_13 ? 8'h39 : _GEN_6422; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6424 = 8'h18 == io_state_in_13 ? 8'h28 : _GEN_6423; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6425 = 8'h19 == io_state_in_13 ? 8'h2b : _GEN_6424; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6426 = 8'h1a == io_state_in_13 ? 8'h2e : _GEN_6425; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6427 = 8'h1b == io_state_in_13 ? 8'h2d : _GEN_6426; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6428 = 8'h1c == io_state_in_13 ? 8'h24 : _GEN_6427; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6429 = 8'h1d == io_state_in_13 ? 8'h27 : _GEN_6428; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6430 = 8'h1e == io_state_in_13 ? 8'h22 : _GEN_6429; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6431 = 8'h1f == io_state_in_13 ? 8'h21 : _GEN_6430; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6432 = 8'h20 == io_state_in_13 ? 8'h60 : _GEN_6431; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6433 = 8'h21 == io_state_in_13 ? 8'h63 : _GEN_6432; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6434 = 8'h22 == io_state_in_13 ? 8'h66 : _GEN_6433; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6435 = 8'h23 == io_state_in_13 ? 8'h65 : _GEN_6434; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6436 = 8'h24 == io_state_in_13 ? 8'h6c : _GEN_6435; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6437 = 8'h25 == io_state_in_13 ? 8'h6f : _GEN_6436; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6438 = 8'h26 == io_state_in_13 ? 8'h6a : _GEN_6437; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6439 = 8'h27 == io_state_in_13 ? 8'h69 : _GEN_6438; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6440 = 8'h28 == io_state_in_13 ? 8'h78 : _GEN_6439; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6441 = 8'h29 == io_state_in_13 ? 8'h7b : _GEN_6440; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6442 = 8'h2a == io_state_in_13 ? 8'h7e : _GEN_6441; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6443 = 8'h2b == io_state_in_13 ? 8'h7d : _GEN_6442; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6444 = 8'h2c == io_state_in_13 ? 8'h74 : _GEN_6443; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6445 = 8'h2d == io_state_in_13 ? 8'h77 : _GEN_6444; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6446 = 8'h2e == io_state_in_13 ? 8'h72 : _GEN_6445; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6447 = 8'h2f == io_state_in_13 ? 8'h71 : _GEN_6446; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6448 = 8'h30 == io_state_in_13 ? 8'h50 : _GEN_6447; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6449 = 8'h31 == io_state_in_13 ? 8'h53 : _GEN_6448; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6450 = 8'h32 == io_state_in_13 ? 8'h56 : _GEN_6449; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6451 = 8'h33 == io_state_in_13 ? 8'h55 : _GEN_6450; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6452 = 8'h34 == io_state_in_13 ? 8'h5c : _GEN_6451; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6453 = 8'h35 == io_state_in_13 ? 8'h5f : _GEN_6452; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6454 = 8'h36 == io_state_in_13 ? 8'h5a : _GEN_6453; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6455 = 8'h37 == io_state_in_13 ? 8'h59 : _GEN_6454; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6456 = 8'h38 == io_state_in_13 ? 8'h48 : _GEN_6455; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6457 = 8'h39 == io_state_in_13 ? 8'h4b : _GEN_6456; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6458 = 8'h3a == io_state_in_13 ? 8'h4e : _GEN_6457; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6459 = 8'h3b == io_state_in_13 ? 8'h4d : _GEN_6458; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6460 = 8'h3c == io_state_in_13 ? 8'h44 : _GEN_6459; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6461 = 8'h3d == io_state_in_13 ? 8'h47 : _GEN_6460; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6462 = 8'h3e == io_state_in_13 ? 8'h42 : _GEN_6461; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6463 = 8'h3f == io_state_in_13 ? 8'h41 : _GEN_6462; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6464 = 8'h40 == io_state_in_13 ? 8'hc0 : _GEN_6463; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6465 = 8'h41 == io_state_in_13 ? 8'hc3 : _GEN_6464; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6466 = 8'h42 == io_state_in_13 ? 8'hc6 : _GEN_6465; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6467 = 8'h43 == io_state_in_13 ? 8'hc5 : _GEN_6466; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6468 = 8'h44 == io_state_in_13 ? 8'hcc : _GEN_6467; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6469 = 8'h45 == io_state_in_13 ? 8'hcf : _GEN_6468; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6470 = 8'h46 == io_state_in_13 ? 8'hca : _GEN_6469; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6471 = 8'h47 == io_state_in_13 ? 8'hc9 : _GEN_6470; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6472 = 8'h48 == io_state_in_13 ? 8'hd8 : _GEN_6471; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6473 = 8'h49 == io_state_in_13 ? 8'hdb : _GEN_6472; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6474 = 8'h4a == io_state_in_13 ? 8'hde : _GEN_6473; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6475 = 8'h4b == io_state_in_13 ? 8'hdd : _GEN_6474; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6476 = 8'h4c == io_state_in_13 ? 8'hd4 : _GEN_6475; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6477 = 8'h4d == io_state_in_13 ? 8'hd7 : _GEN_6476; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6478 = 8'h4e == io_state_in_13 ? 8'hd2 : _GEN_6477; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6479 = 8'h4f == io_state_in_13 ? 8'hd1 : _GEN_6478; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6480 = 8'h50 == io_state_in_13 ? 8'hf0 : _GEN_6479; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6481 = 8'h51 == io_state_in_13 ? 8'hf3 : _GEN_6480; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6482 = 8'h52 == io_state_in_13 ? 8'hf6 : _GEN_6481; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6483 = 8'h53 == io_state_in_13 ? 8'hf5 : _GEN_6482; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6484 = 8'h54 == io_state_in_13 ? 8'hfc : _GEN_6483; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6485 = 8'h55 == io_state_in_13 ? 8'hff : _GEN_6484; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6486 = 8'h56 == io_state_in_13 ? 8'hfa : _GEN_6485; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6487 = 8'h57 == io_state_in_13 ? 8'hf9 : _GEN_6486; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6488 = 8'h58 == io_state_in_13 ? 8'he8 : _GEN_6487; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6489 = 8'h59 == io_state_in_13 ? 8'heb : _GEN_6488; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6490 = 8'h5a == io_state_in_13 ? 8'hee : _GEN_6489; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6491 = 8'h5b == io_state_in_13 ? 8'hed : _GEN_6490; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6492 = 8'h5c == io_state_in_13 ? 8'he4 : _GEN_6491; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6493 = 8'h5d == io_state_in_13 ? 8'he7 : _GEN_6492; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6494 = 8'h5e == io_state_in_13 ? 8'he2 : _GEN_6493; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6495 = 8'h5f == io_state_in_13 ? 8'he1 : _GEN_6494; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6496 = 8'h60 == io_state_in_13 ? 8'ha0 : _GEN_6495; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6497 = 8'h61 == io_state_in_13 ? 8'ha3 : _GEN_6496; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6498 = 8'h62 == io_state_in_13 ? 8'ha6 : _GEN_6497; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6499 = 8'h63 == io_state_in_13 ? 8'ha5 : _GEN_6498; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6500 = 8'h64 == io_state_in_13 ? 8'hac : _GEN_6499; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6501 = 8'h65 == io_state_in_13 ? 8'haf : _GEN_6500; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6502 = 8'h66 == io_state_in_13 ? 8'haa : _GEN_6501; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6503 = 8'h67 == io_state_in_13 ? 8'ha9 : _GEN_6502; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6504 = 8'h68 == io_state_in_13 ? 8'hb8 : _GEN_6503; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6505 = 8'h69 == io_state_in_13 ? 8'hbb : _GEN_6504; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6506 = 8'h6a == io_state_in_13 ? 8'hbe : _GEN_6505; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6507 = 8'h6b == io_state_in_13 ? 8'hbd : _GEN_6506; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6508 = 8'h6c == io_state_in_13 ? 8'hb4 : _GEN_6507; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6509 = 8'h6d == io_state_in_13 ? 8'hb7 : _GEN_6508; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6510 = 8'h6e == io_state_in_13 ? 8'hb2 : _GEN_6509; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6511 = 8'h6f == io_state_in_13 ? 8'hb1 : _GEN_6510; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6512 = 8'h70 == io_state_in_13 ? 8'h90 : _GEN_6511; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6513 = 8'h71 == io_state_in_13 ? 8'h93 : _GEN_6512; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6514 = 8'h72 == io_state_in_13 ? 8'h96 : _GEN_6513; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6515 = 8'h73 == io_state_in_13 ? 8'h95 : _GEN_6514; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6516 = 8'h74 == io_state_in_13 ? 8'h9c : _GEN_6515; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6517 = 8'h75 == io_state_in_13 ? 8'h9f : _GEN_6516; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6518 = 8'h76 == io_state_in_13 ? 8'h9a : _GEN_6517; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6519 = 8'h77 == io_state_in_13 ? 8'h99 : _GEN_6518; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6520 = 8'h78 == io_state_in_13 ? 8'h88 : _GEN_6519; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6521 = 8'h79 == io_state_in_13 ? 8'h8b : _GEN_6520; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6522 = 8'h7a == io_state_in_13 ? 8'h8e : _GEN_6521; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6523 = 8'h7b == io_state_in_13 ? 8'h8d : _GEN_6522; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6524 = 8'h7c == io_state_in_13 ? 8'h84 : _GEN_6523; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6525 = 8'h7d == io_state_in_13 ? 8'h87 : _GEN_6524; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6526 = 8'h7e == io_state_in_13 ? 8'h82 : _GEN_6525; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6527 = 8'h7f == io_state_in_13 ? 8'h81 : _GEN_6526; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6528 = 8'h80 == io_state_in_13 ? 8'h9b : _GEN_6527; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6529 = 8'h81 == io_state_in_13 ? 8'h98 : _GEN_6528; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6530 = 8'h82 == io_state_in_13 ? 8'h9d : _GEN_6529; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6531 = 8'h83 == io_state_in_13 ? 8'h9e : _GEN_6530; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6532 = 8'h84 == io_state_in_13 ? 8'h97 : _GEN_6531; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6533 = 8'h85 == io_state_in_13 ? 8'h94 : _GEN_6532; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6534 = 8'h86 == io_state_in_13 ? 8'h91 : _GEN_6533; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6535 = 8'h87 == io_state_in_13 ? 8'h92 : _GEN_6534; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6536 = 8'h88 == io_state_in_13 ? 8'h83 : _GEN_6535; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6537 = 8'h89 == io_state_in_13 ? 8'h80 : _GEN_6536; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6538 = 8'h8a == io_state_in_13 ? 8'h85 : _GEN_6537; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6539 = 8'h8b == io_state_in_13 ? 8'h86 : _GEN_6538; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6540 = 8'h8c == io_state_in_13 ? 8'h8f : _GEN_6539; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6541 = 8'h8d == io_state_in_13 ? 8'h8c : _GEN_6540; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6542 = 8'h8e == io_state_in_13 ? 8'h89 : _GEN_6541; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6543 = 8'h8f == io_state_in_13 ? 8'h8a : _GEN_6542; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6544 = 8'h90 == io_state_in_13 ? 8'hab : _GEN_6543; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6545 = 8'h91 == io_state_in_13 ? 8'ha8 : _GEN_6544; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6546 = 8'h92 == io_state_in_13 ? 8'had : _GEN_6545; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6547 = 8'h93 == io_state_in_13 ? 8'hae : _GEN_6546; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6548 = 8'h94 == io_state_in_13 ? 8'ha7 : _GEN_6547; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6549 = 8'h95 == io_state_in_13 ? 8'ha4 : _GEN_6548; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6550 = 8'h96 == io_state_in_13 ? 8'ha1 : _GEN_6549; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6551 = 8'h97 == io_state_in_13 ? 8'ha2 : _GEN_6550; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6552 = 8'h98 == io_state_in_13 ? 8'hb3 : _GEN_6551; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6553 = 8'h99 == io_state_in_13 ? 8'hb0 : _GEN_6552; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6554 = 8'h9a == io_state_in_13 ? 8'hb5 : _GEN_6553; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6555 = 8'h9b == io_state_in_13 ? 8'hb6 : _GEN_6554; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6556 = 8'h9c == io_state_in_13 ? 8'hbf : _GEN_6555; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6557 = 8'h9d == io_state_in_13 ? 8'hbc : _GEN_6556; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6558 = 8'h9e == io_state_in_13 ? 8'hb9 : _GEN_6557; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6559 = 8'h9f == io_state_in_13 ? 8'hba : _GEN_6558; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6560 = 8'ha0 == io_state_in_13 ? 8'hfb : _GEN_6559; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6561 = 8'ha1 == io_state_in_13 ? 8'hf8 : _GEN_6560; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6562 = 8'ha2 == io_state_in_13 ? 8'hfd : _GEN_6561; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6563 = 8'ha3 == io_state_in_13 ? 8'hfe : _GEN_6562; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6564 = 8'ha4 == io_state_in_13 ? 8'hf7 : _GEN_6563; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6565 = 8'ha5 == io_state_in_13 ? 8'hf4 : _GEN_6564; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6566 = 8'ha6 == io_state_in_13 ? 8'hf1 : _GEN_6565; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6567 = 8'ha7 == io_state_in_13 ? 8'hf2 : _GEN_6566; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6568 = 8'ha8 == io_state_in_13 ? 8'he3 : _GEN_6567; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6569 = 8'ha9 == io_state_in_13 ? 8'he0 : _GEN_6568; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6570 = 8'haa == io_state_in_13 ? 8'he5 : _GEN_6569; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6571 = 8'hab == io_state_in_13 ? 8'he6 : _GEN_6570; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6572 = 8'hac == io_state_in_13 ? 8'hef : _GEN_6571; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6573 = 8'had == io_state_in_13 ? 8'hec : _GEN_6572; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6574 = 8'hae == io_state_in_13 ? 8'he9 : _GEN_6573; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6575 = 8'haf == io_state_in_13 ? 8'hea : _GEN_6574; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6576 = 8'hb0 == io_state_in_13 ? 8'hcb : _GEN_6575; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6577 = 8'hb1 == io_state_in_13 ? 8'hc8 : _GEN_6576; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6578 = 8'hb2 == io_state_in_13 ? 8'hcd : _GEN_6577; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6579 = 8'hb3 == io_state_in_13 ? 8'hce : _GEN_6578; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6580 = 8'hb4 == io_state_in_13 ? 8'hc7 : _GEN_6579; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6581 = 8'hb5 == io_state_in_13 ? 8'hc4 : _GEN_6580; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6582 = 8'hb6 == io_state_in_13 ? 8'hc1 : _GEN_6581; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6583 = 8'hb7 == io_state_in_13 ? 8'hc2 : _GEN_6582; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6584 = 8'hb8 == io_state_in_13 ? 8'hd3 : _GEN_6583; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6585 = 8'hb9 == io_state_in_13 ? 8'hd0 : _GEN_6584; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6586 = 8'hba == io_state_in_13 ? 8'hd5 : _GEN_6585; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6587 = 8'hbb == io_state_in_13 ? 8'hd6 : _GEN_6586; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6588 = 8'hbc == io_state_in_13 ? 8'hdf : _GEN_6587; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6589 = 8'hbd == io_state_in_13 ? 8'hdc : _GEN_6588; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6590 = 8'hbe == io_state_in_13 ? 8'hd9 : _GEN_6589; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6591 = 8'hbf == io_state_in_13 ? 8'hda : _GEN_6590; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6592 = 8'hc0 == io_state_in_13 ? 8'h5b : _GEN_6591; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6593 = 8'hc1 == io_state_in_13 ? 8'h58 : _GEN_6592; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6594 = 8'hc2 == io_state_in_13 ? 8'h5d : _GEN_6593; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6595 = 8'hc3 == io_state_in_13 ? 8'h5e : _GEN_6594; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6596 = 8'hc4 == io_state_in_13 ? 8'h57 : _GEN_6595; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6597 = 8'hc5 == io_state_in_13 ? 8'h54 : _GEN_6596; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6598 = 8'hc6 == io_state_in_13 ? 8'h51 : _GEN_6597; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6599 = 8'hc7 == io_state_in_13 ? 8'h52 : _GEN_6598; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6600 = 8'hc8 == io_state_in_13 ? 8'h43 : _GEN_6599; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6601 = 8'hc9 == io_state_in_13 ? 8'h40 : _GEN_6600; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6602 = 8'hca == io_state_in_13 ? 8'h45 : _GEN_6601; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6603 = 8'hcb == io_state_in_13 ? 8'h46 : _GEN_6602; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6604 = 8'hcc == io_state_in_13 ? 8'h4f : _GEN_6603; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6605 = 8'hcd == io_state_in_13 ? 8'h4c : _GEN_6604; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6606 = 8'hce == io_state_in_13 ? 8'h49 : _GEN_6605; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6607 = 8'hcf == io_state_in_13 ? 8'h4a : _GEN_6606; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6608 = 8'hd0 == io_state_in_13 ? 8'h6b : _GEN_6607; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6609 = 8'hd1 == io_state_in_13 ? 8'h68 : _GEN_6608; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6610 = 8'hd2 == io_state_in_13 ? 8'h6d : _GEN_6609; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6611 = 8'hd3 == io_state_in_13 ? 8'h6e : _GEN_6610; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6612 = 8'hd4 == io_state_in_13 ? 8'h67 : _GEN_6611; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6613 = 8'hd5 == io_state_in_13 ? 8'h64 : _GEN_6612; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6614 = 8'hd6 == io_state_in_13 ? 8'h61 : _GEN_6613; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6615 = 8'hd7 == io_state_in_13 ? 8'h62 : _GEN_6614; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6616 = 8'hd8 == io_state_in_13 ? 8'h73 : _GEN_6615; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6617 = 8'hd9 == io_state_in_13 ? 8'h70 : _GEN_6616; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6618 = 8'hda == io_state_in_13 ? 8'h75 : _GEN_6617; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6619 = 8'hdb == io_state_in_13 ? 8'h76 : _GEN_6618; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6620 = 8'hdc == io_state_in_13 ? 8'h7f : _GEN_6619; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6621 = 8'hdd == io_state_in_13 ? 8'h7c : _GEN_6620; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6622 = 8'hde == io_state_in_13 ? 8'h79 : _GEN_6621; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6623 = 8'hdf == io_state_in_13 ? 8'h7a : _GEN_6622; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6624 = 8'he0 == io_state_in_13 ? 8'h3b : _GEN_6623; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6625 = 8'he1 == io_state_in_13 ? 8'h38 : _GEN_6624; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6626 = 8'he2 == io_state_in_13 ? 8'h3d : _GEN_6625; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6627 = 8'he3 == io_state_in_13 ? 8'h3e : _GEN_6626; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6628 = 8'he4 == io_state_in_13 ? 8'h37 : _GEN_6627; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6629 = 8'he5 == io_state_in_13 ? 8'h34 : _GEN_6628; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6630 = 8'he6 == io_state_in_13 ? 8'h31 : _GEN_6629; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6631 = 8'he7 == io_state_in_13 ? 8'h32 : _GEN_6630; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6632 = 8'he8 == io_state_in_13 ? 8'h23 : _GEN_6631; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6633 = 8'he9 == io_state_in_13 ? 8'h20 : _GEN_6632; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6634 = 8'hea == io_state_in_13 ? 8'h25 : _GEN_6633; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6635 = 8'heb == io_state_in_13 ? 8'h26 : _GEN_6634; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6636 = 8'hec == io_state_in_13 ? 8'h2f : _GEN_6635; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6637 = 8'hed == io_state_in_13 ? 8'h2c : _GEN_6636; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6638 = 8'hee == io_state_in_13 ? 8'h29 : _GEN_6637; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6639 = 8'hef == io_state_in_13 ? 8'h2a : _GEN_6638; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6640 = 8'hf0 == io_state_in_13 ? 8'hb : _GEN_6639; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6641 = 8'hf1 == io_state_in_13 ? 8'h8 : _GEN_6640; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6642 = 8'hf2 == io_state_in_13 ? 8'hd : _GEN_6641; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6643 = 8'hf3 == io_state_in_13 ? 8'he : _GEN_6642; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6644 = 8'hf4 == io_state_in_13 ? 8'h7 : _GEN_6643; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6645 = 8'hf5 == io_state_in_13 ? 8'h4 : _GEN_6644; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6646 = 8'hf6 == io_state_in_13 ? 8'h1 : _GEN_6645; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6647 = 8'hf7 == io_state_in_13 ? 8'h2 : _GEN_6646; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6648 = 8'hf8 == io_state_in_13 ? 8'h13 : _GEN_6647; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6649 = 8'hf9 == io_state_in_13 ? 8'h10 : _GEN_6648; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6650 = 8'hfa == io_state_in_13 ? 8'h15 : _GEN_6649; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6651 = 8'hfb == io_state_in_13 ? 8'h16 : _GEN_6650; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6652 = 8'hfc == io_state_in_13 ? 8'h1f : _GEN_6651; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6653 = 8'hfd == io_state_in_13 ? 8'h1c : _GEN_6652; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6654 = 8'hfe == io_state_in_13 ? 8'h19 : _GEN_6653; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _GEN_6655 = 8'hff == io_state_in_13 ? 8'h1a : _GEN_6654; // @[MixColumns.scala 140:{43,43}]
  wire [7:0] _tmp_state_12_T = _GEN_6399 ^ _GEN_6655; // @[MixColumns.scala 140:43]
  wire [7:0] _tmp_state_12_T_1 = _tmp_state_12_T ^ io_state_in_14; // @[MixColumns.scala 140:68]
  wire [7:0] _GEN_6657 = 8'h1 == io_state_in_13 ? 8'h2 : 8'h0; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6658 = 8'h2 == io_state_in_13 ? 8'h4 : _GEN_6657; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6659 = 8'h3 == io_state_in_13 ? 8'h6 : _GEN_6658; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6660 = 8'h4 == io_state_in_13 ? 8'h8 : _GEN_6659; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6661 = 8'h5 == io_state_in_13 ? 8'ha : _GEN_6660; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6662 = 8'h6 == io_state_in_13 ? 8'hc : _GEN_6661; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6663 = 8'h7 == io_state_in_13 ? 8'he : _GEN_6662; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6664 = 8'h8 == io_state_in_13 ? 8'h10 : _GEN_6663; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6665 = 8'h9 == io_state_in_13 ? 8'h12 : _GEN_6664; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6666 = 8'ha == io_state_in_13 ? 8'h14 : _GEN_6665; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6667 = 8'hb == io_state_in_13 ? 8'h16 : _GEN_6666; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6668 = 8'hc == io_state_in_13 ? 8'h18 : _GEN_6667; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6669 = 8'hd == io_state_in_13 ? 8'h1a : _GEN_6668; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6670 = 8'he == io_state_in_13 ? 8'h1c : _GEN_6669; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6671 = 8'hf == io_state_in_13 ? 8'h1e : _GEN_6670; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6672 = 8'h10 == io_state_in_13 ? 8'h20 : _GEN_6671; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6673 = 8'h11 == io_state_in_13 ? 8'h22 : _GEN_6672; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6674 = 8'h12 == io_state_in_13 ? 8'h24 : _GEN_6673; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6675 = 8'h13 == io_state_in_13 ? 8'h26 : _GEN_6674; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6676 = 8'h14 == io_state_in_13 ? 8'h28 : _GEN_6675; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6677 = 8'h15 == io_state_in_13 ? 8'h2a : _GEN_6676; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6678 = 8'h16 == io_state_in_13 ? 8'h2c : _GEN_6677; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6679 = 8'h17 == io_state_in_13 ? 8'h2e : _GEN_6678; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6680 = 8'h18 == io_state_in_13 ? 8'h30 : _GEN_6679; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6681 = 8'h19 == io_state_in_13 ? 8'h32 : _GEN_6680; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6682 = 8'h1a == io_state_in_13 ? 8'h34 : _GEN_6681; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6683 = 8'h1b == io_state_in_13 ? 8'h36 : _GEN_6682; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6684 = 8'h1c == io_state_in_13 ? 8'h38 : _GEN_6683; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6685 = 8'h1d == io_state_in_13 ? 8'h3a : _GEN_6684; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6686 = 8'h1e == io_state_in_13 ? 8'h3c : _GEN_6685; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6687 = 8'h1f == io_state_in_13 ? 8'h3e : _GEN_6686; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6688 = 8'h20 == io_state_in_13 ? 8'h40 : _GEN_6687; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6689 = 8'h21 == io_state_in_13 ? 8'h42 : _GEN_6688; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6690 = 8'h22 == io_state_in_13 ? 8'h44 : _GEN_6689; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6691 = 8'h23 == io_state_in_13 ? 8'h46 : _GEN_6690; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6692 = 8'h24 == io_state_in_13 ? 8'h48 : _GEN_6691; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6693 = 8'h25 == io_state_in_13 ? 8'h4a : _GEN_6692; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6694 = 8'h26 == io_state_in_13 ? 8'h4c : _GEN_6693; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6695 = 8'h27 == io_state_in_13 ? 8'h4e : _GEN_6694; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6696 = 8'h28 == io_state_in_13 ? 8'h50 : _GEN_6695; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6697 = 8'h29 == io_state_in_13 ? 8'h52 : _GEN_6696; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6698 = 8'h2a == io_state_in_13 ? 8'h54 : _GEN_6697; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6699 = 8'h2b == io_state_in_13 ? 8'h56 : _GEN_6698; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6700 = 8'h2c == io_state_in_13 ? 8'h58 : _GEN_6699; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6701 = 8'h2d == io_state_in_13 ? 8'h5a : _GEN_6700; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6702 = 8'h2e == io_state_in_13 ? 8'h5c : _GEN_6701; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6703 = 8'h2f == io_state_in_13 ? 8'h5e : _GEN_6702; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6704 = 8'h30 == io_state_in_13 ? 8'h60 : _GEN_6703; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6705 = 8'h31 == io_state_in_13 ? 8'h62 : _GEN_6704; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6706 = 8'h32 == io_state_in_13 ? 8'h64 : _GEN_6705; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6707 = 8'h33 == io_state_in_13 ? 8'h66 : _GEN_6706; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6708 = 8'h34 == io_state_in_13 ? 8'h68 : _GEN_6707; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6709 = 8'h35 == io_state_in_13 ? 8'h6a : _GEN_6708; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6710 = 8'h36 == io_state_in_13 ? 8'h6c : _GEN_6709; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6711 = 8'h37 == io_state_in_13 ? 8'h6e : _GEN_6710; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6712 = 8'h38 == io_state_in_13 ? 8'h70 : _GEN_6711; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6713 = 8'h39 == io_state_in_13 ? 8'h72 : _GEN_6712; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6714 = 8'h3a == io_state_in_13 ? 8'h74 : _GEN_6713; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6715 = 8'h3b == io_state_in_13 ? 8'h76 : _GEN_6714; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6716 = 8'h3c == io_state_in_13 ? 8'h78 : _GEN_6715; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6717 = 8'h3d == io_state_in_13 ? 8'h7a : _GEN_6716; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6718 = 8'h3e == io_state_in_13 ? 8'h7c : _GEN_6717; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6719 = 8'h3f == io_state_in_13 ? 8'h7e : _GEN_6718; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6720 = 8'h40 == io_state_in_13 ? 8'h80 : _GEN_6719; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6721 = 8'h41 == io_state_in_13 ? 8'h82 : _GEN_6720; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6722 = 8'h42 == io_state_in_13 ? 8'h84 : _GEN_6721; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6723 = 8'h43 == io_state_in_13 ? 8'h86 : _GEN_6722; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6724 = 8'h44 == io_state_in_13 ? 8'h88 : _GEN_6723; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6725 = 8'h45 == io_state_in_13 ? 8'h8a : _GEN_6724; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6726 = 8'h46 == io_state_in_13 ? 8'h8c : _GEN_6725; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6727 = 8'h47 == io_state_in_13 ? 8'h8e : _GEN_6726; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6728 = 8'h48 == io_state_in_13 ? 8'h90 : _GEN_6727; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6729 = 8'h49 == io_state_in_13 ? 8'h92 : _GEN_6728; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6730 = 8'h4a == io_state_in_13 ? 8'h94 : _GEN_6729; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6731 = 8'h4b == io_state_in_13 ? 8'h96 : _GEN_6730; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6732 = 8'h4c == io_state_in_13 ? 8'h98 : _GEN_6731; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6733 = 8'h4d == io_state_in_13 ? 8'h9a : _GEN_6732; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6734 = 8'h4e == io_state_in_13 ? 8'h9c : _GEN_6733; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6735 = 8'h4f == io_state_in_13 ? 8'h9e : _GEN_6734; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6736 = 8'h50 == io_state_in_13 ? 8'ha0 : _GEN_6735; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6737 = 8'h51 == io_state_in_13 ? 8'ha2 : _GEN_6736; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6738 = 8'h52 == io_state_in_13 ? 8'ha4 : _GEN_6737; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6739 = 8'h53 == io_state_in_13 ? 8'ha6 : _GEN_6738; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6740 = 8'h54 == io_state_in_13 ? 8'ha8 : _GEN_6739; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6741 = 8'h55 == io_state_in_13 ? 8'haa : _GEN_6740; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6742 = 8'h56 == io_state_in_13 ? 8'hac : _GEN_6741; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6743 = 8'h57 == io_state_in_13 ? 8'hae : _GEN_6742; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6744 = 8'h58 == io_state_in_13 ? 8'hb0 : _GEN_6743; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6745 = 8'h59 == io_state_in_13 ? 8'hb2 : _GEN_6744; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6746 = 8'h5a == io_state_in_13 ? 8'hb4 : _GEN_6745; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6747 = 8'h5b == io_state_in_13 ? 8'hb6 : _GEN_6746; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6748 = 8'h5c == io_state_in_13 ? 8'hb8 : _GEN_6747; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6749 = 8'h5d == io_state_in_13 ? 8'hba : _GEN_6748; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6750 = 8'h5e == io_state_in_13 ? 8'hbc : _GEN_6749; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6751 = 8'h5f == io_state_in_13 ? 8'hbe : _GEN_6750; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6752 = 8'h60 == io_state_in_13 ? 8'hc0 : _GEN_6751; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6753 = 8'h61 == io_state_in_13 ? 8'hc2 : _GEN_6752; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6754 = 8'h62 == io_state_in_13 ? 8'hc4 : _GEN_6753; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6755 = 8'h63 == io_state_in_13 ? 8'hc6 : _GEN_6754; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6756 = 8'h64 == io_state_in_13 ? 8'hc8 : _GEN_6755; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6757 = 8'h65 == io_state_in_13 ? 8'hca : _GEN_6756; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6758 = 8'h66 == io_state_in_13 ? 8'hcc : _GEN_6757; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6759 = 8'h67 == io_state_in_13 ? 8'hce : _GEN_6758; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6760 = 8'h68 == io_state_in_13 ? 8'hd0 : _GEN_6759; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6761 = 8'h69 == io_state_in_13 ? 8'hd2 : _GEN_6760; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6762 = 8'h6a == io_state_in_13 ? 8'hd4 : _GEN_6761; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6763 = 8'h6b == io_state_in_13 ? 8'hd6 : _GEN_6762; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6764 = 8'h6c == io_state_in_13 ? 8'hd8 : _GEN_6763; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6765 = 8'h6d == io_state_in_13 ? 8'hda : _GEN_6764; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6766 = 8'h6e == io_state_in_13 ? 8'hdc : _GEN_6765; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6767 = 8'h6f == io_state_in_13 ? 8'hde : _GEN_6766; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6768 = 8'h70 == io_state_in_13 ? 8'he0 : _GEN_6767; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6769 = 8'h71 == io_state_in_13 ? 8'he2 : _GEN_6768; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6770 = 8'h72 == io_state_in_13 ? 8'he4 : _GEN_6769; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6771 = 8'h73 == io_state_in_13 ? 8'he6 : _GEN_6770; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6772 = 8'h74 == io_state_in_13 ? 8'he8 : _GEN_6771; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6773 = 8'h75 == io_state_in_13 ? 8'hea : _GEN_6772; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6774 = 8'h76 == io_state_in_13 ? 8'hec : _GEN_6773; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6775 = 8'h77 == io_state_in_13 ? 8'hee : _GEN_6774; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6776 = 8'h78 == io_state_in_13 ? 8'hf0 : _GEN_6775; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6777 = 8'h79 == io_state_in_13 ? 8'hf2 : _GEN_6776; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6778 = 8'h7a == io_state_in_13 ? 8'hf4 : _GEN_6777; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6779 = 8'h7b == io_state_in_13 ? 8'hf6 : _GEN_6778; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6780 = 8'h7c == io_state_in_13 ? 8'hf8 : _GEN_6779; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6781 = 8'h7d == io_state_in_13 ? 8'hfa : _GEN_6780; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6782 = 8'h7e == io_state_in_13 ? 8'hfc : _GEN_6781; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6783 = 8'h7f == io_state_in_13 ? 8'hfe : _GEN_6782; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6784 = 8'h80 == io_state_in_13 ? 8'h1b : _GEN_6783; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6785 = 8'h81 == io_state_in_13 ? 8'h19 : _GEN_6784; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6786 = 8'h82 == io_state_in_13 ? 8'h1f : _GEN_6785; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6787 = 8'h83 == io_state_in_13 ? 8'h1d : _GEN_6786; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6788 = 8'h84 == io_state_in_13 ? 8'h13 : _GEN_6787; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6789 = 8'h85 == io_state_in_13 ? 8'h11 : _GEN_6788; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6790 = 8'h86 == io_state_in_13 ? 8'h17 : _GEN_6789; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6791 = 8'h87 == io_state_in_13 ? 8'h15 : _GEN_6790; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6792 = 8'h88 == io_state_in_13 ? 8'hb : _GEN_6791; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6793 = 8'h89 == io_state_in_13 ? 8'h9 : _GEN_6792; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6794 = 8'h8a == io_state_in_13 ? 8'hf : _GEN_6793; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6795 = 8'h8b == io_state_in_13 ? 8'hd : _GEN_6794; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6796 = 8'h8c == io_state_in_13 ? 8'h3 : _GEN_6795; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6797 = 8'h8d == io_state_in_13 ? 8'h1 : _GEN_6796; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6798 = 8'h8e == io_state_in_13 ? 8'h7 : _GEN_6797; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6799 = 8'h8f == io_state_in_13 ? 8'h5 : _GEN_6798; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6800 = 8'h90 == io_state_in_13 ? 8'h3b : _GEN_6799; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6801 = 8'h91 == io_state_in_13 ? 8'h39 : _GEN_6800; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6802 = 8'h92 == io_state_in_13 ? 8'h3f : _GEN_6801; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6803 = 8'h93 == io_state_in_13 ? 8'h3d : _GEN_6802; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6804 = 8'h94 == io_state_in_13 ? 8'h33 : _GEN_6803; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6805 = 8'h95 == io_state_in_13 ? 8'h31 : _GEN_6804; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6806 = 8'h96 == io_state_in_13 ? 8'h37 : _GEN_6805; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6807 = 8'h97 == io_state_in_13 ? 8'h35 : _GEN_6806; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6808 = 8'h98 == io_state_in_13 ? 8'h2b : _GEN_6807; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6809 = 8'h99 == io_state_in_13 ? 8'h29 : _GEN_6808; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6810 = 8'h9a == io_state_in_13 ? 8'h2f : _GEN_6809; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6811 = 8'h9b == io_state_in_13 ? 8'h2d : _GEN_6810; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6812 = 8'h9c == io_state_in_13 ? 8'h23 : _GEN_6811; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6813 = 8'h9d == io_state_in_13 ? 8'h21 : _GEN_6812; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6814 = 8'h9e == io_state_in_13 ? 8'h27 : _GEN_6813; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6815 = 8'h9f == io_state_in_13 ? 8'h25 : _GEN_6814; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6816 = 8'ha0 == io_state_in_13 ? 8'h5b : _GEN_6815; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6817 = 8'ha1 == io_state_in_13 ? 8'h59 : _GEN_6816; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6818 = 8'ha2 == io_state_in_13 ? 8'h5f : _GEN_6817; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6819 = 8'ha3 == io_state_in_13 ? 8'h5d : _GEN_6818; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6820 = 8'ha4 == io_state_in_13 ? 8'h53 : _GEN_6819; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6821 = 8'ha5 == io_state_in_13 ? 8'h51 : _GEN_6820; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6822 = 8'ha6 == io_state_in_13 ? 8'h57 : _GEN_6821; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6823 = 8'ha7 == io_state_in_13 ? 8'h55 : _GEN_6822; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6824 = 8'ha8 == io_state_in_13 ? 8'h4b : _GEN_6823; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6825 = 8'ha9 == io_state_in_13 ? 8'h49 : _GEN_6824; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6826 = 8'haa == io_state_in_13 ? 8'h4f : _GEN_6825; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6827 = 8'hab == io_state_in_13 ? 8'h4d : _GEN_6826; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6828 = 8'hac == io_state_in_13 ? 8'h43 : _GEN_6827; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6829 = 8'had == io_state_in_13 ? 8'h41 : _GEN_6828; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6830 = 8'hae == io_state_in_13 ? 8'h47 : _GEN_6829; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6831 = 8'haf == io_state_in_13 ? 8'h45 : _GEN_6830; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6832 = 8'hb0 == io_state_in_13 ? 8'h7b : _GEN_6831; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6833 = 8'hb1 == io_state_in_13 ? 8'h79 : _GEN_6832; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6834 = 8'hb2 == io_state_in_13 ? 8'h7f : _GEN_6833; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6835 = 8'hb3 == io_state_in_13 ? 8'h7d : _GEN_6834; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6836 = 8'hb4 == io_state_in_13 ? 8'h73 : _GEN_6835; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6837 = 8'hb5 == io_state_in_13 ? 8'h71 : _GEN_6836; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6838 = 8'hb6 == io_state_in_13 ? 8'h77 : _GEN_6837; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6839 = 8'hb7 == io_state_in_13 ? 8'h75 : _GEN_6838; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6840 = 8'hb8 == io_state_in_13 ? 8'h6b : _GEN_6839; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6841 = 8'hb9 == io_state_in_13 ? 8'h69 : _GEN_6840; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6842 = 8'hba == io_state_in_13 ? 8'h6f : _GEN_6841; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6843 = 8'hbb == io_state_in_13 ? 8'h6d : _GEN_6842; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6844 = 8'hbc == io_state_in_13 ? 8'h63 : _GEN_6843; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6845 = 8'hbd == io_state_in_13 ? 8'h61 : _GEN_6844; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6846 = 8'hbe == io_state_in_13 ? 8'h67 : _GEN_6845; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6847 = 8'hbf == io_state_in_13 ? 8'h65 : _GEN_6846; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6848 = 8'hc0 == io_state_in_13 ? 8'h9b : _GEN_6847; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6849 = 8'hc1 == io_state_in_13 ? 8'h99 : _GEN_6848; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6850 = 8'hc2 == io_state_in_13 ? 8'h9f : _GEN_6849; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6851 = 8'hc3 == io_state_in_13 ? 8'h9d : _GEN_6850; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6852 = 8'hc4 == io_state_in_13 ? 8'h93 : _GEN_6851; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6853 = 8'hc5 == io_state_in_13 ? 8'h91 : _GEN_6852; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6854 = 8'hc6 == io_state_in_13 ? 8'h97 : _GEN_6853; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6855 = 8'hc7 == io_state_in_13 ? 8'h95 : _GEN_6854; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6856 = 8'hc8 == io_state_in_13 ? 8'h8b : _GEN_6855; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6857 = 8'hc9 == io_state_in_13 ? 8'h89 : _GEN_6856; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6858 = 8'hca == io_state_in_13 ? 8'h8f : _GEN_6857; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6859 = 8'hcb == io_state_in_13 ? 8'h8d : _GEN_6858; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6860 = 8'hcc == io_state_in_13 ? 8'h83 : _GEN_6859; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6861 = 8'hcd == io_state_in_13 ? 8'h81 : _GEN_6860; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6862 = 8'hce == io_state_in_13 ? 8'h87 : _GEN_6861; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6863 = 8'hcf == io_state_in_13 ? 8'h85 : _GEN_6862; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6864 = 8'hd0 == io_state_in_13 ? 8'hbb : _GEN_6863; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6865 = 8'hd1 == io_state_in_13 ? 8'hb9 : _GEN_6864; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6866 = 8'hd2 == io_state_in_13 ? 8'hbf : _GEN_6865; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6867 = 8'hd3 == io_state_in_13 ? 8'hbd : _GEN_6866; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6868 = 8'hd4 == io_state_in_13 ? 8'hb3 : _GEN_6867; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6869 = 8'hd5 == io_state_in_13 ? 8'hb1 : _GEN_6868; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6870 = 8'hd6 == io_state_in_13 ? 8'hb7 : _GEN_6869; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6871 = 8'hd7 == io_state_in_13 ? 8'hb5 : _GEN_6870; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6872 = 8'hd8 == io_state_in_13 ? 8'hab : _GEN_6871; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6873 = 8'hd9 == io_state_in_13 ? 8'ha9 : _GEN_6872; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6874 = 8'hda == io_state_in_13 ? 8'haf : _GEN_6873; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6875 = 8'hdb == io_state_in_13 ? 8'had : _GEN_6874; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6876 = 8'hdc == io_state_in_13 ? 8'ha3 : _GEN_6875; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6877 = 8'hdd == io_state_in_13 ? 8'ha1 : _GEN_6876; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6878 = 8'hde == io_state_in_13 ? 8'ha7 : _GEN_6877; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6879 = 8'hdf == io_state_in_13 ? 8'ha5 : _GEN_6878; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6880 = 8'he0 == io_state_in_13 ? 8'hdb : _GEN_6879; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6881 = 8'he1 == io_state_in_13 ? 8'hd9 : _GEN_6880; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6882 = 8'he2 == io_state_in_13 ? 8'hdf : _GEN_6881; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6883 = 8'he3 == io_state_in_13 ? 8'hdd : _GEN_6882; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6884 = 8'he4 == io_state_in_13 ? 8'hd3 : _GEN_6883; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6885 = 8'he5 == io_state_in_13 ? 8'hd1 : _GEN_6884; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6886 = 8'he6 == io_state_in_13 ? 8'hd7 : _GEN_6885; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6887 = 8'he7 == io_state_in_13 ? 8'hd5 : _GEN_6886; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6888 = 8'he8 == io_state_in_13 ? 8'hcb : _GEN_6887; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6889 = 8'he9 == io_state_in_13 ? 8'hc9 : _GEN_6888; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6890 = 8'hea == io_state_in_13 ? 8'hcf : _GEN_6889; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6891 = 8'heb == io_state_in_13 ? 8'hcd : _GEN_6890; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6892 = 8'hec == io_state_in_13 ? 8'hc3 : _GEN_6891; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6893 = 8'hed == io_state_in_13 ? 8'hc1 : _GEN_6892; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6894 = 8'hee == io_state_in_13 ? 8'hc7 : _GEN_6893; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6895 = 8'hef == io_state_in_13 ? 8'hc5 : _GEN_6894; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6896 = 8'hf0 == io_state_in_13 ? 8'hfb : _GEN_6895; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6897 = 8'hf1 == io_state_in_13 ? 8'hf9 : _GEN_6896; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6898 = 8'hf2 == io_state_in_13 ? 8'hff : _GEN_6897; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6899 = 8'hf3 == io_state_in_13 ? 8'hfd : _GEN_6898; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6900 = 8'hf4 == io_state_in_13 ? 8'hf3 : _GEN_6899; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6901 = 8'hf5 == io_state_in_13 ? 8'hf1 : _GEN_6900; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6902 = 8'hf6 == io_state_in_13 ? 8'hf7 : _GEN_6901; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6903 = 8'hf7 == io_state_in_13 ? 8'hf5 : _GEN_6902; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6904 = 8'hf8 == io_state_in_13 ? 8'heb : _GEN_6903; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6905 = 8'hf9 == io_state_in_13 ? 8'he9 : _GEN_6904; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6906 = 8'hfa == io_state_in_13 ? 8'hef : _GEN_6905; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6907 = 8'hfb == io_state_in_13 ? 8'hed : _GEN_6906; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6908 = 8'hfc == io_state_in_13 ? 8'he3 : _GEN_6907; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6909 = 8'hfd == io_state_in_13 ? 8'he1 : _GEN_6908; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6910 = 8'hfe == io_state_in_13 ? 8'he7 : _GEN_6909; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _GEN_6911 = 8'hff == io_state_in_13 ? 8'he5 : _GEN_6910; // @[MixColumns.scala 141:{36,36}]
  wire [7:0] _tmp_state_13_T = io_state_in_12 ^ _GEN_6911; // @[MixColumns.scala 141:36]
  wire [7:0] _GEN_6913 = 8'h1 == io_state_in_14 ? 8'h3 : 8'h0; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6914 = 8'h2 == io_state_in_14 ? 8'h6 : _GEN_6913; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6915 = 8'h3 == io_state_in_14 ? 8'h5 : _GEN_6914; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6916 = 8'h4 == io_state_in_14 ? 8'hc : _GEN_6915; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6917 = 8'h5 == io_state_in_14 ? 8'hf : _GEN_6916; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6918 = 8'h6 == io_state_in_14 ? 8'ha : _GEN_6917; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6919 = 8'h7 == io_state_in_14 ? 8'h9 : _GEN_6918; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6920 = 8'h8 == io_state_in_14 ? 8'h18 : _GEN_6919; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6921 = 8'h9 == io_state_in_14 ? 8'h1b : _GEN_6920; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6922 = 8'ha == io_state_in_14 ? 8'h1e : _GEN_6921; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6923 = 8'hb == io_state_in_14 ? 8'h1d : _GEN_6922; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6924 = 8'hc == io_state_in_14 ? 8'h14 : _GEN_6923; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6925 = 8'hd == io_state_in_14 ? 8'h17 : _GEN_6924; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6926 = 8'he == io_state_in_14 ? 8'h12 : _GEN_6925; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6927 = 8'hf == io_state_in_14 ? 8'h11 : _GEN_6926; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6928 = 8'h10 == io_state_in_14 ? 8'h30 : _GEN_6927; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6929 = 8'h11 == io_state_in_14 ? 8'h33 : _GEN_6928; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6930 = 8'h12 == io_state_in_14 ? 8'h36 : _GEN_6929; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6931 = 8'h13 == io_state_in_14 ? 8'h35 : _GEN_6930; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6932 = 8'h14 == io_state_in_14 ? 8'h3c : _GEN_6931; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6933 = 8'h15 == io_state_in_14 ? 8'h3f : _GEN_6932; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6934 = 8'h16 == io_state_in_14 ? 8'h3a : _GEN_6933; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6935 = 8'h17 == io_state_in_14 ? 8'h39 : _GEN_6934; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6936 = 8'h18 == io_state_in_14 ? 8'h28 : _GEN_6935; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6937 = 8'h19 == io_state_in_14 ? 8'h2b : _GEN_6936; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6938 = 8'h1a == io_state_in_14 ? 8'h2e : _GEN_6937; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6939 = 8'h1b == io_state_in_14 ? 8'h2d : _GEN_6938; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6940 = 8'h1c == io_state_in_14 ? 8'h24 : _GEN_6939; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6941 = 8'h1d == io_state_in_14 ? 8'h27 : _GEN_6940; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6942 = 8'h1e == io_state_in_14 ? 8'h22 : _GEN_6941; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6943 = 8'h1f == io_state_in_14 ? 8'h21 : _GEN_6942; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6944 = 8'h20 == io_state_in_14 ? 8'h60 : _GEN_6943; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6945 = 8'h21 == io_state_in_14 ? 8'h63 : _GEN_6944; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6946 = 8'h22 == io_state_in_14 ? 8'h66 : _GEN_6945; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6947 = 8'h23 == io_state_in_14 ? 8'h65 : _GEN_6946; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6948 = 8'h24 == io_state_in_14 ? 8'h6c : _GEN_6947; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6949 = 8'h25 == io_state_in_14 ? 8'h6f : _GEN_6948; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6950 = 8'h26 == io_state_in_14 ? 8'h6a : _GEN_6949; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6951 = 8'h27 == io_state_in_14 ? 8'h69 : _GEN_6950; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6952 = 8'h28 == io_state_in_14 ? 8'h78 : _GEN_6951; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6953 = 8'h29 == io_state_in_14 ? 8'h7b : _GEN_6952; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6954 = 8'h2a == io_state_in_14 ? 8'h7e : _GEN_6953; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6955 = 8'h2b == io_state_in_14 ? 8'h7d : _GEN_6954; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6956 = 8'h2c == io_state_in_14 ? 8'h74 : _GEN_6955; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6957 = 8'h2d == io_state_in_14 ? 8'h77 : _GEN_6956; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6958 = 8'h2e == io_state_in_14 ? 8'h72 : _GEN_6957; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6959 = 8'h2f == io_state_in_14 ? 8'h71 : _GEN_6958; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6960 = 8'h30 == io_state_in_14 ? 8'h50 : _GEN_6959; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6961 = 8'h31 == io_state_in_14 ? 8'h53 : _GEN_6960; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6962 = 8'h32 == io_state_in_14 ? 8'h56 : _GEN_6961; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6963 = 8'h33 == io_state_in_14 ? 8'h55 : _GEN_6962; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6964 = 8'h34 == io_state_in_14 ? 8'h5c : _GEN_6963; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6965 = 8'h35 == io_state_in_14 ? 8'h5f : _GEN_6964; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6966 = 8'h36 == io_state_in_14 ? 8'h5a : _GEN_6965; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6967 = 8'h37 == io_state_in_14 ? 8'h59 : _GEN_6966; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6968 = 8'h38 == io_state_in_14 ? 8'h48 : _GEN_6967; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6969 = 8'h39 == io_state_in_14 ? 8'h4b : _GEN_6968; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6970 = 8'h3a == io_state_in_14 ? 8'h4e : _GEN_6969; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6971 = 8'h3b == io_state_in_14 ? 8'h4d : _GEN_6970; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6972 = 8'h3c == io_state_in_14 ? 8'h44 : _GEN_6971; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6973 = 8'h3d == io_state_in_14 ? 8'h47 : _GEN_6972; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6974 = 8'h3e == io_state_in_14 ? 8'h42 : _GEN_6973; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6975 = 8'h3f == io_state_in_14 ? 8'h41 : _GEN_6974; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6976 = 8'h40 == io_state_in_14 ? 8'hc0 : _GEN_6975; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6977 = 8'h41 == io_state_in_14 ? 8'hc3 : _GEN_6976; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6978 = 8'h42 == io_state_in_14 ? 8'hc6 : _GEN_6977; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6979 = 8'h43 == io_state_in_14 ? 8'hc5 : _GEN_6978; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6980 = 8'h44 == io_state_in_14 ? 8'hcc : _GEN_6979; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6981 = 8'h45 == io_state_in_14 ? 8'hcf : _GEN_6980; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6982 = 8'h46 == io_state_in_14 ? 8'hca : _GEN_6981; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6983 = 8'h47 == io_state_in_14 ? 8'hc9 : _GEN_6982; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6984 = 8'h48 == io_state_in_14 ? 8'hd8 : _GEN_6983; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6985 = 8'h49 == io_state_in_14 ? 8'hdb : _GEN_6984; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6986 = 8'h4a == io_state_in_14 ? 8'hde : _GEN_6985; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6987 = 8'h4b == io_state_in_14 ? 8'hdd : _GEN_6986; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6988 = 8'h4c == io_state_in_14 ? 8'hd4 : _GEN_6987; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6989 = 8'h4d == io_state_in_14 ? 8'hd7 : _GEN_6988; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6990 = 8'h4e == io_state_in_14 ? 8'hd2 : _GEN_6989; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6991 = 8'h4f == io_state_in_14 ? 8'hd1 : _GEN_6990; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6992 = 8'h50 == io_state_in_14 ? 8'hf0 : _GEN_6991; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6993 = 8'h51 == io_state_in_14 ? 8'hf3 : _GEN_6992; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6994 = 8'h52 == io_state_in_14 ? 8'hf6 : _GEN_6993; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6995 = 8'h53 == io_state_in_14 ? 8'hf5 : _GEN_6994; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6996 = 8'h54 == io_state_in_14 ? 8'hfc : _GEN_6995; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6997 = 8'h55 == io_state_in_14 ? 8'hff : _GEN_6996; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6998 = 8'h56 == io_state_in_14 ? 8'hfa : _GEN_6997; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_6999 = 8'h57 == io_state_in_14 ? 8'hf9 : _GEN_6998; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7000 = 8'h58 == io_state_in_14 ? 8'he8 : _GEN_6999; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7001 = 8'h59 == io_state_in_14 ? 8'heb : _GEN_7000; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7002 = 8'h5a == io_state_in_14 ? 8'hee : _GEN_7001; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7003 = 8'h5b == io_state_in_14 ? 8'hed : _GEN_7002; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7004 = 8'h5c == io_state_in_14 ? 8'he4 : _GEN_7003; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7005 = 8'h5d == io_state_in_14 ? 8'he7 : _GEN_7004; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7006 = 8'h5e == io_state_in_14 ? 8'he2 : _GEN_7005; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7007 = 8'h5f == io_state_in_14 ? 8'he1 : _GEN_7006; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7008 = 8'h60 == io_state_in_14 ? 8'ha0 : _GEN_7007; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7009 = 8'h61 == io_state_in_14 ? 8'ha3 : _GEN_7008; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7010 = 8'h62 == io_state_in_14 ? 8'ha6 : _GEN_7009; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7011 = 8'h63 == io_state_in_14 ? 8'ha5 : _GEN_7010; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7012 = 8'h64 == io_state_in_14 ? 8'hac : _GEN_7011; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7013 = 8'h65 == io_state_in_14 ? 8'haf : _GEN_7012; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7014 = 8'h66 == io_state_in_14 ? 8'haa : _GEN_7013; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7015 = 8'h67 == io_state_in_14 ? 8'ha9 : _GEN_7014; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7016 = 8'h68 == io_state_in_14 ? 8'hb8 : _GEN_7015; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7017 = 8'h69 == io_state_in_14 ? 8'hbb : _GEN_7016; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7018 = 8'h6a == io_state_in_14 ? 8'hbe : _GEN_7017; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7019 = 8'h6b == io_state_in_14 ? 8'hbd : _GEN_7018; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7020 = 8'h6c == io_state_in_14 ? 8'hb4 : _GEN_7019; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7021 = 8'h6d == io_state_in_14 ? 8'hb7 : _GEN_7020; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7022 = 8'h6e == io_state_in_14 ? 8'hb2 : _GEN_7021; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7023 = 8'h6f == io_state_in_14 ? 8'hb1 : _GEN_7022; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7024 = 8'h70 == io_state_in_14 ? 8'h90 : _GEN_7023; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7025 = 8'h71 == io_state_in_14 ? 8'h93 : _GEN_7024; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7026 = 8'h72 == io_state_in_14 ? 8'h96 : _GEN_7025; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7027 = 8'h73 == io_state_in_14 ? 8'h95 : _GEN_7026; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7028 = 8'h74 == io_state_in_14 ? 8'h9c : _GEN_7027; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7029 = 8'h75 == io_state_in_14 ? 8'h9f : _GEN_7028; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7030 = 8'h76 == io_state_in_14 ? 8'h9a : _GEN_7029; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7031 = 8'h77 == io_state_in_14 ? 8'h99 : _GEN_7030; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7032 = 8'h78 == io_state_in_14 ? 8'h88 : _GEN_7031; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7033 = 8'h79 == io_state_in_14 ? 8'h8b : _GEN_7032; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7034 = 8'h7a == io_state_in_14 ? 8'h8e : _GEN_7033; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7035 = 8'h7b == io_state_in_14 ? 8'h8d : _GEN_7034; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7036 = 8'h7c == io_state_in_14 ? 8'h84 : _GEN_7035; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7037 = 8'h7d == io_state_in_14 ? 8'h87 : _GEN_7036; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7038 = 8'h7e == io_state_in_14 ? 8'h82 : _GEN_7037; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7039 = 8'h7f == io_state_in_14 ? 8'h81 : _GEN_7038; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7040 = 8'h80 == io_state_in_14 ? 8'h9b : _GEN_7039; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7041 = 8'h81 == io_state_in_14 ? 8'h98 : _GEN_7040; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7042 = 8'h82 == io_state_in_14 ? 8'h9d : _GEN_7041; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7043 = 8'h83 == io_state_in_14 ? 8'h9e : _GEN_7042; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7044 = 8'h84 == io_state_in_14 ? 8'h97 : _GEN_7043; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7045 = 8'h85 == io_state_in_14 ? 8'h94 : _GEN_7044; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7046 = 8'h86 == io_state_in_14 ? 8'h91 : _GEN_7045; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7047 = 8'h87 == io_state_in_14 ? 8'h92 : _GEN_7046; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7048 = 8'h88 == io_state_in_14 ? 8'h83 : _GEN_7047; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7049 = 8'h89 == io_state_in_14 ? 8'h80 : _GEN_7048; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7050 = 8'h8a == io_state_in_14 ? 8'h85 : _GEN_7049; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7051 = 8'h8b == io_state_in_14 ? 8'h86 : _GEN_7050; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7052 = 8'h8c == io_state_in_14 ? 8'h8f : _GEN_7051; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7053 = 8'h8d == io_state_in_14 ? 8'h8c : _GEN_7052; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7054 = 8'h8e == io_state_in_14 ? 8'h89 : _GEN_7053; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7055 = 8'h8f == io_state_in_14 ? 8'h8a : _GEN_7054; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7056 = 8'h90 == io_state_in_14 ? 8'hab : _GEN_7055; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7057 = 8'h91 == io_state_in_14 ? 8'ha8 : _GEN_7056; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7058 = 8'h92 == io_state_in_14 ? 8'had : _GEN_7057; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7059 = 8'h93 == io_state_in_14 ? 8'hae : _GEN_7058; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7060 = 8'h94 == io_state_in_14 ? 8'ha7 : _GEN_7059; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7061 = 8'h95 == io_state_in_14 ? 8'ha4 : _GEN_7060; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7062 = 8'h96 == io_state_in_14 ? 8'ha1 : _GEN_7061; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7063 = 8'h97 == io_state_in_14 ? 8'ha2 : _GEN_7062; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7064 = 8'h98 == io_state_in_14 ? 8'hb3 : _GEN_7063; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7065 = 8'h99 == io_state_in_14 ? 8'hb0 : _GEN_7064; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7066 = 8'h9a == io_state_in_14 ? 8'hb5 : _GEN_7065; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7067 = 8'h9b == io_state_in_14 ? 8'hb6 : _GEN_7066; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7068 = 8'h9c == io_state_in_14 ? 8'hbf : _GEN_7067; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7069 = 8'h9d == io_state_in_14 ? 8'hbc : _GEN_7068; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7070 = 8'h9e == io_state_in_14 ? 8'hb9 : _GEN_7069; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7071 = 8'h9f == io_state_in_14 ? 8'hba : _GEN_7070; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7072 = 8'ha0 == io_state_in_14 ? 8'hfb : _GEN_7071; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7073 = 8'ha1 == io_state_in_14 ? 8'hf8 : _GEN_7072; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7074 = 8'ha2 == io_state_in_14 ? 8'hfd : _GEN_7073; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7075 = 8'ha3 == io_state_in_14 ? 8'hfe : _GEN_7074; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7076 = 8'ha4 == io_state_in_14 ? 8'hf7 : _GEN_7075; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7077 = 8'ha5 == io_state_in_14 ? 8'hf4 : _GEN_7076; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7078 = 8'ha6 == io_state_in_14 ? 8'hf1 : _GEN_7077; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7079 = 8'ha7 == io_state_in_14 ? 8'hf2 : _GEN_7078; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7080 = 8'ha8 == io_state_in_14 ? 8'he3 : _GEN_7079; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7081 = 8'ha9 == io_state_in_14 ? 8'he0 : _GEN_7080; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7082 = 8'haa == io_state_in_14 ? 8'he5 : _GEN_7081; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7083 = 8'hab == io_state_in_14 ? 8'he6 : _GEN_7082; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7084 = 8'hac == io_state_in_14 ? 8'hef : _GEN_7083; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7085 = 8'had == io_state_in_14 ? 8'hec : _GEN_7084; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7086 = 8'hae == io_state_in_14 ? 8'he9 : _GEN_7085; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7087 = 8'haf == io_state_in_14 ? 8'hea : _GEN_7086; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7088 = 8'hb0 == io_state_in_14 ? 8'hcb : _GEN_7087; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7089 = 8'hb1 == io_state_in_14 ? 8'hc8 : _GEN_7088; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7090 = 8'hb2 == io_state_in_14 ? 8'hcd : _GEN_7089; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7091 = 8'hb3 == io_state_in_14 ? 8'hce : _GEN_7090; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7092 = 8'hb4 == io_state_in_14 ? 8'hc7 : _GEN_7091; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7093 = 8'hb5 == io_state_in_14 ? 8'hc4 : _GEN_7092; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7094 = 8'hb6 == io_state_in_14 ? 8'hc1 : _GEN_7093; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7095 = 8'hb7 == io_state_in_14 ? 8'hc2 : _GEN_7094; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7096 = 8'hb8 == io_state_in_14 ? 8'hd3 : _GEN_7095; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7097 = 8'hb9 == io_state_in_14 ? 8'hd0 : _GEN_7096; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7098 = 8'hba == io_state_in_14 ? 8'hd5 : _GEN_7097; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7099 = 8'hbb == io_state_in_14 ? 8'hd6 : _GEN_7098; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7100 = 8'hbc == io_state_in_14 ? 8'hdf : _GEN_7099; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7101 = 8'hbd == io_state_in_14 ? 8'hdc : _GEN_7100; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7102 = 8'hbe == io_state_in_14 ? 8'hd9 : _GEN_7101; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7103 = 8'hbf == io_state_in_14 ? 8'hda : _GEN_7102; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7104 = 8'hc0 == io_state_in_14 ? 8'h5b : _GEN_7103; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7105 = 8'hc1 == io_state_in_14 ? 8'h58 : _GEN_7104; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7106 = 8'hc2 == io_state_in_14 ? 8'h5d : _GEN_7105; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7107 = 8'hc3 == io_state_in_14 ? 8'h5e : _GEN_7106; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7108 = 8'hc4 == io_state_in_14 ? 8'h57 : _GEN_7107; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7109 = 8'hc5 == io_state_in_14 ? 8'h54 : _GEN_7108; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7110 = 8'hc6 == io_state_in_14 ? 8'h51 : _GEN_7109; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7111 = 8'hc7 == io_state_in_14 ? 8'h52 : _GEN_7110; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7112 = 8'hc8 == io_state_in_14 ? 8'h43 : _GEN_7111; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7113 = 8'hc9 == io_state_in_14 ? 8'h40 : _GEN_7112; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7114 = 8'hca == io_state_in_14 ? 8'h45 : _GEN_7113; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7115 = 8'hcb == io_state_in_14 ? 8'h46 : _GEN_7114; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7116 = 8'hcc == io_state_in_14 ? 8'h4f : _GEN_7115; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7117 = 8'hcd == io_state_in_14 ? 8'h4c : _GEN_7116; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7118 = 8'hce == io_state_in_14 ? 8'h49 : _GEN_7117; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7119 = 8'hcf == io_state_in_14 ? 8'h4a : _GEN_7118; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7120 = 8'hd0 == io_state_in_14 ? 8'h6b : _GEN_7119; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7121 = 8'hd1 == io_state_in_14 ? 8'h68 : _GEN_7120; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7122 = 8'hd2 == io_state_in_14 ? 8'h6d : _GEN_7121; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7123 = 8'hd3 == io_state_in_14 ? 8'h6e : _GEN_7122; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7124 = 8'hd4 == io_state_in_14 ? 8'h67 : _GEN_7123; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7125 = 8'hd5 == io_state_in_14 ? 8'h64 : _GEN_7124; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7126 = 8'hd6 == io_state_in_14 ? 8'h61 : _GEN_7125; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7127 = 8'hd7 == io_state_in_14 ? 8'h62 : _GEN_7126; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7128 = 8'hd8 == io_state_in_14 ? 8'h73 : _GEN_7127; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7129 = 8'hd9 == io_state_in_14 ? 8'h70 : _GEN_7128; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7130 = 8'hda == io_state_in_14 ? 8'h75 : _GEN_7129; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7131 = 8'hdb == io_state_in_14 ? 8'h76 : _GEN_7130; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7132 = 8'hdc == io_state_in_14 ? 8'h7f : _GEN_7131; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7133 = 8'hdd == io_state_in_14 ? 8'h7c : _GEN_7132; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7134 = 8'hde == io_state_in_14 ? 8'h79 : _GEN_7133; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7135 = 8'hdf == io_state_in_14 ? 8'h7a : _GEN_7134; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7136 = 8'he0 == io_state_in_14 ? 8'h3b : _GEN_7135; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7137 = 8'he1 == io_state_in_14 ? 8'h38 : _GEN_7136; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7138 = 8'he2 == io_state_in_14 ? 8'h3d : _GEN_7137; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7139 = 8'he3 == io_state_in_14 ? 8'h3e : _GEN_7138; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7140 = 8'he4 == io_state_in_14 ? 8'h37 : _GEN_7139; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7141 = 8'he5 == io_state_in_14 ? 8'h34 : _GEN_7140; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7142 = 8'he6 == io_state_in_14 ? 8'h31 : _GEN_7141; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7143 = 8'he7 == io_state_in_14 ? 8'h32 : _GEN_7142; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7144 = 8'he8 == io_state_in_14 ? 8'h23 : _GEN_7143; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7145 = 8'he9 == io_state_in_14 ? 8'h20 : _GEN_7144; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7146 = 8'hea == io_state_in_14 ? 8'h25 : _GEN_7145; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7147 = 8'heb == io_state_in_14 ? 8'h26 : _GEN_7146; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7148 = 8'hec == io_state_in_14 ? 8'h2f : _GEN_7147; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7149 = 8'hed == io_state_in_14 ? 8'h2c : _GEN_7148; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7150 = 8'hee == io_state_in_14 ? 8'h29 : _GEN_7149; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7151 = 8'hef == io_state_in_14 ? 8'h2a : _GEN_7150; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7152 = 8'hf0 == io_state_in_14 ? 8'hb : _GEN_7151; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7153 = 8'hf1 == io_state_in_14 ? 8'h8 : _GEN_7152; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7154 = 8'hf2 == io_state_in_14 ? 8'hd : _GEN_7153; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7155 = 8'hf3 == io_state_in_14 ? 8'he : _GEN_7154; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7156 = 8'hf4 == io_state_in_14 ? 8'h7 : _GEN_7155; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7157 = 8'hf5 == io_state_in_14 ? 8'h4 : _GEN_7156; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7158 = 8'hf6 == io_state_in_14 ? 8'h1 : _GEN_7157; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7159 = 8'hf7 == io_state_in_14 ? 8'h2 : _GEN_7158; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7160 = 8'hf8 == io_state_in_14 ? 8'h13 : _GEN_7159; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7161 = 8'hf9 == io_state_in_14 ? 8'h10 : _GEN_7160; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7162 = 8'hfa == io_state_in_14 ? 8'h15 : _GEN_7161; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7163 = 8'hfb == io_state_in_14 ? 8'h16 : _GEN_7162; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7164 = 8'hfc == io_state_in_14 ? 8'h1f : _GEN_7163; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7165 = 8'hfd == io_state_in_14 ? 8'h1c : _GEN_7164; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7166 = 8'hfe == io_state_in_14 ? 8'h19 : _GEN_7165; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _GEN_7167 = 8'hff == io_state_in_14 ? 8'h1a : _GEN_7166; // @[MixColumns.scala 141:{61,61}]
  wire [7:0] _tmp_state_13_T_1 = _tmp_state_13_T ^ _GEN_7167; // @[MixColumns.scala 141:61]
  wire [7:0] _tmp_state_14_T = io_state_in_12 ^ io_state_in_13; // @[MixColumns.scala 142:36]
  wire [7:0] _GEN_7169 = 8'h1 == io_state_in_14 ? 8'h2 : 8'h0; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7170 = 8'h2 == io_state_in_14 ? 8'h4 : _GEN_7169; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7171 = 8'h3 == io_state_in_14 ? 8'h6 : _GEN_7170; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7172 = 8'h4 == io_state_in_14 ? 8'h8 : _GEN_7171; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7173 = 8'h5 == io_state_in_14 ? 8'ha : _GEN_7172; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7174 = 8'h6 == io_state_in_14 ? 8'hc : _GEN_7173; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7175 = 8'h7 == io_state_in_14 ? 8'he : _GEN_7174; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7176 = 8'h8 == io_state_in_14 ? 8'h10 : _GEN_7175; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7177 = 8'h9 == io_state_in_14 ? 8'h12 : _GEN_7176; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7178 = 8'ha == io_state_in_14 ? 8'h14 : _GEN_7177; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7179 = 8'hb == io_state_in_14 ? 8'h16 : _GEN_7178; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7180 = 8'hc == io_state_in_14 ? 8'h18 : _GEN_7179; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7181 = 8'hd == io_state_in_14 ? 8'h1a : _GEN_7180; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7182 = 8'he == io_state_in_14 ? 8'h1c : _GEN_7181; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7183 = 8'hf == io_state_in_14 ? 8'h1e : _GEN_7182; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7184 = 8'h10 == io_state_in_14 ? 8'h20 : _GEN_7183; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7185 = 8'h11 == io_state_in_14 ? 8'h22 : _GEN_7184; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7186 = 8'h12 == io_state_in_14 ? 8'h24 : _GEN_7185; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7187 = 8'h13 == io_state_in_14 ? 8'h26 : _GEN_7186; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7188 = 8'h14 == io_state_in_14 ? 8'h28 : _GEN_7187; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7189 = 8'h15 == io_state_in_14 ? 8'h2a : _GEN_7188; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7190 = 8'h16 == io_state_in_14 ? 8'h2c : _GEN_7189; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7191 = 8'h17 == io_state_in_14 ? 8'h2e : _GEN_7190; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7192 = 8'h18 == io_state_in_14 ? 8'h30 : _GEN_7191; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7193 = 8'h19 == io_state_in_14 ? 8'h32 : _GEN_7192; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7194 = 8'h1a == io_state_in_14 ? 8'h34 : _GEN_7193; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7195 = 8'h1b == io_state_in_14 ? 8'h36 : _GEN_7194; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7196 = 8'h1c == io_state_in_14 ? 8'h38 : _GEN_7195; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7197 = 8'h1d == io_state_in_14 ? 8'h3a : _GEN_7196; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7198 = 8'h1e == io_state_in_14 ? 8'h3c : _GEN_7197; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7199 = 8'h1f == io_state_in_14 ? 8'h3e : _GEN_7198; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7200 = 8'h20 == io_state_in_14 ? 8'h40 : _GEN_7199; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7201 = 8'h21 == io_state_in_14 ? 8'h42 : _GEN_7200; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7202 = 8'h22 == io_state_in_14 ? 8'h44 : _GEN_7201; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7203 = 8'h23 == io_state_in_14 ? 8'h46 : _GEN_7202; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7204 = 8'h24 == io_state_in_14 ? 8'h48 : _GEN_7203; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7205 = 8'h25 == io_state_in_14 ? 8'h4a : _GEN_7204; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7206 = 8'h26 == io_state_in_14 ? 8'h4c : _GEN_7205; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7207 = 8'h27 == io_state_in_14 ? 8'h4e : _GEN_7206; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7208 = 8'h28 == io_state_in_14 ? 8'h50 : _GEN_7207; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7209 = 8'h29 == io_state_in_14 ? 8'h52 : _GEN_7208; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7210 = 8'h2a == io_state_in_14 ? 8'h54 : _GEN_7209; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7211 = 8'h2b == io_state_in_14 ? 8'h56 : _GEN_7210; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7212 = 8'h2c == io_state_in_14 ? 8'h58 : _GEN_7211; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7213 = 8'h2d == io_state_in_14 ? 8'h5a : _GEN_7212; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7214 = 8'h2e == io_state_in_14 ? 8'h5c : _GEN_7213; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7215 = 8'h2f == io_state_in_14 ? 8'h5e : _GEN_7214; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7216 = 8'h30 == io_state_in_14 ? 8'h60 : _GEN_7215; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7217 = 8'h31 == io_state_in_14 ? 8'h62 : _GEN_7216; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7218 = 8'h32 == io_state_in_14 ? 8'h64 : _GEN_7217; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7219 = 8'h33 == io_state_in_14 ? 8'h66 : _GEN_7218; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7220 = 8'h34 == io_state_in_14 ? 8'h68 : _GEN_7219; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7221 = 8'h35 == io_state_in_14 ? 8'h6a : _GEN_7220; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7222 = 8'h36 == io_state_in_14 ? 8'h6c : _GEN_7221; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7223 = 8'h37 == io_state_in_14 ? 8'h6e : _GEN_7222; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7224 = 8'h38 == io_state_in_14 ? 8'h70 : _GEN_7223; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7225 = 8'h39 == io_state_in_14 ? 8'h72 : _GEN_7224; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7226 = 8'h3a == io_state_in_14 ? 8'h74 : _GEN_7225; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7227 = 8'h3b == io_state_in_14 ? 8'h76 : _GEN_7226; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7228 = 8'h3c == io_state_in_14 ? 8'h78 : _GEN_7227; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7229 = 8'h3d == io_state_in_14 ? 8'h7a : _GEN_7228; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7230 = 8'h3e == io_state_in_14 ? 8'h7c : _GEN_7229; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7231 = 8'h3f == io_state_in_14 ? 8'h7e : _GEN_7230; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7232 = 8'h40 == io_state_in_14 ? 8'h80 : _GEN_7231; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7233 = 8'h41 == io_state_in_14 ? 8'h82 : _GEN_7232; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7234 = 8'h42 == io_state_in_14 ? 8'h84 : _GEN_7233; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7235 = 8'h43 == io_state_in_14 ? 8'h86 : _GEN_7234; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7236 = 8'h44 == io_state_in_14 ? 8'h88 : _GEN_7235; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7237 = 8'h45 == io_state_in_14 ? 8'h8a : _GEN_7236; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7238 = 8'h46 == io_state_in_14 ? 8'h8c : _GEN_7237; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7239 = 8'h47 == io_state_in_14 ? 8'h8e : _GEN_7238; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7240 = 8'h48 == io_state_in_14 ? 8'h90 : _GEN_7239; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7241 = 8'h49 == io_state_in_14 ? 8'h92 : _GEN_7240; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7242 = 8'h4a == io_state_in_14 ? 8'h94 : _GEN_7241; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7243 = 8'h4b == io_state_in_14 ? 8'h96 : _GEN_7242; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7244 = 8'h4c == io_state_in_14 ? 8'h98 : _GEN_7243; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7245 = 8'h4d == io_state_in_14 ? 8'h9a : _GEN_7244; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7246 = 8'h4e == io_state_in_14 ? 8'h9c : _GEN_7245; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7247 = 8'h4f == io_state_in_14 ? 8'h9e : _GEN_7246; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7248 = 8'h50 == io_state_in_14 ? 8'ha0 : _GEN_7247; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7249 = 8'h51 == io_state_in_14 ? 8'ha2 : _GEN_7248; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7250 = 8'h52 == io_state_in_14 ? 8'ha4 : _GEN_7249; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7251 = 8'h53 == io_state_in_14 ? 8'ha6 : _GEN_7250; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7252 = 8'h54 == io_state_in_14 ? 8'ha8 : _GEN_7251; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7253 = 8'h55 == io_state_in_14 ? 8'haa : _GEN_7252; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7254 = 8'h56 == io_state_in_14 ? 8'hac : _GEN_7253; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7255 = 8'h57 == io_state_in_14 ? 8'hae : _GEN_7254; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7256 = 8'h58 == io_state_in_14 ? 8'hb0 : _GEN_7255; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7257 = 8'h59 == io_state_in_14 ? 8'hb2 : _GEN_7256; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7258 = 8'h5a == io_state_in_14 ? 8'hb4 : _GEN_7257; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7259 = 8'h5b == io_state_in_14 ? 8'hb6 : _GEN_7258; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7260 = 8'h5c == io_state_in_14 ? 8'hb8 : _GEN_7259; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7261 = 8'h5d == io_state_in_14 ? 8'hba : _GEN_7260; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7262 = 8'h5e == io_state_in_14 ? 8'hbc : _GEN_7261; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7263 = 8'h5f == io_state_in_14 ? 8'hbe : _GEN_7262; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7264 = 8'h60 == io_state_in_14 ? 8'hc0 : _GEN_7263; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7265 = 8'h61 == io_state_in_14 ? 8'hc2 : _GEN_7264; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7266 = 8'h62 == io_state_in_14 ? 8'hc4 : _GEN_7265; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7267 = 8'h63 == io_state_in_14 ? 8'hc6 : _GEN_7266; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7268 = 8'h64 == io_state_in_14 ? 8'hc8 : _GEN_7267; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7269 = 8'h65 == io_state_in_14 ? 8'hca : _GEN_7268; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7270 = 8'h66 == io_state_in_14 ? 8'hcc : _GEN_7269; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7271 = 8'h67 == io_state_in_14 ? 8'hce : _GEN_7270; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7272 = 8'h68 == io_state_in_14 ? 8'hd0 : _GEN_7271; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7273 = 8'h69 == io_state_in_14 ? 8'hd2 : _GEN_7272; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7274 = 8'h6a == io_state_in_14 ? 8'hd4 : _GEN_7273; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7275 = 8'h6b == io_state_in_14 ? 8'hd6 : _GEN_7274; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7276 = 8'h6c == io_state_in_14 ? 8'hd8 : _GEN_7275; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7277 = 8'h6d == io_state_in_14 ? 8'hda : _GEN_7276; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7278 = 8'h6e == io_state_in_14 ? 8'hdc : _GEN_7277; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7279 = 8'h6f == io_state_in_14 ? 8'hde : _GEN_7278; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7280 = 8'h70 == io_state_in_14 ? 8'he0 : _GEN_7279; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7281 = 8'h71 == io_state_in_14 ? 8'he2 : _GEN_7280; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7282 = 8'h72 == io_state_in_14 ? 8'he4 : _GEN_7281; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7283 = 8'h73 == io_state_in_14 ? 8'he6 : _GEN_7282; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7284 = 8'h74 == io_state_in_14 ? 8'he8 : _GEN_7283; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7285 = 8'h75 == io_state_in_14 ? 8'hea : _GEN_7284; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7286 = 8'h76 == io_state_in_14 ? 8'hec : _GEN_7285; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7287 = 8'h77 == io_state_in_14 ? 8'hee : _GEN_7286; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7288 = 8'h78 == io_state_in_14 ? 8'hf0 : _GEN_7287; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7289 = 8'h79 == io_state_in_14 ? 8'hf2 : _GEN_7288; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7290 = 8'h7a == io_state_in_14 ? 8'hf4 : _GEN_7289; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7291 = 8'h7b == io_state_in_14 ? 8'hf6 : _GEN_7290; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7292 = 8'h7c == io_state_in_14 ? 8'hf8 : _GEN_7291; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7293 = 8'h7d == io_state_in_14 ? 8'hfa : _GEN_7292; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7294 = 8'h7e == io_state_in_14 ? 8'hfc : _GEN_7293; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7295 = 8'h7f == io_state_in_14 ? 8'hfe : _GEN_7294; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7296 = 8'h80 == io_state_in_14 ? 8'h1b : _GEN_7295; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7297 = 8'h81 == io_state_in_14 ? 8'h19 : _GEN_7296; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7298 = 8'h82 == io_state_in_14 ? 8'h1f : _GEN_7297; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7299 = 8'h83 == io_state_in_14 ? 8'h1d : _GEN_7298; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7300 = 8'h84 == io_state_in_14 ? 8'h13 : _GEN_7299; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7301 = 8'h85 == io_state_in_14 ? 8'h11 : _GEN_7300; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7302 = 8'h86 == io_state_in_14 ? 8'h17 : _GEN_7301; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7303 = 8'h87 == io_state_in_14 ? 8'h15 : _GEN_7302; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7304 = 8'h88 == io_state_in_14 ? 8'hb : _GEN_7303; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7305 = 8'h89 == io_state_in_14 ? 8'h9 : _GEN_7304; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7306 = 8'h8a == io_state_in_14 ? 8'hf : _GEN_7305; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7307 = 8'h8b == io_state_in_14 ? 8'hd : _GEN_7306; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7308 = 8'h8c == io_state_in_14 ? 8'h3 : _GEN_7307; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7309 = 8'h8d == io_state_in_14 ? 8'h1 : _GEN_7308; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7310 = 8'h8e == io_state_in_14 ? 8'h7 : _GEN_7309; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7311 = 8'h8f == io_state_in_14 ? 8'h5 : _GEN_7310; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7312 = 8'h90 == io_state_in_14 ? 8'h3b : _GEN_7311; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7313 = 8'h91 == io_state_in_14 ? 8'h39 : _GEN_7312; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7314 = 8'h92 == io_state_in_14 ? 8'h3f : _GEN_7313; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7315 = 8'h93 == io_state_in_14 ? 8'h3d : _GEN_7314; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7316 = 8'h94 == io_state_in_14 ? 8'h33 : _GEN_7315; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7317 = 8'h95 == io_state_in_14 ? 8'h31 : _GEN_7316; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7318 = 8'h96 == io_state_in_14 ? 8'h37 : _GEN_7317; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7319 = 8'h97 == io_state_in_14 ? 8'h35 : _GEN_7318; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7320 = 8'h98 == io_state_in_14 ? 8'h2b : _GEN_7319; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7321 = 8'h99 == io_state_in_14 ? 8'h29 : _GEN_7320; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7322 = 8'h9a == io_state_in_14 ? 8'h2f : _GEN_7321; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7323 = 8'h9b == io_state_in_14 ? 8'h2d : _GEN_7322; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7324 = 8'h9c == io_state_in_14 ? 8'h23 : _GEN_7323; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7325 = 8'h9d == io_state_in_14 ? 8'h21 : _GEN_7324; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7326 = 8'h9e == io_state_in_14 ? 8'h27 : _GEN_7325; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7327 = 8'h9f == io_state_in_14 ? 8'h25 : _GEN_7326; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7328 = 8'ha0 == io_state_in_14 ? 8'h5b : _GEN_7327; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7329 = 8'ha1 == io_state_in_14 ? 8'h59 : _GEN_7328; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7330 = 8'ha2 == io_state_in_14 ? 8'h5f : _GEN_7329; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7331 = 8'ha3 == io_state_in_14 ? 8'h5d : _GEN_7330; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7332 = 8'ha4 == io_state_in_14 ? 8'h53 : _GEN_7331; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7333 = 8'ha5 == io_state_in_14 ? 8'h51 : _GEN_7332; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7334 = 8'ha6 == io_state_in_14 ? 8'h57 : _GEN_7333; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7335 = 8'ha7 == io_state_in_14 ? 8'h55 : _GEN_7334; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7336 = 8'ha8 == io_state_in_14 ? 8'h4b : _GEN_7335; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7337 = 8'ha9 == io_state_in_14 ? 8'h49 : _GEN_7336; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7338 = 8'haa == io_state_in_14 ? 8'h4f : _GEN_7337; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7339 = 8'hab == io_state_in_14 ? 8'h4d : _GEN_7338; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7340 = 8'hac == io_state_in_14 ? 8'h43 : _GEN_7339; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7341 = 8'had == io_state_in_14 ? 8'h41 : _GEN_7340; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7342 = 8'hae == io_state_in_14 ? 8'h47 : _GEN_7341; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7343 = 8'haf == io_state_in_14 ? 8'h45 : _GEN_7342; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7344 = 8'hb0 == io_state_in_14 ? 8'h7b : _GEN_7343; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7345 = 8'hb1 == io_state_in_14 ? 8'h79 : _GEN_7344; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7346 = 8'hb2 == io_state_in_14 ? 8'h7f : _GEN_7345; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7347 = 8'hb3 == io_state_in_14 ? 8'h7d : _GEN_7346; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7348 = 8'hb4 == io_state_in_14 ? 8'h73 : _GEN_7347; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7349 = 8'hb5 == io_state_in_14 ? 8'h71 : _GEN_7348; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7350 = 8'hb6 == io_state_in_14 ? 8'h77 : _GEN_7349; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7351 = 8'hb7 == io_state_in_14 ? 8'h75 : _GEN_7350; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7352 = 8'hb8 == io_state_in_14 ? 8'h6b : _GEN_7351; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7353 = 8'hb9 == io_state_in_14 ? 8'h69 : _GEN_7352; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7354 = 8'hba == io_state_in_14 ? 8'h6f : _GEN_7353; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7355 = 8'hbb == io_state_in_14 ? 8'h6d : _GEN_7354; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7356 = 8'hbc == io_state_in_14 ? 8'h63 : _GEN_7355; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7357 = 8'hbd == io_state_in_14 ? 8'h61 : _GEN_7356; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7358 = 8'hbe == io_state_in_14 ? 8'h67 : _GEN_7357; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7359 = 8'hbf == io_state_in_14 ? 8'h65 : _GEN_7358; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7360 = 8'hc0 == io_state_in_14 ? 8'h9b : _GEN_7359; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7361 = 8'hc1 == io_state_in_14 ? 8'h99 : _GEN_7360; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7362 = 8'hc2 == io_state_in_14 ? 8'h9f : _GEN_7361; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7363 = 8'hc3 == io_state_in_14 ? 8'h9d : _GEN_7362; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7364 = 8'hc4 == io_state_in_14 ? 8'h93 : _GEN_7363; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7365 = 8'hc5 == io_state_in_14 ? 8'h91 : _GEN_7364; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7366 = 8'hc6 == io_state_in_14 ? 8'h97 : _GEN_7365; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7367 = 8'hc7 == io_state_in_14 ? 8'h95 : _GEN_7366; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7368 = 8'hc8 == io_state_in_14 ? 8'h8b : _GEN_7367; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7369 = 8'hc9 == io_state_in_14 ? 8'h89 : _GEN_7368; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7370 = 8'hca == io_state_in_14 ? 8'h8f : _GEN_7369; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7371 = 8'hcb == io_state_in_14 ? 8'h8d : _GEN_7370; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7372 = 8'hcc == io_state_in_14 ? 8'h83 : _GEN_7371; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7373 = 8'hcd == io_state_in_14 ? 8'h81 : _GEN_7372; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7374 = 8'hce == io_state_in_14 ? 8'h87 : _GEN_7373; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7375 = 8'hcf == io_state_in_14 ? 8'h85 : _GEN_7374; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7376 = 8'hd0 == io_state_in_14 ? 8'hbb : _GEN_7375; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7377 = 8'hd1 == io_state_in_14 ? 8'hb9 : _GEN_7376; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7378 = 8'hd2 == io_state_in_14 ? 8'hbf : _GEN_7377; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7379 = 8'hd3 == io_state_in_14 ? 8'hbd : _GEN_7378; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7380 = 8'hd4 == io_state_in_14 ? 8'hb3 : _GEN_7379; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7381 = 8'hd5 == io_state_in_14 ? 8'hb1 : _GEN_7380; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7382 = 8'hd6 == io_state_in_14 ? 8'hb7 : _GEN_7381; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7383 = 8'hd7 == io_state_in_14 ? 8'hb5 : _GEN_7382; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7384 = 8'hd8 == io_state_in_14 ? 8'hab : _GEN_7383; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7385 = 8'hd9 == io_state_in_14 ? 8'ha9 : _GEN_7384; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7386 = 8'hda == io_state_in_14 ? 8'haf : _GEN_7385; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7387 = 8'hdb == io_state_in_14 ? 8'had : _GEN_7386; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7388 = 8'hdc == io_state_in_14 ? 8'ha3 : _GEN_7387; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7389 = 8'hdd == io_state_in_14 ? 8'ha1 : _GEN_7388; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7390 = 8'hde == io_state_in_14 ? 8'ha7 : _GEN_7389; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7391 = 8'hdf == io_state_in_14 ? 8'ha5 : _GEN_7390; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7392 = 8'he0 == io_state_in_14 ? 8'hdb : _GEN_7391; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7393 = 8'he1 == io_state_in_14 ? 8'hd9 : _GEN_7392; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7394 = 8'he2 == io_state_in_14 ? 8'hdf : _GEN_7393; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7395 = 8'he3 == io_state_in_14 ? 8'hdd : _GEN_7394; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7396 = 8'he4 == io_state_in_14 ? 8'hd3 : _GEN_7395; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7397 = 8'he5 == io_state_in_14 ? 8'hd1 : _GEN_7396; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7398 = 8'he6 == io_state_in_14 ? 8'hd7 : _GEN_7397; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7399 = 8'he7 == io_state_in_14 ? 8'hd5 : _GEN_7398; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7400 = 8'he8 == io_state_in_14 ? 8'hcb : _GEN_7399; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7401 = 8'he9 == io_state_in_14 ? 8'hc9 : _GEN_7400; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7402 = 8'hea == io_state_in_14 ? 8'hcf : _GEN_7401; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7403 = 8'heb == io_state_in_14 ? 8'hcd : _GEN_7402; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7404 = 8'hec == io_state_in_14 ? 8'hc3 : _GEN_7403; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7405 = 8'hed == io_state_in_14 ? 8'hc1 : _GEN_7404; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7406 = 8'hee == io_state_in_14 ? 8'hc7 : _GEN_7405; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7407 = 8'hef == io_state_in_14 ? 8'hc5 : _GEN_7406; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7408 = 8'hf0 == io_state_in_14 ? 8'hfb : _GEN_7407; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7409 = 8'hf1 == io_state_in_14 ? 8'hf9 : _GEN_7408; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7410 = 8'hf2 == io_state_in_14 ? 8'hff : _GEN_7409; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7411 = 8'hf3 == io_state_in_14 ? 8'hfd : _GEN_7410; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7412 = 8'hf4 == io_state_in_14 ? 8'hf3 : _GEN_7411; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7413 = 8'hf5 == io_state_in_14 ? 8'hf1 : _GEN_7412; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7414 = 8'hf6 == io_state_in_14 ? 8'hf7 : _GEN_7413; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7415 = 8'hf7 == io_state_in_14 ? 8'hf5 : _GEN_7414; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7416 = 8'hf8 == io_state_in_14 ? 8'heb : _GEN_7415; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7417 = 8'hf9 == io_state_in_14 ? 8'he9 : _GEN_7416; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7418 = 8'hfa == io_state_in_14 ? 8'hef : _GEN_7417; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7419 = 8'hfb == io_state_in_14 ? 8'hed : _GEN_7418; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7420 = 8'hfc == io_state_in_14 ? 8'he3 : _GEN_7419; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7421 = 8'hfd == io_state_in_14 ? 8'he1 : _GEN_7420; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7422 = 8'hfe == io_state_in_14 ? 8'he7 : _GEN_7421; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _GEN_7423 = 8'hff == io_state_in_14 ? 8'he5 : _GEN_7422; // @[MixColumns.scala 142:{54,54}]
  wire [7:0] _tmp_state_14_T_1 = _tmp_state_14_T ^ _GEN_7423; // @[MixColumns.scala 142:54]
  wire [7:0] _GEN_7425 = 8'h1 == io_state_in_15 ? 8'h3 : 8'h0; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7426 = 8'h2 == io_state_in_15 ? 8'h6 : _GEN_7425; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7427 = 8'h3 == io_state_in_15 ? 8'h5 : _GEN_7426; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7428 = 8'h4 == io_state_in_15 ? 8'hc : _GEN_7427; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7429 = 8'h5 == io_state_in_15 ? 8'hf : _GEN_7428; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7430 = 8'h6 == io_state_in_15 ? 8'ha : _GEN_7429; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7431 = 8'h7 == io_state_in_15 ? 8'h9 : _GEN_7430; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7432 = 8'h8 == io_state_in_15 ? 8'h18 : _GEN_7431; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7433 = 8'h9 == io_state_in_15 ? 8'h1b : _GEN_7432; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7434 = 8'ha == io_state_in_15 ? 8'h1e : _GEN_7433; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7435 = 8'hb == io_state_in_15 ? 8'h1d : _GEN_7434; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7436 = 8'hc == io_state_in_15 ? 8'h14 : _GEN_7435; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7437 = 8'hd == io_state_in_15 ? 8'h17 : _GEN_7436; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7438 = 8'he == io_state_in_15 ? 8'h12 : _GEN_7437; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7439 = 8'hf == io_state_in_15 ? 8'h11 : _GEN_7438; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7440 = 8'h10 == io_state_in_15 ? 8'h30 : _GEN_7439; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7441 = 8'h11 == io_state_in_15 ? 8'h33 : _GEN_7440; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7442 = 8'h12 == io_state_in_15 ? 8'h36 : _GEN_7441; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7443 = 8'h13 == io_state_in_15 ? 8'h35 : _GEN_7442; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7444 = 8'h14 == io_state_in_15 ? 8'h3c : _GEN_7443; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7445 = 8'h15 == io_state_in_15 ? 8'h3f : _GEN_7444; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7446 = 8'h16 == io_state_in_15 ? 8'h3a : _GEN_7445; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7447 = 8'h17 == io_state_in_15 ? 8'h39 : _GEN_7446; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7448 = 8'h18 == io_state_in_15 ? 8'h28 : _GEN_7447; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7449 = 8'h19 == io_state_in_15 ? 8'h2b : _GEN_7448; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7450 = 8'h1a == io_state_in_15 ? 8'h2e : _GEN_7449; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7451 = 8'h1b == io_state_in_15 ? 8'h2d : _GEN_7450; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7452 = 8'h1c == io_state_in_15 ? 8'h24 : _GEN_7451; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7453 = 8'h1d == io_state_in_15 ? 8'h27 : _GEN_7452; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7454 = 8'h1e == io_state_in_15 ? 8'h22 : _GEN_7453; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7455 = 8'h1f == io_state_in_15 ? 8'h21 : _GEN_7454; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7456 = 8'h20 == io_state_in_15 ? 8'h60 : _GEN_7455; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7457 = 8'h21 == io_state_in_15 ? 8'h63 : _GEN_7456; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7458 = 8'h22 == io_state_in_15 ? 8'h66 : _GEN_7457; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7459 = 8'h23 == io_state_in_15 ? 8'h65 : _GEN_7458; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7460 = 8'h24 == io_state_in_15 ? 8'h6c : _GEN_7459; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7461 = 8'h25 == io_state_in_15 ? 8'h6f : _GEN_7460; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7462 = 8'h26 == io_state_in_15 ? 8'h6a : _GEN_7461; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7463 = 8'h27 == io_state_in_15 ? 8'h69 : _GEN_7462; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7464 = 8'h28 == io_state_in_15 ? 8'h78 : _GEN_7463; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7465 = 8'h29 == io_state_in_15 ? 8'h7b : _GEN_7464; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7466 = 8'h2a == io_state_in_15 ? 8'h7e : _GEN_7465; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7467 = 8'h2b == io_state_in_15 ? 8'h7d : _GEN_7466; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7468 = 8'h2c == io_state_in_15 ? 8'h74 : _GEN_7467; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7469 = 8'h2d == io_state_in_15 ? 8'h77 : _GEN_7468; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7470 = 8'h2e == io_state_in_15 ? 8'h72 : _GEN_7469; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7471 = 8'h2f == io_state_in_15 ? 8'h71 : _GEN_7470; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7472 = 8'h30 == io_state_in_15 ? 8'h50 : _GEN_7471; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7473 = 8'h31 == io_state_in_15 ? 8'h53 : _GEN_7472; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7474 = 8'h32 == io_state_in_15 ? 8'h56 : _GEN_7473; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7475 = 8'h33 == io_state_in_15 ? 8'h55 : _GEN_7474; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7476 = 8'h34 == io_state_in_15 ? 8'h5c : _GEN_7475; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7477 = 8'h35 == io_state_in_15 ? 8'h5f : _GEN_7476; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7478 = 8'h36 == io_state_in_15 ? 8'h5a : _GEN_7477; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7479 = 8'h37 == io_state_in_15 ? 8'h59 : _GEN_7478; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7480 = 8'h38 == io_state_in_15 ? 8'h48 : _GEN_7479; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7481 = 8'h39 == io_state_in_15 ? 8'h4b : _GEN_7480; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7482 = 8'h3a == io_state_in_15 ? 8'h4e : _GEN_7481; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7483 = 8'h3b == io_state_in_15 ? 8'h4d : _GEN_7482; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7484 = 8'h3c == io_state_in_15 ? 8'h44 : _GEN_7483; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7485 = 8'h3d == io_state_in_15 ? 8'h47 : _GEN_7484; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7486 = 8'h3e == io_state_in_15 ? 8'h42 : _GEN_7485; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7487 = 8'h3f == io_state_in_15 ? 8'h41 : _GEN_7486; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7488 = 8'h40 == io_state_in_15 ? 8'hc0 : _GEN_7487; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7489 = 8'h41 == io_state_in_15 ? 8'hc3 : _GEN_7488; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7490 = 8'h42 == io_state_in_15 ? 8'hc6 : _GEN_7489; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7491 = 8'h43 == io_state_in_15 ? 8'hc5 : _GEN_7490; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7492 = 8'h44 == io_state_in_15 ? 8'hcc : _GEN_7491; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7493 = 8'h45 == io_state_in_15 ? 8'hcf : _GEN_7492; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7494 = 8'h46 == io_state_in_15 ? 8'hca : _GEN_7493; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7495 = 8'h47 == io_state_in_15 ? 8'hc9 : _GEN_7494; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7496 = 8'h48 == io_state_in_15 ? 8'hd8 : _GEN_7495; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7497 = 8'h49 == io_state_in_15 ? 8'hdb : _GEN_7496; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7498 = 8'h4a == io_state_in_15 ? 8'hde : _GEN_7497; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7499 = 8'h4b == io_state_in_15 ? 8'hdd : _GEN_7498; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7500 = 8'h4c == io_state_in_15 ? 8'hd4 : _GEN_7499; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7501 = 8'h4d == io_state_in_15 ? 8'hd7 : _GEN_7500; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7502 = 8'h4e == io_state_in_15 ? 8'hd2 : _GEN_7501; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7503 = 8'h4f == io_state_in_15 ? 8'hd1 : _GEN_7502; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7504 = 8'h50 == io_state_in_15 ? 8'hf0 : _GEN_7503; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7505 = 8'h51 == io_state_in_15 ? 8'hf3 : _GEN_7504; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7506 = 8'h52 == io_state_in_15 ? 8'hf6 : _GEN_7505; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7507 = 8'h53 == io_state_in_15 ? 8'hf5 : _GEN_7506; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7508 = 8'h54 == io_state_in_15 ? 8'hfc : _GEN_7507; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7509 = 8'h55 == io_state_in_15 ? 8'hff : _GEN_7508; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7510 = 8'h56 == io_state_in_15 ? 8'hfa : _GEN_7509; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7511 = 8'h57 == io_state_in_15 ? 8'hf9 : _GEN_7510; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7512 = 8'h58 == io_state_in_15 ? 8'he8 : _GEN_7511; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7513 = 8'h59 == io_state_in_15 ? 8'heb : _GEN_7512; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7514 = 8'h5a == io_state_in_15 ? 8'hee : _GEN_7513; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7515 = 8'h5b == io_state_in_15 ? 8'hed : _GEN_7514; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7516 = 8'h5c == io_state_in_15 ? 8'he4 : _GEN_7515; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7517 = 8'h5d == io_state_in_15 ? 8'he7 : _GEN_7516; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7518 = 8'h5e == io_state_in_15 ? 8'he2 : _GEN_7517; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7519 = 8'h5f == io_state_in_15 ? 8'he1 : _GEN_7518; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7520 = 8'h60 == io_state_in_15 ? 8'ha0 : _GEN_7519; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7521 = 8'h61 == io_state_in_15 ? 8'ha3 : _GEN_7520; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7522 = 8'h62 == io_state_in_15 ? 8'ha6 : _GEN_7521; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7523 = 8'h63 == io_state_in_15 ? 8'ha5 : _GEN_7522; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7524 = 8'h64 == io_state_in_15 ? 8'hac : _GEN_7523; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7525 = 8'h65 == io_state_in_15 ? 8'haf : _GEN_7524; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7526 = 8'h66 == io_state_in_15 ? 8'haa : _GEN_7525; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7527 = 8'h67 == io_state_in_15 ? 8'ha9 : _GEN_7526; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7528 = 8'h68 == io_state_in_15 ? 8'hb8 : _GEN_7527; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7529 = 8'h69 == io_state_in_15 ? 8'hbb : _GEN_7528; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7530 = 8'h6a == io_state_in_15 ? 8'hbe : _GEN_7529; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7531 = 8'h6b == io_state_in_15 ? 8'hbd : _GEN_7530; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7532 = 8'h6c == io_state_in_15 ? 8'hb4 : _GEN_7531; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7533 = 8'h6d == io_state_in_15 ? 8'hb7 : _GEN_7532; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7534 = 8'h6e == io_state_in_15 ? 8'hb2 : _GEN_7533; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7535 = 8'h6f == io_state_in_15 ? 8'hb1 : _GEN_7534; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7536 = 8'h70 == io_state_in_15 ? 8'h90 : _GEN_7535; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7537 = 8'h71 == io_state_in_15 ? 8'h93 : _GEN_7536; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7538 = 8'h72 == io_state_in_15 ? 8'h96 : _GEN_7537; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7539 = 8'h73 == io_state_in_15 ? 8'h95 : _GEN_7538; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7540 = 8'h74 == io_state_in_15 ? 8'h9c : _GEN_7539; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7541 = 8'h75 == io_state_in_15 ? 8'h9f : _GEN_7540; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7542 = 8'h76 == io_state_in_15 ? 8'h9a : _GEN_7541; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7543 = 8'h77 == io_state_in_15 ? 8'h99 : _GEN_7542; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7544 = 8'h78 == io_state_in_15 ? 8'h88 : _GEN_7543; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7545 = 8'h79 == io_state_in_15 ? 8'h8b : _GEN_7544; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7546 = 8'h7a == io_state_in_15 ? 8'h8e : _GEN_7545; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7547 = 8'h7b == io_state_in_15 ? 8'h8d : _GEN_7546; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7548 = 8'h7c == io_state_in_15 ? 8'h84 : _GEN_7547; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7549 = 8'h7d == io_state_in_15 ? 8'h87 : _GEN_7548; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7550 = 8'h7e == io_state_in_15 ? 8'h82 : _GEN_7549; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7551 = 8'h7f == io_state_in_15 ? 8'h81 : _GEN_7550; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7552 = 8'h80 == io_state_in_15 ? 8'h9b : _GEN_7551; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7553 = 8'h81 == io_state_in_15 ? 8'h98 : _GEN_7552; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7554 = 8'h82 == io_state_in_15 ? 8'h9d : _GEN_7553; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7555 = 8'h83 == io_state_in_15 ? 8'h9e : _GEN_7554; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7556 = 8'h84 == io_state_in_15 ? 8'h97 : _GEN_7555; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7557 = 8'h85 == io_state_in_15 ? 8'h94 : _GEN_7556; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7558 = 8'h86 == io_state_in_15 ? 8'h91 : _GEN_7557; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7559 = 8'h87 == io_state_in_15 ? 8'h92 : _GEN_7558; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7560 = 8'h88 == io_state_in_15 ? 8'h83 : _GEN_7559; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7561 = 8'h89 == io_state_in_15 ? 8'h80 : _GEN_7560; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7562 = 8'h8a == io_state_in_15 ? 8'h85 : _GEN_7561; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7563 = 8'h8b == io_state_in_15 ? 8'h86 : _GEN_7562; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7564 = 8'h8c == io_state_in_15 ? 8'h8f : _GEN_7563; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7565 = 8'h8d == io_state_in_15 ? 8'h8c : _GEN_7564; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7566 = 8'h8e == io_state_in_15 ? 8'h89 : _GEN_7565; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7567 = 8'h8f == io_state_in_15 ? 8'h8a : _GEN_7566; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7568 = 8'h90 == io_state_in_15 ? 8'hab : _GEN_7567; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7569 = 8'h91 == io_state_in_15 ? 8'ha8 : _GEN_7568; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7570 = 8'h92 == io_state_in_15 ? 8'had : _GEN_7569; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7571 = 8'h93 == io_state_in_15 ? 8'hae : _GEN_7570; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7572 = 8'h94 == io_state_in_15 ? 8'ha7 : _GEN_7571; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7573 = 8'h95 == io_state_in_15 ? 8'ha4 : _GEN_7572; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7574 = 8'h96 == io_state_in_15 ? 8'ha1 : _GEN_7573; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7575 = 8'h97 == io_state_in_15 ? 8'ha2 : _GEN_7574; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7576 = 8'h98 == io_state_in_15 ? 8'hb3 : _GEN_7575; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7577 = 8'h99 == io_state_in_15 ? 8'hb0 : _GEN_7576; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7578 = 8'h9a == io_state_in_15 ? 8'hb5 : _GEN_7577; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7579 = 8'h9b == io_state_in_15 ? 8'hb6 : _GEN_7578; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7580 = 8'h9c == io_state_in_15 ? 8'hbf : _GEN_7579; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7581 = 8'h9d == io_state_in_15 ? 8'hbc : _GEN_7580; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7582 = 8'h9e == io_state_in_15 ? 8'hb9 : _GEN_7581; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7583 = 8'h9f == io_state_in_15 ? 8'hba : _GEN_7582; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7584 = 8'ha0 == io_state_in_15 ? 8'hfb : _GEN_7583; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7585 = 8'ha1 == io_state_in_15 ? 8'hf8 : _GEN_7584; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7586 = 8'ha2 == io_state_in_15 ? 8'hfd : _GEN_7585; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7587 = 8'ha3 == io_state_in_15 ? 8'hfe : _GEN_7586; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7588 = 8'ha4 == io_state_in_15 ? 8'hf7 : _GEN_7587; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7589 = 8'ha5 == io_state_in_15 ? 8'hf4 : _GEN_7588; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7590 = 8'ha6 == io_state_in_15 ? 8'hf1 : _GEN_7589; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7591 = 8'ha7 == io_state_in_15 ? 8'hf2 : _GEN_7590; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7592 = 8'ha8 == io_state_in_15 ? 8'he3 : _GEN_7591; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7593 = 8'ha9 == io_state_in_15 ? 8'he0 : _GEN_7592; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7594 = 8'haa == io_state_in_15 ? 8'he5 : _GEN_7593; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7595 = 8'hab == io_state_in_15 ? 8'he6 : _GEN_7594; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7596 = 8'hac == io_state_in_15 ? 8'hef : _GEN_7595; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7597 = 8'had == io_state_in_15 ? 8'hec : _GEN_7596; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7598 = 8'hae == io_state_in_15 ? 8'he9 : _GEN_7597; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7599 = 8'haf == io_state_in_15 ? 8'hea : _GEN_7598; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7600 = 8'hb0 == io_state_in_15 ? 8'hcb : _GEN_7599; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7601 = 8'hb1 == io_state_in_15 ? 8'hc8 : _GEN_7600; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7602 = 8'hb2 == io_state_in_15 ? 8'hcd : _GEN_7601; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7603 = 8'hb3 == io_state_in_15 ? 8'hce : _GEN_7602; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7604 = 8'hb4 == io_state_in_15 ? 8'hc7 : _GEN_7603; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7605 = 8'hb5 == io_state_in_15 ? 8'hc4 : _GEN_7604; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7606 = 8'hb6 == io_state_in_15 ? 8'hc1 : _GEN_7605; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7607 = 8'hb7 == io_state_in_15 ? 8'hc2 : _GEN_7606; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7608 = 8'hb8 == io_state_in_15 ? 8'hd3 : _GEN_7607; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7609 = 8'hb9 == io_state_in_15 ? 8'hd0 : _GEN_7608; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7610 = 8'hba == io_state_in_15 ? 8'hd5 : _GEN_7609; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7611 = 8'hbb == io_state_in_15 ? 8'hd6 : _GEN_7610; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7612 = 8'hbc == io_state_in_15 ? 8'hdf : _GEN_7611; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7613 = 8'hbd == io_state_in_15 ? 8'hdc : _GEN_7612; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7614 = 8'hbe == io_state_in_15 ? 8'hd9 : _GEN_7613; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7615 = 8'hbf == io_state_in_15 ? 8'hda : _GEN_7614; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7616 = 8'hc0 == io_state_in_15 ? 8'h5b : _GEN_7615; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7617 = 8'hc1 == io_state_in_15 ? 8'h58 : _GEN_7616; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7618 = 8'hc2 == io_state_in_15 ? 8'h5d : _GEN_7617; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7619 = 8'hc3 == io_state_in_15 ? 8'h5e : _GEN_7618; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7620 = 8'hc4 == io_state_in_15 ? 8'h57 : _GEN_7619; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7621 = 8'hc5 == io_state_in_15 ? 8'h54 : _GEN_7620; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7622 = 8'hc6 == io_state_in_15 ? 8'h51 : _GEN_7621; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7623 = 8'hc7 == io_state_in_15 ? 8'h52 : _GEN_7622; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7624 = 8'hc8 == io_state_in_15 ? 8'h43 : _GEN_7623; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7625 = 8'hc9 == io_state_in_15 ? 8'h40 : _GEN_7624; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7626 = 8'hca == io_state_in_15 ? 8'h45 : _GEN_7625; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7627 = 8'hcb == io_state_in_15 ? 8'h46 : _GEN_7626; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7628 = 8'hcc == io_state_in_15 ? 8'h4f : _GEN_7627; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7629 = 8'hcd == io_state_in_15 ? 8'h4c : _GEN_7628; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7630 = 8'hce == io_state_in_15 ? 8'h49 : _GEN_7629; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7631 = 8'hcf == io_state_in_15 ? 8'h4a : _GEN_7630; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7632 = 8'hd0 == io_state_in_15 ? 8'h6b : _GEN_7631; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7633 = 8'hd1 == io_state_in_15 ? 8'h68 : _GEN_7632; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7634 = 8'hd2 == io_state_in_15 ? 8'h6d : _GEN_7633; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7635 = 8'hd3 == io_state_in_15 ? 8'h6e : _GEN_7634; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7636 = 8'hd4 == io_state_in_15 ? 8'h67 : _GEN_7635; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7637 = 8'hd5 == io_state_in_15 ? 8'h64 : _GEN_7636; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7638 = 8'hd6 == io_state_in_15 ? 8'h61 : _GEN_7637; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7639 = 8'hd7 == io_state_in_15 ? 8'h62 : _GEN_7638; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7640 = 8'hd8 == io_state_in_15 ? 8'h73 : _GEN_7639; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7641 = 8'hd9 == io_state_in_15 ? 8'h70 : _GEN_7640; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7642 = 8'hda == io_state_in_15 ? 8'h75 : _GEN_7641; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7643 = 8'hdb == io_state_in_15 ? 8'h76 : _GEN_7642; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7644 = 8'hdc == io_state_in_15 ? 8'h7f : _GEN_7643; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7645 = 8'hdd == io_state_in_15 ? 8'h7c : _GEN_7644; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7646 = 8'hde == io_state_in_15 ? 8'h79 : _GEN_7645; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7647 = 8'hdf == io_state_in_15 ? 8'h7a : _GEN_7646; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7648 = 8'he0 == io_state_in_15 ? 8'h3b : _GEN_7647; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7649 = 8'he1 == io_state_in_15 ? 8'h38 : _GEN_7648; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7650 = 8'he2 == io_state_in_15 ? 8'h3d : _GEN_7649; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7651 = 8'he3 == io_state_in_15 ? 8'h3e : _GEN_7650; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7652 = 8'he4 == io_state_in_15 ? 8'h37 : _GEN_7651; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7653 = 8'he5 == io_state_in_15 ? 8'h34 : _GEN_7652; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7654 = 8'he6 == io_state_in_15 ? 8'h31 : _GEN_7653; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7655 = 8'he7 == io_state_in_15 ? 8'h32 : _GEN_7654; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7656 = 8'he8 == io_state_in_15 ? 8'h23 : _GEN_7655; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7657 = 8'he9 == io_state_in_15 ? 8'h20 : _GEN_7656; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7658 = 8'hea == io_state_in_15 ? 8'h25 : _GEN_7657; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7659 = 8'heb == io_state_in_15 ? 8'h26 : _GEN_7658; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7660 = 8'hec == io_state_in_15 ? 8'h2f : _GEN_7659; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7661 = 8'hed == io_state_in_15 ? 8'h2c : _GEN_7660; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7662 = 8'hee == io_state_in_15 ? 8'h29 : _GEN_7661; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7663 = 8'hef == io_state_in_15 ? 8'h2a : _GEN_7662; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7664 = 8'hf0 == io_state_in_15 ? 8'hb : _GEN_7663; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7665 = 8'hf1 == io_state_in_15 ? 8'h8 : _GEN_7664; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7666 = 8'hf2 == io_state_in_15 ? 8'hd : _GEN_7665; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7667 = 8'hf3 == io_state_in_15 ? 8'he : _GEN_7666; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7668 = 8'hf4 == io_state_in_15 ? 8'h7 : _GEN_7667; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7669 = 8'hf5 == io_state_in_15 ? 8'h4 : _GEN_7668; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7670 = 8'hf6 == io_state_in_15 ? 8'h1 : _GEN_7669; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7671 = 8'hf7 == io_state_in_15 ? 8'h2 : _GEN_7670; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7672 = 8'hf8 == io_state_in_15 ? 8'h13 : _GEN_7671; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7673 = 8'hf9 == io_state_in_15 ? 8'h10 : _GEN_7672; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7674 = 8'hfa == io_state_in_15 ? 8'h15 : _GEN_7673; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7675 = 8'hfb == io_state_in_15 ? 8'h16 : _GEN_7674; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7676 = 8'hfc == io_state_in_15 ? 8'h1f : _GEN_7675; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7677 = 8'hfd == io_state_in_15 ? 8'h1c : _GEN_7676; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7678 = 8'hfe == io_state_in_15 ? 8'h19 : _GEN_7677; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7679 = 8'hff == io_state_in_15 ? 8'h1a : _GEN_7678; // @[MixColumns.scala 142:{79,79}]
  wire [7:0] _GEN_7681 = 8'h1 == io_state_in_12 ? 8'h3 : 8'h0; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7682 = 8'h2 == io_state_in_12 ? 8'h6 : _GEN_7681; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7683 = 8'h3 == io_state_in_12 ? 8'h5 : _GEN_7682; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7684 = 8'h4 == io_state_in_12 ? 8'hc : _GEN_7683; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7685 = 8'h5 == io_state_in_12 ? 8'hf : _GEN_7684; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7686 = 8'h6 == io_state_in_12 ? 8'ha : _GEN_7685; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7687 = 8'h7 == io_state_in_12 ? 8'h9 : _GEN_7686; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7688 = 8'h8 == io_state_in_12 ? 8'h18 : _GEN_7687; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7689 = 8'h9 == io_state_in_12 ? 8'h1b : _GEN_7688; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7690 = 8'ha == io_state_in_12 ? 8'h1e : _GEN_7689; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7691 = 8'hb == io_state_in_12 ? 8'h1d : _GEN_7690; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7692 = 8'hc == io_state_in_12 ? 8'h14 : _GEN_7691; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7693 = 8'hd == io_state_in_12 ? 8'h17 : _GEN_7692; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7694 = 8'he == io_state_in_12 ? 8'h12 : _GEN_7693; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7695 = 8'hf == io_state_in_12 ? 8'h11 : _GEN_7694; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7696 = 8'h10 == io_state_in_12 ? 8'h30 : _GEN_7695; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7697 = 8'h11 == io_state_in_12 ? 8'h33 : _GEN_7696; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7698 = 8'h12 == io_state_in_12 ? 8'h36 : _GEN_7697; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7699 = 8'h13 == io_state_in_12 ? 8'h35 : _GEN_7698; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7700 = 8'h14 == io_state_in_12 ? 8'h3c : _GEN_7699; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7701 = 8'h15 == io_state_in_12 ? 8'h3f : _GEN_7700; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7702 = 8'h16 == io_state_in_12 ? 8'h3a : _GEN_7701; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7703 = 8'h17 == io_state_in_12 ? 8'h39 : _GEN_7702; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7704 = 8'h18 == io_state_in_12 ? 8'h28 : _GEN_7703; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7705 = 8'h19 == io_state_in_12 ? 8'h2b : _GEN_7704; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7706 = 8'h1a == io_state_in_12 ? 8'h2e : _GEN_7705; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7707 = 8'h1b == io_state_in_12 ? 8'h2d : _GEN_7706; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7708 = 8'h1c == io_state_in_12 ? 8'h24 : _GEN_7707; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7709 = 8'h1d == io_state_in_12 ? 8'h27 : _GEN_7708; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7710 = 8'h1e == io_state_in_12 ? 8'h22 : _GEN_7709; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7711 = 8'h1f == io_state_in_12 ? 8'h21 : _GEN_7710; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7712 = 8'h20 == io_state_in_12 ? 8'h60 : _GEN_7711; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7713 = 8'h21 == io_state_in_12 ? 8'h63 : _GEN_7712; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7714 = 8'h22 == io_state_in_12 ? 8'h66 : _GEN_7713; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7715 = 8'h23 == io_state_in_12 ? 8'h65 : _GEN_7714; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7716 = 8'h24 == io_state_in_12 ? 8'h6c : _GEN_7715; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7717 = 8'h25 == io_state_in_12 ? 8'h6f : _GEN_7716; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7718 = 8'h26 == io_state_in_12 ? 8'h6a : _GEN_7717; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7719 = 8'h27 == io_state_in_12 ? 8'h69 : _GEN_7718; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7720 = 8'h28 == io_state_in_12 ? 8'h78 : _GEN_7719; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7721 = 8'h29 == io_state_in_12 ? 8'h7b : _GEN_7720; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7722 = 8'h2a == io_state_in_12 ? 8'h7e : _GEN_7721; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7723 = 8'h2b == io_state_in_12 ? 8'h7d : _GEN_7722; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7724 = 8'h2c == io_state_in_12 ? 8'h74 : _GEN_7723; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7725 = 8'h2d == io_state_in_12 ? 8'h77 : _GEN_7724; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7726 = 8'h2e == io_state_in_12 ? 8'h72 : _GEN_7725; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7727 = 8'h2f == io_state_in_12 ? 8'h71 : _GEN_7726; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7728 = 8'h30 == io_state_in_12 ? 8'h50 : _GEN_7727; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7729 = 8'h31 == io_state_in_12 ? 8'h53 : _GEN_7728; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7730 = 8'h32 == io_state_in_12 ? 8'h56 : _GEN_7729; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7731 = 8'h33 == io_state_in_12 ? 8'h55 : _GEN_7730; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7732 = 8'h34 == io_state_in_12 ? 8'h5c : _GEN_7731; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7733 = 8'h35 == io_state_in_12 ? 8'h5f : _GEN_7732; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7734 = 8'h36 == io_state_in_12 ? 8'h5a : _GEN_7733; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7735 = 8'h37 == io_state_in_12 ? 8'h59 : _GEN_7734; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7736 = 8'h38 == io_state_in_12 ? 8'h48 : _GEN_7735; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7737 = 8'h39 == io_state_in_12 ? 8'h4b : _GEN_7736; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7738 = 8'h3a == io_state_in_12 ? 8'h4e : _GEN_7737; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7739 = 8'h3b == io_state_in_12 ? 8'h4d : _GEN_7738; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7740 = 8'h3c == io_state_in_12 ? 8'h44 : _GEN_7739; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7741 = 8'h3d == io_state_in_12 ? 8'h47 : _GEN_7740; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7742 = 8'h3e == io_state_in_12 ? 8'h42 : _GEN_7741; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7743 = 8'h3f == io_state_in_12 ? 8'h41 : _GEN_7742; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7744 = 8'h40 == io_state_in_12 ? 8'hc0 : _GEN_7743; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7745 = 8'h41 == io_state_in_12 ? 8'hc3 : _GEN_7744; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7746 = 8'h42 == io_state_in_12 ? 8'hc6 : _GEN_7745; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7747 = 8'h43 == io_state_in_12 ? 8'hc5 : _GEN_7746; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7748 = 8'h44 == io_state_in_12 ? 8'hcc : _GEN_7747; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7749 = 8'h45 == io_state_in_12 ? 8'hcf : _GEN_7748; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7750 = 8'h46 == io_state_in_12 ? 8'hca : _GEN_7749; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7751 = 8'h47 == io_state_in_12 ? 8'hc9 : _GEN_7750; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7752 = 8'h48 == io_state_in_12 ? 8'hd8 : _GEN_7751; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7753 = 8'h49 == io_state_in_12 ? 8'hdb : _GEN_7752; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7754 = 8'h4a == io_state_in_12 ? 8'hde : _GEN_7753; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7755 = 8'h4b == io_state_in_12 ? 8'hdd : _GEN_7754; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7756 = 8'h4c == io_state_in_12 ? 8'hd4 : _GEN_7755; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7757 = 8'h4d == io_state_in_12 ? 8'hd7 : _GEN_7756; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7758 = 8'h4e == io_state_in_12 ? 8'hd2 : _GEN_7757; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7759 = 8'h4f == io_state_in_12 ? 8'hd1 : _GEN_7758; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7760 = 8'h50 == io_state_in_12 ? 8'hf0 : _GEN_7759; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7761 = 8'h51 == io_state_in_12 ? 8'hf3 : _GEN_7760; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7762 = 8'h52 == io_state_in_12 ? 8'hf6 : _GEN_7761; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7763 = 8'h53 == io_state_in_12 ? 8'hf5 : _GEN_7762; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7764 = 8'h54 == io_state_in_12 ? 8'hfc : _GEN_7763; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7765 = 8'h55 == io_state_in_12 ? 8'hff : _GEN_7764; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7766 = 8'h56 == io_state_in_12 ? 8'hfa : _GEN_7765; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7767 = 8'h57 == io_state_in_12 ? 8'hf9 : _GEN_7766; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7768 = 8'h58 == io_state_in_12 ? 8'he8 : _GEN_7767; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7769 = 8'h59 == io_state_in_12 ? 8'heb : _GEN_7768; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7770 = 8'h5a == io_state_in_12 ? 8'hee : _GEN_7769; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7771 = 8'h5b == io_state_in_12 ? 8'hed : _GEN_7770; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7772 = 8'h5c == io_state_in_12 ? 8'he4 : _GEN_7771; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7773 = 8'h5d == io_state_in_12 ? 8'he7 : _GEN_7772; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7774 = 8'h5e == io_state_in_12 ? 8'he2 : _GEN_7773; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7775 = 8'h5f == io_state_in_12 ? 8'he1 : _GEN_7774; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7776 = 8'h60 == io_state_in_12 ? 8'ha0 : _GEN_7775; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7777 = 8'h61 == io_state_in_12 ? 8'ha3 : _GEN_7776; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7778 = 8'h62 == io_state_in_12 ? 8'ha6 : _GEN_7777; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7779 = 8'h63 == io_state_in_12 ? 8'ha5 : _GEN_7778; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7780 = 8'h64 == io_state_in_12 ? 8'hac : _GEN_7779; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7781 = 8'h65 == io_state_in_12 ? 8'haf : _GEN_7780; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7782 = 8'h66 == io_state_in_12 ? 8'haa : _GEN_7781; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7783 = 8'h67 == io_state_in_12 ? 8'ha9 : _GEN_7782; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7784 = 8'h68 == io_state_in_12 ? 8'hb8 : _GEN_7783; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7785 = 8'h69 == io_state_in_12 ? 8'hbb : _GEN_7784; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7786 = 8'h6a == io_state_in_12 ? 8'hbe : _GEN_7785; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7787 = 8'h6b == io_state_in_12 ? 8'hbd : _GEN_7786; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7788 = 8'h6c == io_state_in_12 ? 8'hb4 : _GEN_7787; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7789 = 8'h6d == io_state_in_12 ? 8'hb7 : _GEN_7788; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7790 = 8'h6e == io_state_in_12 ? 8'hb2 : _GEN_7789; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7791 = 8'h6f == io_state_in_12 ? 8'hb1 : _GEN_7790; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7792 = 8'h70 == io_state_in_12 ? 8'h90 : _GEN_7791; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7793 = 8'h71 == io_state_in_12 ? 8'h93 : _GEN_7792; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7794 = 8'h72 == io_state_in_12 ? 8'h96 : _GEN_7793; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7795 = 8'h73 == io_state_in_12 ? 8'h95 : _GEN_7794; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7796 = 8'h74 == io_state_in_12 ? 8'h9c : _GEN_7795; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7797 = 8'h75 == io_state_in_12 ? 8'h9f : _GEN_7796; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7798 = 8'h76 == io_state_in_12 ? 8'h9a : _GEN_7797; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7799 = 8'h77 == io_state_in_12 ? 8'h99 : _GEN_7798; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7800 = 8'h78 == io_state_in_12 ? 8'h88 : _GEN_7799; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7801 = 8'h79 == io_state_in_12 ? 8'h8b : _GEN_7800; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7802 = 8'h7a == io_state_in_12 ? 8'h8e : _GEN_7801; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7803 = 8'h7b == io_state_in_12 ? 8'h8d : _GEN_7802; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7804 = 8'h7c == io_state_in_12 ? 8'h84 : _GEN_7803; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7805 = 8'h7d == io_state_in_12 ? 8'h87 : _GEN_7804; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7806 = 8'h7e == io_state_in_12 ? 8'h82 : _GEN_7805; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7807 = 8'h7f == io_state_in_12 ? 8'h81 : _GEN_7806; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7808 = 8'h80 == io_state_in_12 ? 8'h9b : _GEN_7807; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7809 = 8'h81 == io_state_in_12 ? 8'h98 : _GEN_7808; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7810 = 8'h82 == io_state_in_12 ? 8'h9d : _GEN_7809; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7811 = 8'h83 == io_state_in_12 ? 8'h9e : _GEN_7810; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7812 = 8'h84 == io_state_in_12 ? 8'h97 : _GEN_7811; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7813 = 8'h85 == io_state_in_12 ? 8'h94 : _GEN_7812; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7814 = 8'h86 == io_state_in_12 ? 8'h91 : _GEN_7813; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7815 = 8'h87 == io_state_in_12 ? 8'h92 : _GEN_7814; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7816 = 8'h88 == io_state_in_12 ? 8'h83 : _GEN_7815; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7817 = 8'h89 == io_state_in_12 ? 8'h80 : _GEN_7816; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7818 = 8'h8a == io_state_in_12 ? 8'h85 : _GEN_7817; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7819 = 8'h8b == io_state_in_12 ? 8'h86 : _GEN_7818; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7820 = 8'h8c == io_state_in_12 ? 8'h8f : _GEN_7819; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7821 = 8'h8d == io_state_in_12 ? 8'h8c : _GEN_7820; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7822 = 8'h8e == io_state_in_12 ? 8'h89 : _GEN_7821; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7823 = 8'h8f == io_state_in_12 ? 8'h8a : _GEN_7822; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7824 = 8'h90 == io_state_in_12 ? 8'hab : _GEN_7823; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7825 = 8'h91 == io_state_in_12 ? 8'ha8 : _GEN_7824; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7826 = 8'h92 == io_state_in_12 ? 8'had : _GEN_7825; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7827 = 8'h93 == io_state_in_12 ? 8'hae : _GEN_7826; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7828 = 8'h94 == io_state_in_12 ? 8'ha7 : _GEN_7827; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7829 = 8'h95 == io_state_in_12 ? 8'ha4 : _GEN_7828; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7830 = 8'h96 == io_state_in_12 ? 8'ha1 : _GEN_7829; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7831 = 8'h97 == io_state_in_12 ? 8'ha2 : _GEN_7830; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7832 = 8'h98 == io_state_in_12 ? 8'hb3 : _GEN_7831; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7833 = 8'h99 == io_state_in_12 ? 8'hb0 : _GEN_7832; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7834 = 8'h9a == io_state_in_12 ? 8'hb5 : _GEN_7833; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7835 = 8'h9b == io_state_in_12 ? 8'hb6 : _GEN_7834; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7836 = 8'h9c == io_state_in_12 ? 8'hbf : _GEN_7835; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7837 = 8'h9d == io_state_in_12 ? 8'hbc : _GEN_7836; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7838 = 8'h9e == io_state_in_12 ? 8'hb9 : _GEN_7837; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7839 = 8'h9f == io_state_in_12 ? 8'hba : _GEN_7838; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7840 = 8'ha0 == io_state_in_12 ? 8'hfb : _GEN_7839; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7841 = 8'ha1 == io_state_in_12 ? 8'hf8 : _GEN_7840; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7842 = 8'ha2 == io_state_in_12 ? 8'hfd : _GEN_7841; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7843 = 8'ha3 == io_state_in_12 ? 8'hfe : _GEN_7842; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7844 = 8'ha4 == io_state_in_12 ? 8'hf7 : _GEN_7843; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7845 = 8'ha5 == io_state_in_12 ? 8'hf4 : _GEN_7844; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7846 = 8'ha6 == io_state_in_12 ? 8'hf1 : _GEN_7845; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7847 = 8'ha7 == io_state_in_12 ? 8'hf2 : _GEN_7846; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7848 = 8'ha8 == io_state_in_12 ? 8'he3 : _GEN_7847; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7849 = 8'ha9 == io_state_in_12 ? 8'he0 : _GEN_7848; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7850 = 8'haa == io_state_in_12 ? 8'he5 : _GEN_7849; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7851 = 8'hab == io_state_in_12 ? 8'he6 : _GEN_7850; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7852 = 8'hac == io_state_in_12 ? 8'hef : _GEN_7851; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7853 = 8'had == io_state_in_12 ? 8'hec : _GEN_7852; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7854 = 8'hae == io_state_in_12 ? 8'he9 : _GEN_7853; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7855 = 8'haf == io_state_in_12 ? 8'hea : _GEN_7854; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7856 = 8'hb0 == io_state_in_12 ? 8'hcb : _GEN_7855; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7857 = 8'hb1 == io_state_in_12 ? 8'hc8 : _GEN_7856; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7858 = 8'hb2 == io_state_in_12 ? 8'hcd : _GEN_7857; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7859 = 8'hb3 == io_state_in_12 ? 8'hce : _GEN_7858; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7860 = 8'hb4 == io_state_in_12 ? 8'hc7 : _GEN_7859; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7861 = 8'hb5 == io_state_in_12 ? 8'hc4 : _GEN_7860; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7862 = 8'hb6 == io_state_in_12 ? 8'hc1 : _GEN_7861; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7863 = 8'hb7 == io_state_in_12 ? 8'hc2 : _GEN_7862; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7864 = 8'hb8 == io_state_in_12 ? 8'hd3 : _GEN_7863; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7865 = 8'hb9 == io_state_in_12 ? 8'hd0 : _GEN_7864; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7866 = 8'hba == io_state_in_12 ? 8'hd5 : _GEN_7865; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7867 = 8'hbb == io_state_in_12 ? 8'hd6 : _GEN_7866; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7868 = 8'hbc == io_state_in_12 ? 8'hdf : _GEN_7867; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7869 = 8'hbd == io_state_in_12 ? 8'hdc : _GEN_7868; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7870 = 8'hbe == io_state_in_12 ? 8'hd9 : _GEN_7869; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7871 = 8'hbf == io_state_in_12 ? 8'hda : _GEN_7870; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7872 = 8'hc0 == io_state_in_12 ? 8'h5b : _GEN_7871; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7873 = 8'hc1 == io_state_in_12 ? 8'h58 : _GEN_7872; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7874 = 8'hc2 == io_state_in_12 ? 8'h5d : _GEN_7873; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7875 = 8'hc3 == io_state_in_12 ? 8'h5e : _GEN_7874; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7876 = 8'hc4 == io_state_in_12 ? 8'h57 : _GEN_7875; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7877 = 8'hc5 == io_state_in_12 ? 8'h54 : _GEN_7876; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7878 = 8'hc6 == io_state_in_12 ? 8'h51 : _GEN_7877; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7879 = 8'hc7 == io_state_in_12 ? 8'h52 : _GEN_7878; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7880 = 8'hc8 == io_state_in_12 ? 8'h43 : _GEN_7879; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7881 = 8'hc9 == io_state_in_12 ? 8'h40 : _GEN_7880; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7882 = 8'hca == io_state_in_12 ? 8'h45 : _GEN_7881; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7883 = 8'hcb == io_state_in_12 ? 8'h46 : _GEN_7882; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7884 = 8'hcc == io_state_in_12 ? 8'h4f : _GEN_7883; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7885 = 8'hcd == io_state_in_12 ? 8'h4c : _GEN_7884; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7886 = 8'hce == io_state_in_12 ? 8'h49 : _GEN_7885; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7887 = 8'hcf == io_state_in_12 ? 8'h4a : _GEN_7886; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7888 = 8'hd0 == io_state_in_12 ? 8'h6b : _GEN_7887; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7889 = 8'hd1 == io_state_in_12 ? 8'h68 : _GEN_7888; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7890 = 8'hd2 == io_state_in_12 ? 8'h6d : _GEN_7889; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7891 = 8'hd3 == io_state_in_12 ? 8'h6e : _GEN_7890; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7892 = 8'hd4 == io_state_in_12 ? 8'h67 : _GEN_7891; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7893 = 8'hd5 == io_state_in_12 ? 8'h64 : _GEN_7892; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7894 = 8'hd6 == io_state_in_12 ? 8'h61 : _GEN_7893; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7895 = 8'hd7 == io_state_in_12 ? 8'h62 : _GEN_7894; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7896 = 8'hd8 == io_state_in_12 ? 8'h73 : _GEN_7895; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7897 = 8'hd9 == io_state_in_12 ? 8'h70 : _GEN_7896; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7898 = 8'hda == io_state_in_12 ? 8'h75 : _GEN_7897; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7899 = 8'hdb == io_state_in_12 ? 8'h76 : _GEN_7898; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7900 = 8'hdc == io_state_in_12 ? 8'h7f : _GEN_7899; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7901 = 8'hdd == io_state_in_12 ? 8'h7c : _GEN_7900; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7902 = 8'hde == io_state_in_12 ? 8'h79 : _GEN_7901; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7903 = 8'hdf == io_state_in_12 ? 8'h7a : _GEN_7902; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7904 = 8'he0 == io_state_in_12 ? 8'h3b : _GEN_7903; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7905 = 8'he1 == io_state_in_12 ? 8'h38 : _GEN_7904; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7906 = 8'he2 == io_state_in_12 ? 8'h3d : _GEN_7905; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7907 = 8'he3 == io_state_in_12 ? 8'h3e : _GEN_7906; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7908 = 8'he4 == io_state_in_12 ? 8'h37 : _GEN_7907; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7909 = 8'he5 == io_state_in_12 ? 8'h34 : _GEN_7908; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7910 = 8'he6 == io_state_in_12 ? 8'h31 : _GEN_7909; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7911 = 8'he7 == io_state_in_12 ? 8'h32 : _GEN_7910; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7912 = 8'he8 == io_state_in_12 ? 8'h23 : _GEN_7911; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7913 = 8'he9 == io_state_in_12 ? 8'h20 : _GEN_7912; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7914 = 8'hea == io_state_in_12 ? 8'h25 : _GEN_7913; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7915 = 8'heb == io_state_in_12 ? 8'h26 : _GEN_7914; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7916 = 8'hec == io_state_in_12 ? 8'h2f : _GEN_7915; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7917 = 8'hed == io_state_in_12 ? 8'h2c : _GEN_7916; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7918 = 8'hee == io_state_in_12 ? 8'h29 : _GEN_7917; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7919 = 8'hef == io_state_in_12 ? 8'h2a : _GEN_7918; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7920 = 8'hf0 == io_state_in_12 ? 8'hb : _GEN_7919; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7921 = 8'hf1 == io_state_in_12 ? 8'h8 : _GEN_7920; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7922 = 8'hf2 == io_state_in_12 ? 8'hd : _GEN_7921; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7923 = 8'hf3 == io_state_in_12 ? 8'he : _GEN_7922; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7924 = 8'hf4 == io_state_in_12 ? 8'h7 : _GEN_7923; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7925 = 8'hf5 == io_state_in_12 ? 8'h4 : _GEN_7924; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7926 = 8'hf6 == io_state_in_12 ? 8'h1 : _GEN_7925; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7927 = 8'hf7 == io_state_in_12 ? 8'h2 : _GEN_7926; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7928 = 8'hf8 == io_state_in_12 ? 8'h13 : _GEN_7927; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7929 = 8'hf9 == io_state_in_12 ? 8'h10 : _GEN_7928; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7930 = 8'hfa == io_state_in_12 ? 8'h15 : _GEN_7929; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7931 = 8'hfb == io_state_in_12 ? 8'h16 : _GEN_7930; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7932 = 8'hfc == io_state_in_12 ? 8'h1f : _GEN_7931; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7933 = 8'hfd == io_state_in_12 ? 8'h1c : _GEN_7932; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7934 = 8'hfe == io_state_in_12 ? 8'h19 : _GEN_7933; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _GEN_7935 = 8'hff == io_state_in_12 ? 8'h1a : _GEN_7934; // @[MixColumns.scala 143:{43,43}]
  wire [7:0] _tmp_state_15_T = _GEN_7935 ^ io_state_in_13; // @[MixColumns.scala 143:43]
  wire [7:0] _tmp_state_15_T_1 = _tmp_state_15_T ^ io_state_in_14; // @[MixColumns.scala 143:61]
  wire [7:0] _GEN_7937 = 8'h1 == io_state_in_15 ? 8'h2 : 8'h0; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7938 = 8'h2 == io_state_in_15 ? 8'h4 : _GEN_7937; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7939 = 8'h3 == io_state_in_15 ? 8'h6 : _GEN_7938; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7940 = 8'h4 == io_state_in_15 ? 8'h8 : _GEN_7939; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7941 = 8'h5 == io_state_in_15 ? 8'ha : _GEN_7940; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7942 = 8'h6 == io_state_in_15 ? 8'hc : _GEN_7941; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7943 = 8'h7 == io_state_in_15 ? 8'he : _GEN_7942; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7944 = 8'h8 == io_state_in_15 ? 8'h10 : _GEN_7943; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7945 = 8'h9 == io_state_in_15 ? 8'h12 : _GEN_7944; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7946 = 8'ha == io_state_in_15 ? 8'h14 : _GEN_7945; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7947 = 8'hb == io_state_in_15 ? 8'h16 : _GEN_7946; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7948 = 8'hc == io_state_in_15 ? 8'h18 : _GEN_7947; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7949 = 8'hd == io_state_in_15 ? 8'h1a : _GEN_7948; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7950 = 8'he == io_state_in_15 ? 8'h1c : _GEN_7949; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7951 = 8'hf == io_state_in_15 ? 8'h1e : _GEN_7950; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7952 = 8'h10 == io_state_in_15 ? 8'h20 : _GEN_7951; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7953 = 8'h11 == io_state_in_15 ? 8'h22 : _GEN_7952; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7954 = 8'h12 == io_state_in_15 ? 8'h24 : _GEN_7953; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7955 = 8'h13 == io_state_in_15 ? 8'h26 : _GEN_7954; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7956 = 8'h14 == io_state_in_15 ? 8'h28 : _GEN_7955; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7957 = 8'h15 == io_state_in_15 ? 8'h2a : _GEN_7956; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7958 = 8'h16 == io_state_in_15 ? 8'h2c : _GEN_7957; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7959 = 8'h17 == io_state_in_15 ? 8'h2e : _GEN_7958; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7960 = 8'h18 == io_state_in_15 ? 8'h30 : _GEN_7959; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7961 = 8'h19 == io_state_in_15 ? 8'h32 : _GEN_7960; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7962 = 8'h1a == io_state_in_15 ? 8'h34 : _GEN_7961; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7963 = 8'h1b == io_state_in_15 ? 8'h36 : _GEN_7962; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7964 = 8'h1c == io_state_in_15 ? 8'h38 : _GEN_7963; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7965 = 8'h1d == io_state_in_15 ? 8'h3a : _GEN_7964; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7966 = 8'h1e == io_state_in_15 ? 8'h3c : _GEN_7965; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7967 = 8'h1f == io_state_in_15 ? 8'h3e : _GEN_7966; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7968 = 8'h20 == io_state_in_15 ? 8'h40 : _GEN_7967; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7969 = 8'h21 == io_state_in_15 ? 8'h42 : _GEN_7968; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7970 = 8'h22 == io_state_in_15 ? 8'h44 : _GEN_7969; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7971 = 8'h23 == io_state_in_15 ? 8'h46 : _GEN_7970; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7972 = 8'h24 == io_state_in_15 ? 8'h48 : _GEN_7971; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7973 = 8'h25 == io_state_in_15 ? 8'h4a : _GEN_7972; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7974 = 8'h26 == io_state_in_15 ? 8'h4c : _GEN_7973; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7975 = 8'h27 == io_state_in_15 ? 8'h4e : _GEN_7974; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7976 = 8'h28 == io_state_in_15 ? 8'h50 : _GEN_7975; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7977 = 8'h29 == io_state_in_15 ? 8'h52 : _GEN_7976; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7978 = 8'h2a == io_state_in_15 ? 8'h54 : _GEN_7977; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7979 = 8'h2b == io_state_in_15 ? 8'h56 : _GEN_7978; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7980 = 8'h2c == io_state_in_15 ? 8'h58 : _GEN_7979; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7981 = 8'h2d == io_state_in_15 ? 8'h5a : _GEN_7980; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7982 = 8'h2e == io_state_in_15 ? 8'h5c : _GEN_7981; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7983 = 8'h2f == io_state_in_15 ? 8'h5e : _GEN_7982; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7984 = 8'h30 == io_state_in_15 ? 8'h60 : _GEN_7983; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7985 = 8'h31 == io_state_in_15 ? 8'h62 : _GEN_7984; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7986 = 8'h32 == io_state_in_15 ? 8'h64 : _GEN_7985; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7987 = 8'h33 == io_state_in_15 ? 8'h66 : _GEN_7986; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7988 = 8'h34 == io_state_in_15 ? 8'h68 : _GEN_7987; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7989 = 8'h35 == io_state_in_15 ? 8'h6a : _GEN_7988; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7990 = 8'h36 == io_state_in_15 ? 8'h6c : _GEN_7989; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7991 = 8'h37 == io_state_in_15 ? 8'h6e : _GEN_7990; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7992 = 8'h38 == io_state_in_15 ? 8'h70 : _GEN_7991; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7993 = 8'h39 == io_state_in_15 ? 8'h72 : _GEN_7992; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7994 = 8'h3a == io_state_in_15 ? 8'h74 : _GEN_7993; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7995 = 8'h3b == io_state_in_15 ? 8'h76 : _GEN_7994; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7996 = 8'h3c == io_state_in_15 ? 8'h78 : _GEN_7995; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7997 = 8'h3d == io_state_in_15 ? 8'h7a : _GEN_7996; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7998 = 8'h3e == io_state_in_15 ? 8'h7c : _GEN_7997; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_7999 = 8'h3f == io_state_in_15 ? 8'h7e : _GEN_7998; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8000 = 8'h40 == io_state_in_15 ? 8'h80 : _GEN_7999; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8001 = 8'h41 == io_state_in_15 ? 8'h82 : _GEN_8000; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8002 = 8'h42 == io_state_in_15 ? 8'h84 : _GEN_8001; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8003 = 8'h43 == io_state_in_15 ? 8'h86 : _GEN_8002; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8004 = 8'h44 == io_state_in_15 ? 8'h88 : _GEN_8003; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8005 = 8'h45 == io_state_in_15 ? 8'h8a : _GEN_8004; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8006 = 8'h46 == io_state_in_15 ? 8'h8c : _GEN_8005; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8007 = 8'h47 == io_state_in_15 ? 8'h8e : _GEN_8006; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8008 = 8'h48 == io_state_in_15 ? 8'h90 : _GEN_8007; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8009 = 8'h49 == io_state_in_15 ? 8'h92 : _GEN_8008; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8010 = 8'h4a == io_state_in_15 ? 8'h94 : _GEN_8009; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8011 = 8'h4b == io_state_in_15 ? 8'h96 : _GEN_8010; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8012 = 8'h4c == io_state_in_15 ? 8'h98 : _GEN_8011; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8013 = 8'h4d == io_state_in_15 ? 8'h9a : _GEN_8012; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8014 = 8'h4e == io_state_in_15 ? 8'h9c : _GEN_8013; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8015 = 8'h4f == io_state_in_15 ? 8'h9e : _GEN_8014; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8016 = 8'h50 == io_state_in_15 ? 8'ha0 : _GEN_8015; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8017 = 8'h51 == io_state_in_15 ? 8'ha2 : _GEN_8016; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8018 = 8'h52 == io_state_in_15 ? 8'ha4 : _GEN_8017; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8019 = 8'h53 == io_state_in_15 ? 8'ha6 : _GEN_8018; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8020 = 8'h54 == io_state_in_15 ? 8'ha8 : _GEN_8019; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8021 = 8'h55 == io_state_in_15 ? 8'haa : _GEN_8020; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8022 = 8'h56 == io_state_in_15 ? 8'hac : _GEN_8021; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8023 = 8'h57 == io_state_in_15 ? 8'hae : _GEN_8022; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8024 = 8'h58 == io_state_in_15 ? 8'hb0 : _GEN_8023; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8025 = 8'h59 == io_state_in_15 ? 8'hb2 : _GEN_8024; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8026 = 8'h5a == io_state_in_15 ? 8'hb4 : _GEN_8025; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8027 = 8'h5b == io_state_in_15 ? 8'hb6 : _GEN_8026; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8028 = 8'h5c == io_state_in_15 ? 8'hb8 : _GEN_8027; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8029 = 8'h5d == io_state_in_15 ? 8'hba : _GEN_8028; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8030 = 8'h5e == io_state_in_15 ? 8'hbc : _GEN_8029; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8031 = 8'h5f == io_state_in_15 ? 8'hbe : _GEN_8030; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8032 = 8'h60 == io_state_in_15 ? 8'hc0 : _GEN_8031; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8033 = 8'h61 == io_state_in_15 ? 8'hc2 : _GEN_8032; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8034 = 8'h62 == io_state_in_15 ? 8'hc4 : _GEN_8033; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8035 = 8'h63 == io_state_in_15 ? 8'hc6 : _GEN_8034; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8036 = 8'h64 == io_state_in_15 ? 8'hc8 : _GEN_8035; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8037 = 8'h65 == io_state_in_15 ? 8'hca : _GEN_8036; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8038 = 8'h66 == io_state_in_15 ? 8'hcc : _GEN_8037; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8039 = 8'h67 == io_state_in_15 ? 8'hce : _GEN_8038; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8040 = 8'h68 == io_state_in_15 ? 8'hd0 : _GEN_8039; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8041 = 8'h69 == io_state_in_15 ? 8'hd2 : _GEN_8040; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8042 = 8'h6a == io_state_in_15 ? 8'hd4 : _GEN_8041; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8043 = 8'h6b == io_state_in_15 ? 8'hd6 : _GEN_8042; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8044 = 8'h6c == io_state_in_15 ? 8'hd8 : _GEN_8043; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8045 = 8'h6d == io_state_in_15 ? 8'hda : _GEN_8044; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8046 = 8'h6e == io_state_in_15 ? 8'hdc : _GEN_8045; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8047 = 8'h6f == io_state_in_15 ? 8'hde : _GEN_8046; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8048 = 8'h70 == io_state_in_15 ? 8'he0 : _GEN_8047; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8049 = 8'h71 == io_state_in_15 ? 8'he2 : _GEN_8048; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8050 = 8'h72 == io_state_in_15 ? 8'he4 : _GEN_8049; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8051 = 8'h73 == io_state_in_15 ? 8'he6 : _GEN_8050; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8052 = 8'h74 == io_state_in_15 ? 8'he8 : _GEN_8051; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8053 = 8'h75 == io_state_in_15 ? 8'hea : _GEN_8052; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8054 = 8'h76 == io_state_in_15 ? 8'hec : _GEN_8053; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8055 = 8'h77 == io_state_in_15 ? 8'hee : _GEN_8054; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8056 = 8'h78 == io_state_in_15 ? 8'hf0 : _GEN_8055; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8057 = 8'h79 == io_state_in_15 ? 8'hf2 : _GEN_8056; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8058 = 8'h7a == io_state_in_15 ? 8'hf4 : _GEN_8057; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8059 = 8'h7b == io_state_in_15 ? 8'hf6 : _GEN_8058; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8060 = 8'h7c == io_state_in_15 ? 8'hf8 : _GEN_8059; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8061 = 8'h7d == io_state_in_15 ? 8'hfa : _GEN_8060; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8062 = 8'h7e == io_state_in_15 ? 8'hfc : _GEN_8061; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8063 = 8'h7f == io_state_in_15 ? 8'hfe : _GEN_8062; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8064 = 8'h80 == io_state_in_15 ? 8'h1b : _GEN_8063; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8065 = 8'h81 == io_state_in_15 ? 8'h19 : _GEN_8064; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8066 = 8'h82 == io_state_in_15 ? 8'h1f : _GEN_8065; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8067 = 8'h83 == io_state_in_15 ? 8'h1d : _GEN_8066; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8068 = 8'h84 == io_state_in_15 ? 8'h13 : _GEN_8067; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8069 = 8'h85 == io_state_in_15 ? 8'h11 : _GEN_8068; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8070 = 8'h86 == io_state_in_15 ? 8'h17 : _GEN_8069; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8071 = 8'h87 == io_state_in_15 ? 8'h15 : _GEN_8070; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8072 = 8'h88 == io_state_in_15 ? 8'hb : _GEN_8071; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8073 = 8'h89 == io_state_in_15 ? 8'h9 : _GEN_8072; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8074 = 8'h8a == io_state_in_15 ? 8'hf : _GEN_8073; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8075 = 8'h8b == io_state_in_15 ? 8'hd : _GEN_8074; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8076 = 8'h8c == io_state_in_15 ? 8'h3 : _GEN_8075; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8077 = 8'h8d == io_state_in_15 ? 8'h1 : _GEN_8076; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8078 = 8'h8e == io_state_in_15 ? 8'h7 : _GEN_8077; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8079 = 8'h8f == io_state_in_15 ? 8'h5 : _GEN_8078; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8080 = 8'h90 == io_state_in_15 ? 8'h3b : _GEN_8079; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8081 = 8'h91 == io_state_in_15 ? 8'h39 : _GEN_8080; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8082 = 8'h92 == io_state_in_15 ? 8'h3f : _GEN_8081; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8083 = 8'h93 == io_state_in_15 ? 8'h3d : _GEN_8082; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8084 = 8'h94 == io_state_in_15 ? 8'h33 : _GEN_8083; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8085 = 8'h95 == io_state_in_15 ? 8'h31 : _GEN_8084; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8086 = 8'h96 == io_state_in_15 ? 8'h37 : _GEN_8085; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8087 = 8'h97 == io_state_in_15 ? 8'h35 : _GEN_8086; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8088 = 8'h98 == io_state_in_15 ? 8'h2b : _GEN_8087; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8089 = 8'h99 == io_state_in_15 ? 8'h29 : _GEN_8088; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8090 = 8'h9a == io_state_in_15 ? 8'h2f : _GEN_8089; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8091 = 8'h9b == io_state_in_15 ? 8'h2d : _GEN_8090; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8092 = 8'h9c == io_state_in_15 ? 8'h23 : _GEN_8091; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8093 = 8'h9d == io_state_in_15 ? 8'h21 : _GEN_8092; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8094 = 8'h9e == io_state_in_15 ? 8'h27 : _GEN_8093; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8095 = 8'h9f == io_state_in_15 ? 8'h25 : _GEN_8094; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8096 = 8'ha0 == io_state_in_15 ? 8'h5b : _GEN_8095; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8097 = 8'ha1 == io_state_in_15 ? 8'h59 : _GEN_8096; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8098 = 8'ha2 == io_state_in_15 ? 8'h5f : _GEN_8097; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8099 = 8'ha3 == io_state_in_15 ? 8'h5d : _GEN_8098; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8100 = 8'ha4 == io_state_in_15 ? 8'h53 : _GEN_8099; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8101 = 8'ha5 == io_state_in_15 ? 8'h51 : _GEN_8100; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8102 = 8'ha6 == io_state_in_15 ? 8'h57 : _GEN_8101; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8103 = 8'ha7 == io_state_in_15 ? 8'h55 : _GEN_8102; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8104 = 8'ha8 == io_state_in_15 ? 8'h4b : _GEN_8103; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8105 = 8'ha9 == io_state_in_15 ? 8'h49 : _GEN_8104; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8106 = 8'haa == io_state_in_15 ? 8'h4f : _GEN_8105; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8107 = 8'hab == io_state_in_15 ? 8'h4d : _GEN_8106; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8108 = 8'hac == io_state_in_15 ? 8'h43 : _GEN_8107; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8109 = 8'had == io_state_in_15 ? 8'h41 : _GEN_8108; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8110 = 8'hae == io_state_in_15 ? 8'h47 : _GEN_8109; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8111 = 8'haf == io_state_in_15 ? 8'h45 : _GEN_8110; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8112 = 8'hb0 == io_state_in_15 ? 8'h7b : _GEN_8111; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8113 = 8'hb1 == io_state_in_15 ? 8'h79 : _GEN_8112; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8114 = 8'hb2 == io_state_in_15 ? 8'h7f : _GEN_8113; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8115 = 8'hb3 == io_state_in_15 ? 8'h7d : _GEN_8114; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8116 = 8'hb4 == io_state_in_15 ? 8'h73 : _GEN_8115; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8117 = 8'hb5 == io_state_in_15 ? 8'h71 : _GEN_8116; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8118 = 8'hb6 == io_state_in_15 ? 8'h77 : _GEN_8117; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8119 = 8'hb7 == io_state_in_15 ? 8'h75 : _GEN_8118; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8120 = 8'hb8 == io_state_in_15 ? 8'h6b : _GEN_8119; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8121 = 8'hb9 == io_state_in_15 ? 8'h69 : _GEN_8120; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8122 = 8'hba == io_state_in_15 ? 8'h6f : _GEN_8121; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8123 = 8'hbb == io_state_in_15 ? 8'h6d : _GEN_8122; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8124 = 8'hbc == io_state_in_15 ? 8'h63 : _GEN_8123; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8125 = 8'hbd == io_state_in_15 ? 8'h61 : _GEN_8124; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8126 = 8'hbe == io_state_in_15 ? 8'h67 : _GEN_8125; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8127 = 8'hbf == io_state_in_15 ? 8'h65 : _GEN_8126; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8128 = 8'hc0 == io_state_in_15 ? 8'h9b : _GEN_8127; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8129 = 8'hc1 == io_state_in_15 ? 8'h99 : _GEN_8128; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8130 = 8'hc2 == io_state_in_15 ? 8'h9f : _GEN_8129; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8131 = 8'hc3 == io_state_in_15 ? 8'h9d : _GEN_8130; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8132 = 8'hc4 == io_state_in_15 ? 8'h93 : _GEN_8131; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8133 = 8'hc5 == io_state_in_15 ? 8'h91 : _GEN_8132; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8134 = 8'hc6 == io_state_in_15 ? 8'h97 : _GEN_8133; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8135 = 8'hc7 == io_state_in_15 ? 8'h95 : _GEN_8134; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8136 = 8'hc8 == io_state_in_15 ? 8'h8b : _GEN_8135; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8137 = 8'hc9 == io_state_in_15 ? 8'h89 : _GEN_8136; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8138 = 8'hca == io_state_in_15 ? 8'h8f : _GEN_8137; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8139 = 8'hcb == io_state_in_15 ? 8'h8d : _GEN_8138; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8140 = 8'hcc == io_state_in_15 ? 8'h83 : _GEN_8139; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8141 = 8'hcd == io_state_in_15 ? 8'h81 : _GEN_8140; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8142 = 8'hce == io_state_in_15 ? 8'h87 : _GEN_8141; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8143 = 8'hcf == io_state_in_15 ? 8'h85 : _GEN_8142; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8144 = 8'hd0 == io_state_in_15 ? 8'hbb : _GEN_8143; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8145 = 8'hd1 == io_state_in_15 ? 8'hb9 : _GEN_8144; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8146 = 8'hd2 == io_state_in_15 ? 8'hbf : _GEN_8145; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8147 = 8'hd3 == io_state_in_15 ? 8'hbd : _GEN_8146; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8148 = 8'hd4 == io_state_in_15 ? 8'hb3 : _GEN_8147; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8149 = 8'hd5 == io_state_in_15 ? 8'hb1 : _GEN_8148; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8150 = 8'hd6 == io_state_in_15 ? 8'hb7 : _GEN_8149; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8151 = 8'hd7 == io_state_in_15 ? 8'hb5 : _GEN_8150; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8152 = 8'hd8 == io_state_in_15 ? 8'hab : _GEN_8151; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8153 = 8'hd9 == io_state_in_15 ? 8'ha9 : _GEN_8152; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8154 = 8'hda == io_state_in_15 ? 8'haf : _GEN_8153; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8155 = 8'hdb == io_state_in_15 ? 8'had : _GEN_8154; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8156 = 8'hdc == io_state_in_15 ? 8'ha3 : _GEN_8155; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8157 = 8'hdd == io_state_in_15 ? 8'ha1 : _GEN_8156; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8158 = 8'hde == io_state_in_15 ? 8'ha7 : _GEN_8157; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8159 = 8'hdf == io_state_in_15 ? 8'ha5 : _GEN_8158; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8160 = 8'he0 == io_state_in_15 ? 8'hdb : _GEN_8159; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8161 = 8'he1 == io_state_in_15 ? 8'hd9 : _GEN_8160; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8162 = 8'he2 == io_state_in_15 ? 8'hdf : _GEN_8161; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8163 = 8'he3 == io_state_in_15 ? 8'hdd : _GEN_8162; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8164 = 8'he4 == io_state_in_15 ? 8'hd3 : _GEN_8163; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8165 = 8'he5 == io_state_in_15 ? 8'hd1 : _GEN_8164; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8166 = 8'he6 == io_state_in_15 ? 8'hd7 : _GEN_8165; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8167 = 8'he7 == io_state_in_15 ? 8'hd5 : _GEN_8166; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8168 = 8'he8 == io_state_in_15 ? 8'hcb : _GEN_8167; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8169 = 8'he9 == io_state_in_15 ? 8'hc9 : _GEN_8168; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8170 = 8'hea == io_state_in_15 ? 8'hcf : _GEN_8169; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8171 = 8'heb == io_state_in_15 ? 8'hcd : _GEN_8170; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8172 = 8'hec == io_state_in_15 ? 8'hc3 : _GEN_8171; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8173 = 8'hed == io_state_in_15 ? 8'hc1 : _GEN_8172; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8174 = 8'hee == io_state_in_15 ? 8'hc7 : _GEN_8173; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8175 = 8'hef == io_state_in_15 ? 8'hc5 : _GEN_8174; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8176 = 8'hf0 == io_state_in_15 ? 8'hfb : _GEN_8175; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8177 = 8'hf1 == io_state_in_15 ? 8'hf9 : _GEN_8176; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8178 = 8'hf2 == io_state_in_15 ? 8'hff : _GEN_8177; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8179 = 8'hf3 == io_state_in_15 ? 8'hfd : _GEN_8178; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8180 = 8'hf4 == io_state_in_15 ? 8'hf3 : _GEN_8179; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8181 = 8'hf5 == io_state_in_15 ? 8'hf1 : _GEN_8180; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8182 = 8'hf6 == io_state_in_15 ? 8'hf7 : _GEN_8181; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8183 = 8'hf7 == io_state_in_15 ? 8'hf5 : _GEN_8182; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8184 = 8'hf8 == io_state_in_15 ? 8'heb : _GEN_8183; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8185 = 8'hf9 == io_state_in_15 ? 8'he9 : _GEN_8184; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8186 = 8'hfa == io_state_in_15 ? 8'hef : _GEN_8185; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8187 = 8'hfb == io_state_in_15 ? 8'hed : _GEN_8186; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8188 = 8'hfc == io_state_in_15 ? 8'he3 : _GEN_8187; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8189 = 8'hfd == io_state_in_15 ? 8'he1 : _GEN_8188; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8190 = 8'hfe == io_state_in_15 ? 8'he7 : _GEN_8189; // @[MixColumns.scala 143:{79,79}]
  wire [7:0] _GEN_8191 = 8'hff == io_state_in_15 ? 8'he5 : _GEN_8190; // @[MixColumns.scala 143:{79,79}]
  assign io_state_out_0 = _tmp_state_0_T_1 ^ io_state_in_3; // @[MixColumns.scala 125:82]
  assign io_state_out_1 = _tmp_state_1_T_1 ^ io_state_in_3; // @[MixColumns.scala 126:82]
  assign io_state_out_2 = _tmp_state_2_T_1 ^ _GEN_1535; // @[MixColumns.scala 127:75]
  assign io_state_out_3 = _tmp_state_3_T_1 ^ _GEN_2047; // @[MixColumns.scala 128:75]
  assign io_state_out_4 = _tmp_state_4_T_1 ^ io_state_in_7; // @[MixColumns.scala 130:82]
  assign io_state_out_5 = _tmp_state_5_T_1 ^ io_state_in_7; // @[MixColumns.scala 131:82]
  assign io_state_out_6 = _tmp_state_6_T_1 ^ _GEN_3583; // @[MixColumns.scala 132:75]
  assign io_state_out_7 = _tmp_state_7_T_1 ^ _GEN_4095; // @[MixColumns.scala 133:75]
  assign io_state_out_8 = _tmp_state_8_T_1 ^ io_state_in_11; // @[MixColumns.scala 135:83]
  assign io_state_out_9 = _tmp_state_9_T_1 ^ io_state_in_11; // @[MixColumns.scala 136:83]
  assign io_state_out_10 = _tmp_state_10_T_1 ^ _GEN_5631; // @[MixColumns.scala 137:77]
  assign io_state_out_11 = _tmp_state_11_T_1 ^ _GEN_6143; // @[MixColumns.scala 138:77]
  assign io_state_out_12 = _tmp_state_12_T_1 ^ io_state_in_15; // @[MixColumns.scala 140:86]
  assign io_state_out_13 = _tmp_state_13_T_1 ^ io_state_in_15; // @[MixColumns.scala 141:86]
  assign io_state_out_14 = _tmp_state_14_T_1 ^ _GEN_7679; // @[MixColumns.scala 142:79]
  assign io_state_out_15 = _tmp_state_15_T_1 ^ _GEN_8191; // @[MixColumns.scala 143:79]
endmodule
module Cipher(
  input        clock,
  input        reset,
  input  [7:0] io_plaintext_0,
  input  [7:0] io_plaintext_1,
  input  [7:0] io_plaintext_2,
  input  [7:0] io_plaintext_3,
  input  [7:0] io_plaintext_4,
  input  [7:0] io_plaintext_5,
  input  [7:0] io_plaintext_6,
  input  [7:0] io_plaintext_7,
  input  [7:0] io_plaintext_8,
  input  [7:0] io_plaintext_9,
  input  [7:0] io_plaintext_10,
  input  [7:0] io_plaintext_11,
  input  [7:0] io_plaintext_12,
  input  [7:0] io_plaintext_13,
  input  [7:0] io_plaintext_14,
  input  [7:0] io_plaintext_15,
  input  [7:0] io_roundKey_0,
  input  [7:0] io_roundKey_1,
  input  [7:0] io_roundKey_2,
  input  [7:0] io_roundKey_3,
  input  [7:0] io_roundKey_4,
  input  [7:0] io_roundKey_5,
  input  [7:0] io_roundKey_6,
  input  [7:0] io_roundKey_7,
  input  [7:0] io_roundKey_8,
  input  [7:0] io_roundKey_9,
  input  [7:0] io_roundKey_10,
  input  [7:0] io_roundKey_11,
  input  [7:0] io_roundKey_12,
  input  [7:0] io_roundKey_13,
  input  [7:0] io_roundKey_14,
  input  [7:0] io_roundKey_15,
  input        io_start,
  output [7:0] io_state_out_0,
  output [7:0] io_state_out_1,
  output [7:0] io_state_out_2,
  output [7:0] io_state_out_3,
  output [7:0] io_state_out_4,
  output [7:0] io_state_out_5,
  output [7:0] io_state_out_6,
  output [7:0] io_state_out_7,
  output [7:0] io_state_out_8,
  output [7:0] io_state_out_9,
  output [7:0] io_state_out_10,
  output [7:0] io_state_out_11,
  output [7:0] io_state_out_12,
  output [7:0] io_state_out_13,
  output [7:0] io_state_out_14,
  output [7:0] io_state_out_15,
  output       io_state_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] AddRoundKeyModule_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire [7:0] AddRoundKeyModule_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire [7:0] SubBytesModule_io_state_in_0; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_1; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_2; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_3; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_4; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_5; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_6; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_7; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_8; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_9; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_10; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_11; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_12; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_13; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_14; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_in_15; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_0; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_1; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_2; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_3; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_4; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_5; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_6; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_7; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_8; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_9; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_10; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_11; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_12; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_13; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_14; // @[SubBytes.scala 41:81]
  wire [7:0] SubBytesModule_io_state_out_15; // @[SubBytes.scala 41:81]
  wire [7:0] ShiftRowsModule_io_state_in_0; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_1; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_2; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_3; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_4; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_5; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_6; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_7; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_8; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_9; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_10; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_11; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_12; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_13; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_14; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_in_15; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_0; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_1; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_2; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_3; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_4; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_5; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_6; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_7; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_8; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_9; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_10; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_11; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_12; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_13; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_14; // @[ShiftRows.scala 35:34]
  wire [7:0] ShiftRowsModule_io_state_out_15; // @[ShiftRows.scala 35:34]
  wire [7:0] MixColumnsModule_io_state_in_0; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_1; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_2; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_3; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_4; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_5; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_6; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_7; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_8; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_9; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_10; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_11; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_12; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_13; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_14; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_in_15; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_0; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_1; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_2; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_3; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_4; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_5; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_6; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_7; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_8; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_9; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_10; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_11; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_12; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_13; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_14; // @[MixColumns.scala 153:61]
  wire [7:0] MixColumnsModule_io_state_out_15; // @[MixColumns.scala 153:61]
  reg [7:0] state_0; // @[Cipher.scala 31:22]
  reg [7:0] state_1; // @[Cipher.scala 31:22]
  reg [7:0] state_2; // @[Cipher.scala 31:22]
  reg [7:0] state_3; // @[Cipher.scala 31:22]
  reg [7:0] state_4; // @[Cipher.scala 31:22]
  reg [7:0] state_5; // @[Cipher.scala 31:22]
  reg [7:0] state_6; // @[Cipher.scala 31:22]
  reg [7:0] state_7; // @[Cipher.scala 31:22]
  reg [7:0] state_8; // @[Cipher.scala 31:22]
  reg [7:0] state_9; // @[Cipher.scala 31:22]
  reg [7:0] state_10; // @[Cipher.scala 31:22]
  reg [7:0] state_11; // @[Cipher.scala 31:22]
  reg [7:0] state_12; // @[Cipher.scala 31:22]
  reg [7:0] state_13; // @[Cipher.scala 31:22]
  reg [7:0] state_14; // @[Cipher.scala 31:22]
  reg [7:0] state_15; // @[Cipher.scala 31:22]
  reg [3:0] rounds; // @[Cipher.scala 32:23]
  reg [1:0] STM; // @[Cipher.scala 36:20]
  wire [3:0] _rounds_T_1 = rounds + 4'h1; // @[Cipher.scala 46:24]
  wire  _T_3 = rounds == 4'ha; // @[Cipher.scala 51:19]
  wire [1:0] _GEN_1 = rounds == 4'ha ? 2'h0 : STM; // @[Cipher.scala 51:29 52:13 36:20]
  wire [7:0] _T_6_0 = _T_3 ? ShiftRowsModule_io_state_out_0 : MixColumnsModule_io_state_out_0; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_1 = _T_3 ? ShiftRowsModule_io_state_out_1 : MixColumnsModule_io_state_out_1; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_2 = _T_3 ? ShiftRowsModule_io_state_out_2 : MixColumnsModule_io_state_out_2; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_3 = _T_3 ? ShiftRowsModule_io_state_out_3 : MixColumnsModule_io_state_out_3; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_4 = _T_3 ? ShiftRowsModule_io_state_out_4 : MixColumnsModule_io_state_out_4; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_5 = _T_3 ? ShiftRowsModule_io_state_out_5 : MixColumnsModule_io_state_out_5; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_6 = _T_3 ? ShiftRowsModule_io_state_out_6 : MixColumnsModule_io_state_out_6; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_7 = _T_3 ? ShiftRowsModule_io_state_out_7 : MixColumnsModule_io_state_out_7; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_8 = _T_3 ? ShiftRowsModule_io_state_out_8 : MixColumnsModule_io_state_out_8; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_9 = _T_3 ? ShiftRowsModule_io_state_out_9 : MixColumnsModule_io_state_out_9; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_10 = _T_3 ? ShiftRowsModule_io_state_out_10 : MixColumnsModule_io_state_out_10; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_11 = _T_3 ? ShiftRowsModule_io_state_out_11 : MixColumnsModule_io_state_out_11; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_12 = _T_3 ? ShiftRowsModule_io_state_out_12 : MixColumnsModule_io_state_out_12; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_13 = _T_3 ? ShiftRowsModule_io_state_out_13 : MixColumnsModule_io_state_out_13; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_14 = _T_3 ? ShiftRowsModule_io_state_out_14 : MixColumnsModule_io_state_out_14; // @[Cipher.scala 68:8]
  wire [7:0] _T_6_15 = _T_3 ? ShiftRowsModule_io_state_out_15 : MixColumnsModule_io_state_out_15; // @[Cipher.scala 68:8]
  wire  _io_state_out_valid_T = rounds == 4'hb; // @[Cipher.scala 74:32]
  AddRoundKey AddRoundKeyModule ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKeyModule_io_state_in_0),
    .io_state_in_1(AddRoundKeyModule_io_state_in_1),
    .io_state_in_2(AddRoundKeyModule_io_state_in_2),
    .io_state_in_3(AddRoundKeyModule_io_state_in_3),
    .io_state_in_4(AddRoundKeyModule_io_state_in_4),
    .io_state_in_5(AddRoundKeyModule_io_state_in_5),
    .io_state_in_6(AddRoundKeyModule_io_state_in_6),
    .io_state_in_7(AddRoundKeyModule_io_state_in_7),
    .io_state_in_8(AddRoundKeyModule_io_state_in_8),
    .io_state_in_9(AddRoundKeyModule_io_state_in_9),
    .io_state_in_10(AddRoundKeyModule_io_state_in_10),
    .io_state_in_11(AddRoundKeyModule_io_state_in_11),
    .io_state_in_12(AddRoundKeyModule_io_state_in_12),
    .io_state_in_13(AddRoundKeyModule_io_state_in_13),
    .io_state_in_14(AddRoundKeyModule_io_state_in_14),
    .io_state_in_15(AddRoundKeyModule_io_state_in_15),
    .io_roundKey_0(AddRoundKeyModule_io_roundKey_0),
    .io_roundKey_1(AddRoundKeyModule_io_roundKey_1),
    .io_roundKey_2(AddRoundKeyModule_io_roundKey_2),
    .io_roundKey_3(AddRoundKeyModule_io_roundKey_3),
    .io_roundKey_4(AddRoundKeyModule_io_roundKey_4),
    .io_roundKey_5(AddRoundKeyModule_io_roundKey_5),
    .io_roundKey_6(AddRoundKeyModule_io_roundKey_6),
    .io_roundKey_7(AddRoundKeyModule_io_roundKey_7),
    .io_roundKey_8(AddRoundKeyModule_io_roundKey_8),
    .io_roundKey_9(AddRoundKeyModule_io_roundKey_9),
    .io_roundKey_10(AddRoundKeyModule_io_roundKey_10),
    .io_roundKey_11(AddRoundKeyModule_io_roundKey_11),
    .io_roundKey_12(AddRoundKeyModule_io_roundKey_12),
    .io_roundKey_13(AddRoundKeyModule_io_roundKey_13),
    .io_roundKey_14(AddRoundKeyModule_io_roundKey_14),
    .io_roundKey_15(AddRoundKeyModule_io_roundKey_15),
    .io_state_out_0(AddRoundKeyModule_io_state_out_0),
    .io_state_out_1(AddRoundKeyModule_io_state_out_1),
    .io_state_out_2(AddRoundKeyModule_io_state_out_2),
    .io_state_out_3(AddRoundKeyModule_io_state_out_3),
    .io_state_out_4(AddRoundKeyModule_io_state_out_4),
    .io_state_out_5(AddRoundKeyModule_io_state_out_5),
    .io_state_out_6(AddRoundKeyModule_io_state_out_6),
    .io_state_out_7(AddRoundKeyModule_io_state_out_7),
    .io_state_out_8(AddRoundKeyModule_io_state_out_8),
    .io_state_out_9(AddRoundKeyModule_io_state_out_9),
    .io_state_out_10(AddRoundKeyModule_io_state_out_10),
    .io_state_out_11(AddRoundKeyModule_io_state_out_11),
    .io_state_out_12(AddRoundKeyModule_io_state_out_12),
    .io_state_out_13(AddRoundKeyModule_io_state_out_13),
    .io_state_out_14(AddRoundKeyModule_io_state_out_14),
    .io_state_out_15(AddRoundKeyModule_io_state_out_15)
  );
  SubBytes SubBytesModule ( // @[SubBytes.scala 41:81]
    .io_state_in_0(SubBytesModule_io_state_in_0),
    .io_state_in_1(SubBytesModule_io_state_in_1),
    .io_state_in_2(SubBytesModule_io_state_in_2),
    .io_state_in_3(SubBytesModule_io_state_in_3),
    .io_state_in_4(SubBytesModule_io_state_in_4),
    .io_state_in_5(SubBytesModule_io_state_in_5),
    .io_state_in_6(SubBytesModule_io_state_in_6),
    .io_state_in_7(SubBytesModule_io_state_in_7),
    .io_state_in_8(SubBytesModule_io_state_in_8),
    .io_state_in_9(SubBytesModule_io_state_in_9),
    .io_state_in_10(SubBytesModule_io_state_in_10),
    .io_state_in_11(SubBytesModule_io_state_in_11),
    .io_state_in_12(SubBytesModule_io_state_in_12),
    .io_state_in_13(SubBytesModule_io_state_in_13),
    .io_state_in_14(SubBytesModule_io_state_in_14),
    .io_state_in_15(SubBytesModule_io_state_in_15),
    .io_state_out_0(SubBytesModule_io_state_out_0),
    .io_state_out_1(SubBytesModule_io_state_out_1),
    .io_state_out_2(SubBytesModule_io_state_out_2),
    .io_state_out_3(SubBytesModule_io_state_out_3),
    .io_state_out_4(SubBytesModule_io_state_out_4),
    .io_state_out_5(SubBytesModule_io_state_out_5),
    .io_state_out_6(SubBytesModule_io_state_out_6),
    .io_state_out_7(SubBytesModule_io_state_out_7),
    .io_state_out_8(SubBytesModule_io_state_out_8),
    .io_state_out_9(SubBytesModule_io_state_out_9),
    .io_state_out_10(SubBytesModule_io_state_out_10),
    .io_state_out_11(SubBytesModule_io_state_out_11),
    .io_state_out_12(SubBytesModule_io_state_out_12),
    .io_state_out_13(SubBytesModule_io_state_out_13),
    .io_state_out_14(SubBytesModule_io_state_out_14),
    .io_state_out_15(SubBytesModule_io_state_out_15)
  );
  ShiftRows ShiftRowsModule ( // @[ShiftRows.scala 35:34]
    .io_state_in_0(ShiftRowsModule_io_state_in_0),
    .io_state_in_1(ShiftRowsModule_io_state_in_1),
    .io_state_in_2(ShiftRowsModule_io_state_in_2),
    .io_state_in_3(ShiftRowsModule_io_state_in_3),
    .io_state_in_4(ShiftRowsModule_io_state_in_4),
    .io_state_in_5(ShiftRowsModule_io_state_in_5),
    .io_state_in_6(ShiftRowsModule_io_state_in_6),
    .io_state_in_7(ShiftRowsModule_io_state_in_7),
    .io_state_in_8(ShiftRowsModule_io_state_in_8),
    .io_state_in_9(ShiftRowsModule_io_state_in_9),
    .io_state_in_10(ShiftRowsModule_io_state_in_10),
    .io_state_in_11(ShiftRowsModule_io_state_in_11),
    .io_state_in_12(ShiftRowsModule_io_state_in_12),
    .io_state_in_13(ShiftRowsModule_io_state_in_13),
    .io_state_in_14(ShiftRowsModule_io_state_in_14),
    .io_state_in_15(ShiftRowsModule_io_state_in_15),
    .io_state_out_0(ShiftRowsModule_io_state_out_0),
    .io_state_out_1(ShiftRowsModule_io_state_out_1),
    .io_state_out_2(ShiftRowsModule_io_state_out_2),
    .io_state_out_3(ShiftRowsModule_io_state_out_3),
    .io_state_out_4(ShiftRowsModule_io_state_out_4),
    .io_state_out_5(ShiftRowsModule_io_state_out_5),
    .io_state_out_6(ShiftRowsModule_io_state_out_6),
    .io_state_out_7(ShiftRowsModule_io_state_out_7),
    .io_state_out_8(ShiftRowsModule_io_state_out_8),
    .io_state_out_9(ShiftRowsModule_io_state_out_9),
    .io_state_out_10(ShiftRowsModule_io_state_out_10),
    .io_state_out_11(ShiftRowsModule_io_state_out_11),
    .io_state_out_12(ShiftRowsModule_io_state_out_12),
    .io_state_out_13(ShiftRowsModule_io_state_out_13),
    .io_state_out_14(ShiftRowsModule_io_state_out_14),
    .io_state_out_15(ShiftRowsModule_io_state_out_15)
  );
  MixColumns MixColumnsModule ( // @[MixColumns.scala 153:61]
    .io_state_in_0(MixColumnsModule_io_state_in_0),
    .io_state_in_1(MixColumnsModule_io_state_in_1),
    .io_state_in_2(MixColumnsModule_io_state_in_2),
    .io_state_in_3(MixColumnsModule_io_state_in_3),
    .io_state_in_4(MixColumnsModule_io_state_in_4),
    .io_state_in_5(MixColumnsModule_io_state_in_5),
    .io_state_in_6(MixColumnsModule_io_state_in_6),
    .io_state_in_7(MixColumnsModule_io_state_in_7),
    .io_state_in_8(MixColumnsModule_io_state_in_8),
    .io_state_in_9(MixColumnsModule_io_state_in_9),
    .io_state_in_10(MixColumnsModule_io_state_in_10),
    .io_state_in_11(MixColumnsModule_io_state_in_11),
    .io_state_in_12(MixColumnsModule_io_state_in_12),
    .io_state_in_13(MixColumnsModule_io_state_in_13),
    .io_state_in_14(MixColumnsModule_io_state_in_14),
    .io_state_in_15(MixColumnsModule_io_state_in_15),
    .io_state_out_0(MixColumnsModule_io_state_out_0),
    .io_state_out_1(MixColumnsModule_io_state_out_1),
    .io_state_out_2(MixColumnsModule_io_state_out_2),
    .io_state_out_3(MixColumnsModule_io_state_out_3),
    .io_state_out_4(MixColumnsModule_io_state_out_4),
    .io_state_out_5(MixColumnsModule_io_state_out_5),
    .io_state_out_6(MixColumnsModule_io_state_out_6),
    .io_state_out_7(MixColumnsModule_io_state_out_7),
    .io_state_out_8(MixColumnsModule_io_state_out_8),
    .io_state_out_9(MixColumnsModule_io_state_out_9),
    .io_state_out_10(MixColumnsModule_io_state_out_10),
    .io_state_out_11(MixColumnsModule_io_state_out_11),
    .io_state_out_12(MixColumnsModule_io_state_out_12),
    .io_state_out_13(MixColumnsModule_io_state_out_13),
    .io_state_out_14(MixColumnsModule_io_state_out_14),
    .io_state_out_15(MixColumnsModule_io_state_out_15)
  );
  assign io_state_out_0 = _io_state_out_valid_T ? state_0 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_1 = _io_state_out_valid_T ? state_1 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_2 = _io_state_out_valid_T ? state_2 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_3 = _io_state_out_valid_T ? state_3 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_4 = _io_state_out_valid_T ? state_4 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_5 = _io_state_out_valid_T ? state_5 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_6 = _io_state_out_valid_T ? state_6 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_7 = _io_state_out_valid_T ? state_7 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_8 = _io_state_out_valid_T ? state_8 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_9 = _io_state_out_valid_T ? state_9 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_10 = _io_state_out_valid_T ? state_10 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_11 = _io_state_out_valid_T ? state_11 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_12 = _io_state_out_valid_T ? state_12 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_13 = _io_state_out_valid_T ? state_13 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_14 = _io_state_out_valid_T ? state_14 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_15 = _io_state_out_valid_T ? state_15 : 8'h0; // @[Cipher.scala 75:22]
  assign io_state_out_valid = rounds == 4'hb; // @[Cipher.scala 74:32]
  assign AddRoundKeyModule_io_state_in_0 = STM == 2'h1 ? io_plaintext_0 : _T_6_0; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_1 = STM == 2'h1 ? io_plaintext_1 : _T_6_1; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_2 = STM == 2'h1 ? io_plaintext_2 : _T_6_2; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_3 = STM == 2'h1 ? io_plaintext_3 : _T_6_3; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_4 = STM == 2'h1 ? io_plaintext_4 : _T_6_4; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_5 = STM == 2'h1 ? io_plaintext_5 : _T_6_5; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_6 = STM == 2'h1 ? io_plaintext_6 : _T_6_6; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_7 = STM == 2'h1 ? io_plaintext_7 : _T_6_7; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_8 = STM == 2'h1 ? io_plaintext_8 : _T_6_8; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_9 = STM == 2'h1 ? io_plaintext_9 : _T_6_9; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_10 = STM == 2'h1 ? io_plaintext_10 : _T_6_10; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_11 = STM == 2'h1 ? io_plaintext_11 : _T_6_11; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_12 = STM == 2'h1 ? io_plaintext_12 : _T_6_12; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_13 = STM == 2'h1 ? io_plaintext_13 : _T_6_13; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_14 = STM == 2'h1 ? io_plaintext_14 : _T_6_14; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_state_in_15 = STM == 2'h1 ? io_plaintext_15 : _T_6_15; // @[Cipher.scala 67:39]
  assign AddRoundKeyModule_io_roundKey_0 = io_roundKey_0; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_1 = io_roundKey_1; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_2 = io_roundKey_2; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_3 = io_roundKey_3; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_4 = io_roundKey_4; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_5 = io_roundKey_5; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_6 = io_roundKey_6; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_7 = io_roundKey_7; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_8 = io_roundKey_8; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_9 = io_roundKey_9; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_10 = io_roundKey_10; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_11 = io_roundKey_11; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_12 = io_roundKey_12; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_13 = io_roundKey_13; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_14 = io_roundKey_14; // @[Cipher.scala 69:33]
  assign AddRoundKeyModule_io_roundKey_15 = io_roundKey_15; // @[Cipher.scala 69:33]
  assign SubBytesModule_io_state_in_0 = state_0; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_1 = state_1; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_2 = state_2; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_3 = state_3; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_4 = state_4; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_5 = state_5; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_6 = state_6; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_7 = state_7; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_8 = state_8; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_9 = state_9; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_10 = state_10; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_11 = state_11; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_12 = state_12; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_13 = state_13; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_14 = state_14; // @[Cipher.scala 58:30]
  assign SubBytesModule_io_state_in_15 = state_15; // @[Cipher.scala 58:30]
  assign ShiftRowsModule_io_state_in_0 = SubBytesModule_io_state_out_0; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_1 = SubBytesModule_io_state_out_1; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_2 = SubBytesModule_io_state_out_2; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_3 = SubBytesModule_io_state_out_3; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_4 = SubBytesModule_io_state_out_4; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_5 = SubBytesModule_io_state_out_5; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_6 = SubBytesModule_io_state_out_6; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_7 = SubBytesModule_io_state_out_7; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_8 = SubBytesModule_io_state_out_8; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_9 = SubBytesModule_io_state_out_9; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_10 = SubBytesModule_io_state_out_10; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_11 = SubBytesModule_io_state_out_11; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_12 = SubBytesModule_io_state_out_12; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_13 = SubBytesModule_io_state_out_13; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_14 = SubBytesModule_io_state_out_14; // @[Cipher.scala 61:31]
  assign ShiftRowsModule_io_state_in_15 = SubBytesModule_io_state_out_15; // @[Cipher.scala 61:31]
  assign MixColumnsModule_io_state_in_0 = ShiftRowsModule_io_state_out_0; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_1 = ShiftRowsModule_io_state_out_1; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_2 = ShiftRowsModule_io_state_out_2; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_3 = ShiftRowsModule_io_state_out_3; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_4 = ShiftRowsModule_io_state_out_4; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_5 = ShiftRowsModule_io_state_out_5; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_6 = ShiftRowsModule_io_state_out_6; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_7 = ShiftRowsModule_io_state_out_7; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_8 = ShiftRowsModule_io_state_out_8; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_9 = ShiftRowsModule_io_state_out_9; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_10 = ShiftRowsModule_io_state_out_10; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_11 = ShiftRowsModule_io_state_out_11; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_12 = ShiftRowsModule_io_state_out_12; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_13 = ShiftRowsModule_io_state_out_13; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_14 = ShiftRowsModule_io_state_out_14; // @[Cipher.scala 64:32]
  assign MixColumnsModule_io_state_in_15 = ShiftRowsModule_io_state_out_15; // @[Cipher.scala 64:32]
  always @(posedge clock) begin
    if (reset) begin // @[Cipher.scala 31:22]
      state_0 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_0 <= AddRoundKeyModule_io_state_out_0;
    end else begin
      state_0 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_1 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_1 <= AddRoundKeyModule_io_state_out_1;
    end else begin
      state_1 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_2 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_2 <= AddRoundKeyModule_io_state_out_2;
    end else begin
      state_2 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_3 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_3 <= AddRoundKeyModule_io_state_out_3;
    end else begin
      state_3 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_4 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_4 <= AddRoundKeyModule_io_state_out_4;
    end else begin
      state_4 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_5 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_5 <= AddRoundKeyModule_io_state_out_5;
    end else begin
      state_5 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_6 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_6 <= AddRoundKeyModule_io_state_out_6;
    end else begin
      state_6 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_7 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_7 <= AddRoundKeyModule_io_state_out_7;
    end else begin
      state_7 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_8 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_8 <= AddRoundKeyModule_io_state_out_8;
    end else begin
      state_8 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_9 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_9 <= AddRoundKeyModule_io_state_out_9;
    end else begin
      state_9 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_10 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_10 <= AddRoundKeyModule_io_state_out_10;
    end else begin
      state_10 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_11 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_11 <= AddRoundKeyModule_io_state_out_11;
    end else begin
      state_11 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_12 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_12 <= AddRoundKeyModule_io_state_out_12;
    end else begin
      state_12 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_13 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_13 <= AddRoundKeyModule_io_state_out_13;
    end else begin
      state_13 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_14 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_14 <= AddRoundKeyModule_io_state_out_14;
    end else begin
      state_14 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 31:22]
      state_15 <= 8'h0; // @[Cipher.scala 31:22]
    end else if (STM != 2'h0) begin // @[Cipher.scala 71:15]
      state_15 <= AddRoundKeyModule_io_state_out_15;
    end else begin
      state_15 <= 8'h0;
    end
    if (reset) begin // @[Cipher.scala 32:23]
      rounds <= 4'h0; // @[Cipher.scala 32:23]
    end else if (2'h0 == STM) begin // @[Cipher.scala 38:15]
      rounds <= 4'h0; // @[Cipher.scala 43:14]
    end else if (2'h1 == STM) begin // @[Cipher.scala 38:15]
      rounds <= _rounds_T_1; // @[Cipher.scala 46:14]
    end else if (2'h2 == STM) begin // @[Cipher.scala 38:15]
      rounds <= _rounds_T_1; // @[Cipher.scala 50:14]
    end
    if (reset) begin // @[Cipher.scala 36:20]
      STM <= 2'h0; // @[Cipher.scala 36:20]
    end else if (2'h0 == STM) begin // @[Cipher.scala 38:15]
      if (io_start) begin // @[Cipher.scala 40:22]
        STM <= 2'h1; // @[Cipher.scala 41:13]
      end
    end else if (2'h1 == STM) begin // @[Cipher.scala 38:15]
      STM <= 2'h2; // @[Cipher.scala 47:11]
    end else if (2'h2 == STM) begin // @[Cipher.scala 38:15]
      STM <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  rounds = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  STM = _RAND_17[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AESEncrypt256(
  input          clock,
  input          reset,
  input          io_input_valid,
  input  [127:0] io_input_op1,
  input  [127:0] io_input_op2,
  output [255:0] io_output_text,
  output         io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  cipher_A_clock; // @[AESEncrypt.scala 95:26]
  wire  cipher_A_reset; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_0; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_1; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_2; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_3; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_4; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_5; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_6; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_7; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_8; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_9; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_10; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_11; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_12; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_13; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_14; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_plaintext_15; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_0; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_1; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_2; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_3; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_4; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_5; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_6; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_7; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_8; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_9; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_10; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_11; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_12; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_13; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_14; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_roundKey_15; // @[AESEncrypt.scala 95:26]
  wire  cipher_A_io_start; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_0; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_1; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_2; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_3; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_4; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_5; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_6; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_7; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_8; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_9; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_10; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_11; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_12; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_13; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_14; // @[AESEncrypt.scala 95:26]
  wire [7:0] cipher_A_io_state_out_15; // @[AESEncrypt.scala 95:26]
  wire  cipher_A_io_state_out_valid; // @[AESEncrypt.scala 95:26]
  wire  cipher_B_clock; // @[AESEncrypt.scala 96:26]
  wire  cipher_B_reset; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_0; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_1; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_2; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_3; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_4; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_5; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_6; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_7; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_8; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_9; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_10; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_11; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_12; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_13; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_14; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_plaintext_15; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_0; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_1; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_2; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_3; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_4; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_5; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_6; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_7; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_8; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_9; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_10; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_11; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_12; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_13; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_14; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_roundKey_15; // @[AESEncrypt.scala 96:26]
  wire  cipher_B_io_start; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_0; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_1; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_2; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_3; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_4; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_5; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_6; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_7; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_8; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_9; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_10; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_11; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_12; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_13; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_14; // @[AESEncrypt.scala 96:26]
  wire [7:0] cipher_B_io_state_out_15; // @[AESEncrypt.scala 96:26]
  wire  cipher_B_io_state_out_valid; // @[AESEncrypt.scala 96:26]
  reg [3:0] address; // @[AESEncrypt.scala 86:26]
  reg  tmp; // @[AESEncrypt.scala 88:22]
  wire [3:0] _address_T_1 = address + 4'h1; // @[AESEncrypt.scala 93:26]
  wire  _GEN_2 = io_input_valid & ~tmp | tmp; // @[AESEncrypt.scala 89:34 91:15 88:22]
  wire [7:0] _GEN_4 = 4'h1 == address ? 8'hd6 : 8'h0; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_5 = 4'h2 == address ? 8'hb6 : _GEN_4; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_6 = 4'h3 == address ? 8'hb6 : _GEN_5; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_7 = 4'h4 == address ? 8'h47 : _GEN_6; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_8 = 4'h5 == address ? 8'h3c : _GEN_7; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_9 = 4'h6 == address ? 8'h5e : _GEN_8; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_10 = 4'h7 == address ? 8'h14 : _GEN_9; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_11 = 4'h8 == address ? 8'h47 : _GEN_10; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_12 = 4'h9 == address ? 8'h54 : _GEN_11; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_15 = 4'h1 == address ? 8'haa : 8'h1; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_16 = 4'h2 == address ? 8'h92 : _GEN_15; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_17 = 4'h3 == address ? 8'hff : _GEN_16; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_18 = 4'h4 == address ? 8'hf7 : _GEN_17; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_19 = 4'h5 == address ? 8'haa : _GEN_18; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_20 = 4'h6 == address ? 8'h39 : _GEN_19; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_21 = 4'h7 == address ? 8'hf9 : _GEN_20; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_22 = 4'h8 == address ? 8'h43 : _GEN_21; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_23 = 4'h9 == address ? 8'h99 : _GEN_22; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_26 = 4'h1 == address ? 8'h74 : 8'h2; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_27 = 4'h2 == address ? 8'hcf : _GEN_26; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_28 = 4'h3 == address ? 8'h74 : _GEN_27; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_29 = 4'h4 == address ? 8'hf7 : _GEN_28; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_30 = 4'h5 == address ? 8'ha3 : _GEN_29; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_31 = 4'h6 == address ? 8'hf : _GEN_30; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_32 = 4'h7 == address ? 8'h70 : _GEN_31; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_33 = 4'h8 == address ? 8'h87 : _GEN_32; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_34 = 4'h9 == address ? 8'h32 : _GEN_33; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_37 = 4'h1 == address ? 8'hfd : 8'h3; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_38 = 4'h2 == address ? 8'hb : _GEN_37; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_39 = 4'h3 == address ? 8'h4e : _GEN_38; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_40 = 4'h4 == address ? 8'hbc : _GEN_39; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_41 = 4'h5 == address ? 8'he8 : _GEN_40; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_42 = 4'h6 == address ? 8'h7d : _GEN_41; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_43 = 4'h7 == address ? 8'h1a : _GEN_42; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_44 = 4'h8 == address ? 8'h35 : _GEN_43; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_45 = 4'h9 == address ? 8'hd1 : _GEN_44; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_48 = 4'h1 == address ? 8'hd2 : 8'h4; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_49 = 4'h2 == address ? 8'h64 : _GEN_48; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_50 = 4'h3 == address ? 8'hd2 : _GEN_49; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_51 = 4'h4 == address ? 8'h95 : _GEN_50; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_52 = 4'h5 == address ? 8'ha9 : _GEN_51; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_53 = 4'h6 == address ? 8'hf7 : _GEN_52; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_54 = 4'h7 == address ? 8'he3 : _GEN_53; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_55 = 4'h8 == address ? 8'ha4 : _GEN_54; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_56 = 4'h9 == address ? 8'hf0 : _GEN_55; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_59 = 4'h1 == address ? 8'haf : 8'h5; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_60 = 4'h2 == address ? 8'h3d : _GEN_59; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_61 = 4'h3 == address ? 8'hc2 : _GEN_60; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_62 = 4'h4 == address ? 8'h35 : _GEN_61; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_63 = 4'h5 == address ? 8'h9f : _GEN_62; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_64 = 4'h6 == address ? 8'ha6 : _GEN_63; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_65 = 4'h7 == address ? 8'h5f : _GEN_64; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_66 = 4'h8 == address ? 8'h1c : _GEN_65; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_67 = 4'h9 == address ? 8'h85 : _GEN_66; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_70 = 4'h1 == address ? 8'h72 : 8'h6; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_71 = 4'h2 == address ? 8'hbd : _GEN_70; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_72 = 4'h3 == address ? 8'hc9 : _GEN_71; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_73 = 4'h4 == address ? 8'h3e : _GEN_72; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_74 = 4'h5 == address ? 8'h9d : _GEN_73; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_75 = 4'h6 == address ? 8'h92 : _GEN_74; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_76 = 4'h7 == address ? 8'he2 : _GEN_75; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_77 = 4'h8 == address ? 8'h65 : _GEN_76; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_78 = 4'h9 == address ? 8'h57 : _GEN_77; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_81 = 4'h1 == address ? 8'hfa : 8'h7; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_82 = 4'h2 == address ? 8'hf1 : _GEN_81; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_83 = 4'h3 == address ? 8'hbf : _GEN_82; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_84 = 4'h4 == address ? 8'h3 : _GEN_83; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_85 = 4'h5 == address ? 8'heb : _GEN_84; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_86 = 4'h6 == address ? 8'h96 : _GEN_85; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_87 = 4'h7 == address ? 8'h8c : _GEN_86; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_88 = 4'h8 == address ? 8'hb9 : _GEN_87; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_89 = 4'h9 == address ? 8'h68 : _GEN_88; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_92 = 4'h1 == address ? 8'hda : 8'h8; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_93 = 4'h2 == address ? 8'hbe : _GEN_92; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_94 = 4'h3 == address ? 8'h6c : _GEN_93; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_95 = 4'h4 == address ? 8'hf9 : _GEN_94; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_96 = 4'h5 == address ? 8'h50 : _GEN_95; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_97 = 4'h6 == address ? 8'ha7 : _GEN_96; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_98 = 4'h7 == address ? 8'h44 : _GEN_97; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_99 = 4'h8 == address ? 8'he0 : _GEN_98; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_100 = 4'h9 == address ? 8'h10 : _GEN_99; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_103 = 4'h1 == address ? 8'ha6 : 8'h9; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_104 = 4'h2 == address ? 8'h9b : _GEN_103; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_105 = 4'h3 == address ? 8'h59 : _GEN_104; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_106 = 4'h4 == address ? 8'h6c : _GEN_105; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_107 = 4'h5 == address ? 8'hf3 : _GEN_106; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_108 = 4'h6 == address ? 8'h55 : _GEN_107; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_109 = 4'h7 == address ? 8'ha : _GEN_108; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_110 = 4'h8 == address ? 8'h16 : _GEN_109; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_111 = 4'h9 == address ? 8'h93 : _GEN_110; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_114 = 4'h1 == address ? 8'h78 : 8'ha; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_115 = 4'h2 == address ? 8'hc5 : _GEN_114; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_116 = 4'h3 == address ? 8'hc : _GEN_115; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_117 = 4'h4 == address ? 8'h32 : _GEN_116; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_118 = 4'h5 == address ? 8'haf : _GEN_117; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_119 = 4'h6 == address ? 8'h3d : _GEN_118; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_120 = 4'h7 == address ? 8'hdf : _GEN_119; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_121 = 4'h8 == address ? 8'hba : _GEN_120; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_122 = 4'h9 == address ? 8'hed : _GEN_121; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_125 = 4'h1 == address ? 8'hf1 : 8'hb; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_126 = 4'h2 == address ? 8'h0 : _GEN_125; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_127 = 4'h3 == address ? 8'hbf : _GEN_126; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_128 = 4'h4 == address ? 8'hbc : _GEN_127; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_129 = 4'h5 == address ? 8'h57 : _GEN_128; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_130 = 4'h6 == address ? 8'hc1 : _GEN_129; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_131 = 4'h7 == address ? 8'h4d : _GEN_130; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_132 = 4'h8 == address ? 8'hf4 : _GEN_131; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_133 = 4'h9 == address ? 8'h9c : _GEN_132; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_136 = 4'h1 == address ? 8'hd6 : 8'hc; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_137 = 4'h2 == address ? 8'h68 : _GEN_136; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_138 = 4'h3 == address ? 8'h4 : _GEN_137; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_139 = 4'h4 == address ? 8'hfd : _GEN_138; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_140 = 4'h5 == address ? 8'had : _GEN_139; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_141 = 4'h6 == address ? 8'ha : _GEN_140; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_142 = 4'h7 == address ? 8'h4e : _GEN_141; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_143 = 4'h8 == address ? 8'hae : _GEN_142; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_144 = 4'h9 == address ? 8'hbe : _GEN_143; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_147 = 4'h1 == address ? 8'hab : 8'hd; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_148 = 4'h2 == address ? 8'h30 : _GEN_147; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_149 = 4'h3 == address ? 8'h69 : _GEN_148; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_150 = 4'h4 == address ? 8'h5 : _GEN_149; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_151 = 4'h5 == address ? 8'hf6 : _GEN_150; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_152 = 4'h6 == address ? 8'ha3 : _GEN_151; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_153 = 4'h7 == address ? 8'ha9 : _GEN_152; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_154 = 4'h8 == address ? 8'hbf : _GEN_153; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_155 = 4'h9 == address ? 8'h2c : _GEN_154; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_158 = 4'h1 == address ? 8'h76 : 8'he; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_159 = 4'h2 == address ? 8'hb3 : _GEN_158; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_160 = 4'h3 == address ? 8'hbf : _GEN_159; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_161 = 4'h4 == address ? 8'h8d : _GEN_160; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_162 = 4'h5 == address ? 8'h22 : _GEN_161; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_163 = 4'h6 == address ? 8'h1f : _GEN_162; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_164 = 4'h7 == address ? 8'hc0 : _GEN_163; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_165 = 4'h8 == address ? 8'h7a : _GEN_164; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_166 = 4'h9 == address ? 8'h97 : _GEN_165; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_169 = 4'h1 == address ? 8'hfe : 8'hf; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_170 = 4'h2 == address ? 8'hfe : _GEN_169; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_171 = 4'h3 == address ? 8'h41 : _GEN_170; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_172 = 4'h4 == address ? 8'hfd : _GEN_171; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_173 = 4'h5 == address ? 8'haa : _GEN_172; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_174 = 4'h6 == address ? 8'h6b : _GEN_173; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_175 = 4'h7 == address ? 8'h26 : _GEN_174; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_176 = 4'h8 == address ? 8'hd2 : _GEN_175; // @[AESEncrypt.scala 102:{26,26}]
  wire [7:0] _GEN_177 = 4'h9 == address ? 8'h4e : _GEN_176; // @[AESEncrypt.scala 102:{26,26}]
  wire [63:0] io_output_text_lo = {cipher_B_io_state_out_8,cipher_B_io_state_out_9,cipher_B_io_state_out_10,
    cipher_B_io_state_out_11,cipher_B_io_state_out_12,cipher_B_io_state_out_13,cipher_B_io_state_out_14,
    cipher_B_io_state_out_15}; // @[Cat.scala 31:58]
  wire [127:0] _io_output_text_T = {cipher_B_io_state_out_0,cipher_B_io_state_out_1,cipher_B_io_state_out_2,
    cipher_B_io_state_out_3,cipher_B_io_state_out_4,cipher_B_io_state_out_5,cipher_B_io_state_out_6,
    cipher_B_io_state_out_7,io_output_text_lo}; // @[Cat.scala 31:58]
  wire [63:0] io_output_text_lo_1 = {cipher_A_io_state_out_8,cipher_A_io_state_out_9,cipher_A_io_state_out_10,
    cipher_A_io_state_out_11,cipher_A_io_state_out_12,cipher_A_io_state_out_13,cipher_A_io_state_out_14,
    cipher_A_io_state_out_15}; // @[Cat.scala 31:58]
  wire [127:0] _io_output_text_T_1 = {cipher_A_io_state_out_0,cipher_A_io_state_out_1,cipher_A_io_state_out_2,
    cipher_A_io_state_out_3,cipher_A_io_state_out_4,cipher_A_io_state_out_5,cipher_A_io_state_out_6,
    cipher_A_io_state_out_7,io_output_text_lo_1}; // @[Cat.scala 31:58]
  Cipher cipher_A ( // @[AESEncrypt.scala 95:26]
    .clock(cipher_A_clock),
    .reset(cipher_A_reset),
    .io_plaintext_0(cipher_A_io_plaintext_0),
    .io_plaintext_1(cipher_A_io_plaintext_1),
    .io_plaintext_2(cipher_A_io_plaintext_2),
    .io_plaintext_3(cipher_A_io_plaintext_3),
    .io_plaintext_4(cipher_A_io_plaintext_4),
    .io_plaintext_5(cipher_A_io_plaintext_5),
    .io_plaintext_6(cipher_A_io_plaintext_6),
    .io_plaintext_7(cipher_A_io_plaintext_7),
    .io_plaintext_8(cipher_A_io_plaintext_8),
    .io_plaintext_9(cipher_A_io_plaintext_9),
    .io_plaintext_10(cipher_A_io_plaintext_10),
    .io_plaintext_11(cipher_A_io_plaintext_11),
    .io_plaintext_12(cipher_A_io_plaintext_12),
    .io_plaintext_13(cipher_A_io_plaintext_13),
    .io_plaintext_14(cipher_A_io_plaintext_14),
    .io_plaintext_15(cipher_A_io_plaintext_15),
    .io_roundKey_0(cipher_A_io_roundKey_0),
    .io_roundKey_1(cipher_A_io_roundKey_1),
    .io_roundKey_2(cipher_A_io_roundKey_2),
    .io_roundKey_3(cipher_A_io_roundKey_3),
    .io_roundKey_4(cipher_A_io_roundKey_4),
    .io_roundKey_5(cipher_A_io_roundKey_5),
    .io_roundKey_6(cipher_A_io_roundKey_6),
    .io_roundKey_7(cipher_A_io_roundKey_7),
    .io_roundKey_8(cipher_A_io_roundKey_8),
    .io_roundKey_9(cipher_A_io_roundKey_9),
    .io_roundKey_10(cipher_A_io_roundKey_10),
    .io_roundKey_11(cipher_A_io_roundKey_11),
    .io_roundKey_12(cipher_A_io_roundKey_12),
    .io_roundKey_13(cipher_A_io_roundKey_13),
    .io_roundKey_14(cipher_A_io_roundKey_14),
    .io_roundKey_15(cipher_A_io_roundKey_15),
    .io_start(cipher_A_io_start),
    .io_state_out_0(cipher_A_io_state_out_0),
    .io_state_out_1(cipher_A_io_state_out_1),
    .io_state_out_2(cipher_A_io_state_out_2),
    .io_state_out_3(cipher_A_io_state_out_3),
    .io_state_out_4(cipher_A_io_state_out_4),
    .io_state_out_5(cipher_A_io_state_out_5),
    .io_state_out_6(cipher_A_io_state_out_6),
    .io_state_out_7(cipher_A_io_state_out_7),
    .io_state_out_8(cipher_A_io_state_out_8),
    .io_state_out_9(cipher_A_io_state_out_9),
    .io_state_out_10(cipher_A_io_state_out_10),
    .io_state_out_11(cipher_A_io_state_out_11),
    .io_state_out_12(cipher_A_io_state_out_12),
    .io_state_out_13(cipher_A_io_state_out_13),
    .io_state_out_14(cipher_A_io_state_out_14),
    .io_state_out_15(cipher_A_io_state_out_15),
    .io_state_out_valid(cipher_A_io_state_out_valid)
  );
  Cipher cipher_B ( // @[AESEncrypt.scala 96:26]
    .clock(cipher_B_clock),
    .reset(cipher_B_reset),
    .io_plaintext_0(cipher_B_io_plaintext_0),
    .io_plaintext_1(cipher_B_io_plaintext_1),
    .io_plaintext_2(cipher_B_io_plaintext_2),
    .io_plaintext_3(cipher_B_io_plaintext_3),
    .io_plaintext_4(cipher_B_io_plaintext_4),
    .io_plaintext_5(cipher_B_io_plaintext_5),
    .io_plaintext_6(cipher_B_io_plaintext_6),
    .io_plaintext_7(cipher_B_io_plaintext_7),
    .io_plaintext_8(cipher_B_io_plaintext_8),
    .io_plaintext_9(cipher_B_io_plaintext_9),
    .io_plaintext_10(cipher_B_io_plaintext_10),
    .io_plaintext_11(cipher_B_io_plaintext_11),
    .io_plaintext_12(cipher_B_io_plaintext_12),
    .io_plaintext_13(cipher_B_io_plaintext_13),
    .io_plaintext_14(cipher_B_io_plaintext_14),
    .io_plaintext_15(cipher_B_io_plaintext_15),
    .io_roundKey_0(cipher_B_io_roundKey_0),
    .io_roundKey_1(cipher_B_io_roundKey_1),
    .io_roundKey_2(cipher_B_io_roundKey_2),
    .io_roundKey_3(cipher_B_io_roundKey_3),
    .io_roundKey_4(cipher_B_io_roundKey_4),
    .io_roundKey_5(cipher_B_io_roundKey_5),
    .io_roundKey_6(cipher_B_io_roundKey_6),
    .io_roundKey_7(cipher_B_io_roundKey_7),
    .io_roundKey_8(cipher_B_io_roundKey_8),
    .io_roundKey_9(cipher_B_io_roundKey_9),
    .io_roundKey_10(cipher_B_io_roundKey_10),
    .io_roundKey_11(cipher_B_io_roundKey_11),
    .io_roundKey_12(cipher_B_io_roundKey_12),
    .io_roundKey_13(cipher_B_io_roundKey_13),
    .io_roundKey_14(cipher_B_io_roundKey_14),
    .io_roundKey_15(cipher_B_io_roundKey_15),
    .io_start(cipher_B_io_start),
    .io_state_out_0(cipher_B_io_state_out_0),
    .io_state_out_1(cipher_B_io_state_out_1),
    .io_state_out_2(cipher_B_io_state_out_2),
    .io_state_out_3(cipher_B_io_state_out_3),
    .io_state_out_4(cipher_B_io_state_out_4),
    .io_state_out_5(cipher_B_io_state_out_5),
    .io_state_out_6(cipher_B_io_state_out_6),
    .io_state_out_7(cipher_B_io_state_out_7),
    .io_state_out_8(cipher_B_io_state_out_8),
    .io_state_out_9(cipher_B_io_state_out_9),
    .io_state_out_10(cipher_B_io_state_out_10),
    .io_state_out_11(cipher_B_io_state_out_11),
    .io_state_out_12(cipher_B_io_state_out_12),
    .io_state_out_13(cipher_B_io_state_out_13),
    .io_state_out_14(cipher_B_io_state_out_14),
    .io_state_out_15(cipher_B_io_state_out_15),
    .io_state_out_valid(cipher_B_io_state_out_valid)
  );
  assign io_output_text = {_io_output_text_T,_io_output_text_T_1}; // @[Cat.scala 31:58]
  assign io_output_valid = cipher_A_io_state_out_valid & cipher_B_io_state_out_valid; // @[AESEncrypt.scala 107:52]
  assign cipher_A_clock = clock;
  assign cipher_A_reset = reset;
  assign cipher_A_io_plaintext_0 = io_input_op1[127:120]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_1 = io_input_op1[119:112]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_2 = io_input_op1[111:104]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_3 = io_input_op1[103:96]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_4 = io_input_op1[95:88]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_5 = io_input_op1[87:80]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_6 = io_input_op1[79:72]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_7 = io_input_op1[71:64]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_8 = io_input_op1[63:56]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_9 = io_input_op1[55:48]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_10 = io_input_op1[47:40]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_11 = io_input_op1[39:32]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_12 = io_input_op1[31:24]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_13 = io_input_op1[23:16]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_14 = io_input_op1[15:8]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_plaintext_15 = io_input_op1[7:0]; // @[AESEncrypt.scala 30:39]
  assign cipher_A_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_A_io_start = io_input_valid; // @[AESEncrypt.scala 98:23]
  assign cipher_B_clock = clock;
  assign cipher_B_reset = reset;
  assign cipher_B_io_plaintext_0 = io_input_op2[127:120]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_1 = io_input_op2[119:112]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_2 = io_input_op2[111:104]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_3 = io_input_op2[103:96]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_4 = io_input_op2[95:88]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_5 = io_input_op2[87:80]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_6 = io_input_op2[79:72]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_7 = io_input_op2[71:64]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_8 = io_input_op2[63:56]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_9 = io_input_op2[55:48]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_10 = io_input_op2[47:40]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_11 = io_input_op2[39:32]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_12 = io_input_op2[31:24]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_13 = io_input_op2[23:16]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_14 = io_input_op2[15:8]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_plaintext_15 = io_input_op2[7:0]; // @[AESEncrypt.scala 31:39]
  assign cipher_B_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESEncrypt.scala 102:{26,26}]
  assign cipher_B_io_start = io_input_valid; // @[AESEncrypt.scala 99:23]
  always @(posedge clock) begin
    if (reset) begin // @[AESEncrypt.scala 86:26]
      address <= 4'h0; // @[AESEncrypt.scala 86:26]
    end else if (io_input_valid & ~tmp) begin // @[AESEncrypt.scala 89:34]
      address <= 4'h0; // @[AESEncrypt.scala 90:15]
    end else if (address != 4'ha) begin // @[AESEncrypt.scala 92:33]
      address <= _address_T_1; // @[AESEncrypt.scala 93:15]
    end
    if (reset) begin // @[AESEncrypt.scala 88:22]
      tmp <= 1'h0; // @[AESEncrypt.scala 88:22]
    end else begin
      tmp <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  address = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  tmp = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AESEncrypt(
  input          clock,
  input          reset,
  input          io_input_valid,
  input  [127:0] io_input_text,
  output [127:0] io_output_text,
  output         io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  cipher_clock; // @[AESEncrypt.scala 176:24]
  wire  cipher_reset; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_0; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_1; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_2; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_3; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_4; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_5; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_6; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_7; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_8; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_9; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_10; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_11; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_12; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_13; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_14; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_plaintext_15; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_0; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_1; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_2; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_3; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_4; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_5; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_6; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_7; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_8; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_9; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_10; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_11; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_12; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_13; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_14; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_roundKey_15; // @[AESEncrypt.scala 176:24]
  wire  cipher_io_start; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_0; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_1; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_2; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_3; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_4; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_5; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_6; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_7; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_8; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_9; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_10; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_11; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_12; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_13; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_14; // @[AESEncrypt.scala 176:24]
  wire [7:0] cipher_io_state_out_15; // @[AESEncrypt.scala 176:24]
  wire  cipher_io_state_out_valid; // @[AESEncrypt.scala 176:24]
  reg [3:0] address; // @[AESEncrypt.scala 167:26]
  reg  tmp; // @[AESEncrypt.scala 169:22]
  wire [3:0] _address_T_1 = address + 4'h1; // @[AESEncrypt.scala 174:26]
  wire  _GEN_2 = io_input_valid & ~tmp | tmp; // @[AESEncrypt.scala 170:34 172:15 169:22]
  wire [7:0] _GEN_4 = 4'h1 == address ? 8'hd6 : 8'h0; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_5 = 4'h2 == address ? 8'hb6 : _GEN_4; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_6 = 4'h3 == address ? 8'hb6 : _GEN_5; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_7 = 4'h4 == address ? 8'h47 : _GEN_6; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_8 = 4'h5 == address ? 8'h3c : _GEN_7; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_9 = 4'h6 == address ? 8'h5e : _GEN_8; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_10 = 4'h7 == address ? 8'h14 : _GEN_9; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_11 = 4'h8 == address ? 8'h47 : _GEN_10; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_12 = 4'h9 == address ? 8'h54 : _GEN_11; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_15 = 4'h1 == address ? 8'haa : 8'h1; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_16 = 4'h2 == address ? 8'h92 : _GEN_15; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_17 = 4'h3 == address ? 8'hff : _GEN_16; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_18 = 4'h4 == address ? 8'hf7 : _GEN_17; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_19 = 4'h5 == address ? 8'haa : _GEN_18; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_20 = 4'h6 == address ? 8'h39 : _GEN_19; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_21 = 4'h7 == address ? 8'hf9 : _GEN_20; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_22 = 4'h8 == address ? 8'h43 : _GEN_21; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_23 = 4'h9 == address ? 8'h99 : _GEN_22; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_26 = 4'h1 == address ? 8'h74 : 8'h2; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_27 = 4'h2 == address ? 8'hcf : _GEN_26; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_28 = 4'h3 == address ? 8'h74 : _GEN_27; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_29 = 4'h4 == address ? 8'hf7 : _GEN_28; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_30 = 4'h5 == address ? 8'ha3 : _GEN_29; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_31 = 4'h6 == address ? 8'hf : _GEN_30; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_32 = 4'h7 == address ? 8'h70 : _GEN_31; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_33 = 4'h8 == address ? 8'h87 : _GEN_32; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_34 = 4'h9 == address ? 8'h32 : _GEN_33; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_37 = 4'h1 == address ? 8'hfd : 8'h3; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_38 = 4'h2 == address ? 8'hb : _GEN_37; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_39 = 4'h3 == address ? 8'h4e : _GEN_38; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_40 = 4'h4 == address ? 8'hbc : _GEN_39; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_41 = 4'h5 == address ? 8'he8 : _GEN_40; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_42 = 4'h6 == address ? 8'h7d : _GEN_41; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_43 = 4'h7 == address ? 8'h1a : _GEN_42; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_44 = 4'h8 == address ? 8'h35 : _GEN_43; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_45 = 4'h9 == address ? 8'hd1 : _GEN_44; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_48 = 4'h1 == address ? 8'hd2 : 8'h4; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_49 = 4'h2 == address ? 8'h64 : _GEN_48; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_50 = 4'h3 == address ? 8'hd2 : _GEN_49; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_51 = 4'h4 == address ? 8'h95 : _GEN_50; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_52 = 4'h5 == address ? 8'ha9 : _GEN_51; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_53 = 4'h6 == address ? 8'hf7 : _GEN_52; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_54 = 4'h7 == address ? 8'he3 : _GEN_53; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_55 = 4'h8 == address ? 8'ha4 : _GEN_54; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_56 = 4'h9 == address ? 8'hf0 : _GEN_55; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_59 = 4'h1 == address ? 8'haf : 8'h5; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_60 = 4'h2 == address ? 8'h3d : _GEN_59; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_61 = 4'h3 == address ? 8'hc2 : _GEN_60; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_62 = 4'h4 == address ? 8'h35 : _GEN_61; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_63 = 4'h5 == address ? 8'h9f : _GEN_62; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_64 = 4'h6 == address ? 8'ha6 : _GEN_63; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_65 = 4'h7 == address ? 8'h5f : _GEN_64; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_66 = 4'h8 == address ? 8'h1c : _GEN_65; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_67 = 4'h9 == address ? 8'h85 : _GEN_66; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_70 = 4'h1 == address ? 8'h72 : 8'h6; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_71 = 4'h2 == address ? 8'hbd : _GEN_70; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_72 = 4'h3 == address ? 8'hc9 : _GEN_71; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_73 = 4'h4 == address ? 8'h3e : _GEN_72; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_74 = 4'h5 == address ? 8'h9d : _GEN_73; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_75 = 4'h6 == address ? 8'h92 : _GEN_74; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_76 = 4'h7 == address ? 8'he2 : _GEN_75; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_77 = 4'h8 == address ? 8'h65 : _GEN_76; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_78 = 4'h9 == address ? 8'h57 : _GEN_77; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_81 = 4'h1 == address ? 8'hfa : 8'h7; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_82 = 4'h2 == address ? 8'hf1 : _GEN_81; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_83 = 4'h3 == address ? 8'hbf : _GEN_82; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_84 = 4'h4 == address ? 8'h3 : _GEN_83; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_85 = 4'h5 == address ? 8'heb : _GEN_84; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_86 = 4'h6 == address ? 8'h96 : _GEN_85; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_87 = 4'h7 == address ? 8'h8c : _GEN_86; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_88 = 4'h8 == address ? 8'hb9 : _GEN_87; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_89 = 4'h9 == address ? 8'h68 : _GEN_88; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_92 = 4'h1 == address ? 8'hda : 8'h8; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_93 = 4'h2 == address ? 8'hbe : _GEN_92; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_94 = 4'h3 == address ? 8'h6c : _GEN_93; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_95 = 4'h4 == address ? 8'hf9 : _GEN_94; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_96 = 4'h5 == address ? 8'h50 : _GEN_95; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_97 = 4'h6 == address ? 8'ha7 : _GEN_96; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_98 = 4'h7 == address ? 8'h44 : _GEN_97; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_99 = 4'h8 == address ? 8'he0 : _GEN_98; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_100 = 4'h9 == address ? 8'h10 : _GEN_99; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_103 = 4'h1 == address ? 8'ha6 : 8'h9; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_104 = 4'h2 == address ? 8'h9b : _GEN_103; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_105 = 4'h3 == address ? 8'h59 : _GEN_104; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_106 = 4'h4 == address ? 8'h6c : _GEN_105; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_107 = 4'h5 == address ? 8'hf3 : _GEN_106; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_108 = 4'h6 == address ? 8'h55 : _GEN_107; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_109 = 4'h7 == address ? 8'ha : _GEN_108; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_110 = 4'h8 == address ? 8'h16 : _GEN_109; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_111 = 4'h9 == address ? 8'h93 : _GEN_110; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_114 = 4'h1 == address ? 8'h78 : 8'ha; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_115 = 4'h2 == address ? 8'hc5 : _GEN_114; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_116 = 4'h3 == address ? 8'hc : _GEN_115; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_117 = 4'h4 == address ? 8'h32 : _GEN_116; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_118 = 4'h5 == address ? 8'haf : _GEN_117; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_119 = 4'h6 == address ? 8'h3d : _GEN_118; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_120 = 4'h7 == address ? 8'hdf : _GEN_119; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_121 = 4'h8 == address ? 8'hba : _GEN_120; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_122 = 4'h9 == address ? 8'hed : _GEN_121; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_125 = 4'h1 == address ? 8'hf1 : 8'hb; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_126 = 4'h2 == address ? 8'h0 : _GEN_125; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_127 = 4'h3 == address ? 8'hbf : _GEN_126; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_128 = 4'h4 == address ? 8'hbc : _GEN_127; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_129 = 4'h5 == address ? 8'h57 : _GEN_128; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_130 = 4'h6 == address ? 8'hc1 : _GEN_129; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_131 = 4'h7 == address ? 8'h4d : _GEN_130; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_132 = 4'h8 == address ? 8'hf4 : _GEN_131; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_133 = 4'h9 == address ? 8'h9c : _GEN_132; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_136 = 4'h1 == address ? 8'hd6 : 8'hc; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_137 = 4'h2 == address ? 8'h68 : _GEN_136; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_138 = 4'h3 == address ? 8'h4 : _GEN_137; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_139 = 4'h4 == address ? 8'hfd : _GEN_138; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_140 = 4'h5 == address ? 8'had : _GEN_139; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_141 = 4'h6 == address ? 8'ha : _GEN_140; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_142 = 4'h7 == address ? 8'h4e : _GEN_141; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_143 = 4'h8 == address ? 8'hae : _GEN_142; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_144 = 4'h9 == address ? 8'hbe : _GEN_143; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_147 = 4'h1 == address ? 8'hab : 8'hd; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_148 = 4'h2 == address ? 8'h30 : _GEN_147; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_149 = 4'h3 == address ? 8'h69 : _GEN_148; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_150 = 4'h4 == address ? 8'h5 : _GEN_149; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_151 = 4'h5 == address ? 8'hf6 : _GEN_150; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_152 = 4'h6 == address ? 8'ha3 : _GEN_151; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_153 = 4'h7 == address ? 8'ha9 : _GEN_152; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_154 = 4'h8 == address ? 8'hbf : _GEN_153; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_155 = 4'h9 == address ? 8'h2c : _GEN_154; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_158 = 4'h1 == address ? 8'h76 : 8'he; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_159 = 4'h2 == address ? 8'hb3 : _GEN_158; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_160 = 4'h3 == address ? 8'hbf : _GEN_159; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_161 = 4'h4 == address ? 8'h8d : _GEN_160; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_162 = 4'h5 == address ? 8'h22 : _GEN_161; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_163 = 4'h6 == address ? 8'h1f : _GEN_162; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_164 = 4'h7 == address ? 8'hc0 : _GEN_163; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_165 = 4'h8 == address ? 8'h7a : _GEN_164; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_166 = 4'h9 == address ? 8'h97 : _GEN_165; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_169 = 4'h1 == address ? 8'hfe : 8'hf; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_170 = 4'h2 == address ? 8'hfe : _GEN_169; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_171 = 4'h3 == address ? 8'h41 : _GEN_170; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_172 = 4'h4 == address ? 8'hfd : _GEN_171; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_173 = 4'h5 == address ? 8'haa : _GEN_172; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_174 = 4'h6 == address ? 8'h6b : _GEN_173; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_175 = 4'h7 == address ? 8'h26 : _GEN_174; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_176 = 4'h8 == address ? 8'hd2 : _GEN_175; // @[AESEncrypt.scala 179:{24,24}]
  wire [7:0] _GEN_177 = 4'h9 == address ? 8'h4e : _GEN_176; // @[AESEncrypt.scala 179:{24,24}]
  wire [63:0] io_output_text_lo = {cipher_io_state_out_8,cipher_io_state_out_9,cipher_io_state_out_10,
    cipher_io_state_out_11,cipher_io_state_out_12,cipher_io_state_out_13,cipher_io_state_out_14,cipher_io_state_out_15}; // @[Cat.scala 31:58]
  wire [63:0] io_output_text_hi = {cipher_io_state_out_0,cipher_io_state_out_1,cipher_io_state_out_2,
    cipher_io_state_out_3,cipher_io_state_out_4,cipher_io_state_out_5,cipher_io_state_out_6,cipher_io_state_out_7}; // @[Cat.scala 31:58]
  Cipher cipher ( // @[AESEncrypt.scala 176:24]
    .clock(cipher_clock),
    .reset(cipher_reset),
    .io_plaintext_0(cipher_io_plaintext_0),
    .io_plaintext_1(cipher_io_plaintext_1),
    .io_plaintext_2(cipher_io_plaintext_2),
    .io_plaintext_3(cipher_io_plaintext_3),
    .io_plaintext_4(cipher_io_plaintext_4),
    .io_plaintext_5(cipher_io_plaintext_5),
    .io_plaintext_6(cipher_io_plaintext_6),
    .io_plaintext_7(cipher_io_plaintext_7),
    .io_plaintext_8(cipher_io_plaintext_8),
    .io_plaintext_9(cipher_io_plaintext_9),
    .io_plaintext_10(cipher_io_plaintext_10),
    .io_plaintext_11(cipher_io_plaintext_11),
    .io_plaintext_12(cipher_io_plaintext_12),
    .io_plaintext_13(cipher_io_plaintext_13),
    .io_plaintext_14(cipher_io_plaintext_14),
    .io_plaintext_15(cipher_io_plaintext_15),
    .io_roundKey_0(cipher_io_roundKey_0),
    .io_roundKey_1(cipher_io_roundKey_1),
    .io_roundKey_2(cipher_io_roundKey_2),
    .io_roundKey_3(cipher_io_roundKey_3),
    .io_roundKey_4(cipher_io_roundKey_4),
    .io_roundKey_5(cipher_io_roundKey_5),
    .io_roundKey_6(cipher_io_roundKey_6),
    .io_roundKey_7(cipher_io_roundKey_7),
    .io_roundKey_8(cipher_io_roundKey_8),
    .io_roundKey_9(cipher_io_roundKey_9),
    .io_roundKey_10(cipher_io_roundKey_10),
    .io_roundKey_11(cipher_io_roundKey_11),
    .io_roundKey_12(cipher_io_roundKey_12),
    .io_roundKey_13(cipher_io_roundKey_13),
    .io_roundKey_14(cipher_io_roundKey_14),
    .io_roundKey_15(cipher_io_roundKey_15),
    .io_start(cipher_io_start),
    .io_state_out_0(cipher_io_state_out_0),
    .io_state_out_1(cipher_io_state_out_1),
    .io_state_out_2(cipher_io_state_out_2),
    .io_state_out_3(cipher_io_state_out_3),
    .io_state_out_4(cipher_io_state_out_4),
    .io_state_out_5(cipher_io_state_out_5),
    .io_state_out_6(cipher_io_state_out_6),
    .io_state_out_7(cipher_io_state_out_7),
    .io_state_out_8(cipher_io_state_out_8),
    .io_state_out_9(cipher_io_state_out_9),
    .io_state_out_10(cipher_io_state_out_10),
    .io_state_out_11(cipher_io_state_out_11),
    .io_state_out_12(cipher_io_state_out_12),
    .io_state_out_13(cipher_io_state_out_13),
    .io_state_out_14(cipher_io_state_out_14),
    .io_state_out_15(cipher_io_state_out_15),
    .io_state_out_valid(cipher_io_state_out_valid)
  );
  assign io_output_text = {io_output_text_hi,io_output_text_lo}; // @[Cat.scala 31:58]
  assign io_output_valid = cipher_io_state_out_valid; // @[AESEncrypt.scala 183:21]
  assign cipher_clock = clock;
  assign cipher_reset = reset;
  assign cipher_io_plaintext_0 = io_input_text[127:120]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_1 = io_input_text[119:112]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_2 = io_input_text[111:104]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_3 = io_input_text[103:96]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_4 = io_input_text[95:88]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_5 = io_input_text[87:80]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_6 = io_input_text[79:72]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_7 = io_input_text[71:64]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_8 = io_input_text[63:56]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_9 = io_input_text[55:48]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_10 = io_input_text[47:40]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_11 = io_input_text[39:32]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_12 = io_input_text[31:24]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_13 = io_input_text[23:16]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_14 = io_input_text[15:8]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_plaintext_15 = io_input_text[7:0]; // @[AESEncrypt.scala 133:39]
  assign cipher_io_roundKey_0 = 4'ha == address ? 8'h13 : _GEN_12; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_1 = 4'ha == address ? 8'h11 : _GEN_23; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_2 = 4'ha == address ? 8'h1d : _GEN_34; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_3 = 4'ha == address ? 8'h7f : _GEN_45; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_4 = 4'ha == address ? 8'he3 : _GEN_56; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_5 = 4'ha == address ? 8'h94 : _GEN_67; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_6 = 4'ha == address ? 8'h4a : _GEN_78; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_7 = 4'ha == address ? 8'h17 : _GEN_89; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_8 = 4'ha == address ? 8'hf3 : _GEN_100; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_9 = 4'ha == address ? 8'h7 : _GEN_111; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_10 = 4'ha == address ? 8'ha7 : _GEN_122; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_11 = 4'ha == address ? 8'h8b : _GEN_133; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_12 = 4'ha == address ? 8'h4d : _GEN_144; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_13 = 4'ha == address ? 8'h2b : _GEN_155; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_14 = 4'ha == address ? 8'h30 : _GEN_166; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_roundKey_15 = 4'ha == address ? 8'hc5 : _GEN_177; // @[AESEncrypt.scala 179:{24,24}]
  assign cipher_io_start = io_input_valid; // @[AESEncrypt.scala 177:21]
  always @(posedge clock) begin
    if (reset) begin // @[AESEncrypt.scala 167:26]
      address <= 4'h0; // @[AESEncrypt.scala 167:26]
    end else if (io_input_valid & ~tmp) begin // @[AESEncrypt.scala 170:34]
      address <= 4'h0; // @[AESEncrypt.scala 171:15]
    end else if (address != 4'ha) begin // @[AESEncrypt.scala 173:33]
      address <= _address_T_1; // @[AESEncrypt.scala 174:15]
    end
    if (reset) begin // @[AESEncrypt.scala 169:22]
      tmp <= 1'h0; // @[AESEncrypt.scala 169:22]
    end else begin
      tmp <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  address = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  tmp = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Plaintext_Reverse_Connector(
  input  [315:0] io_op1,
  input  [315:0] io_op2,
  input  [7:0]   io_inst,
  output [7:0]   io_out_0,
  output [7:0]   io_out_1,
  output [7:0]   io_out_2,
  output [7:0]   io_out_3,
  output [7:0]   io_out_4,
  output [7:0]   io_out_5,
  output [7:0]   io_out_6,
  output [7:0]   io_out_7,
  output [7:0]   io_out_8,
  output [7:0]   io_out_9,
  output [7:0]   io_out_10,
  output [7:0]   io_out_11,
  output [7:0]   io_out_12,
  output [7:0]   io_out_13,
  output [7:0]   io_out_14,
  output [7:0]   io_out_15
);
  wire [59:0] op1_hash = io_op1[315:256]; // @[SE.scala 66:41]
  wire [59:0] op2_hash = io_op2[315:256]; // @[SE.scala 67:41]
  wire [127:0] connect_result = {op1_hash,op2_hash,io_inst}; // @[Cat.scala 31:58]
  assign io_out_0 = connect_result[7:0]; // @[SE.scala 74:60]
  assign io_out_1 = connect_result[15:8]; // @[SE.scala 74:60]
  assign io_out_2 = connect_result[23:16]; // @[SE.scala 74:60]
  assign io_out_3 = connect_result[31:24]; // @[SE.scala 74:60]
  assign io_out_4 = connect_result[39:32]; // @[SE.scala 74:60]
  assign io_out_5 = connect_result[47:40]; // @[SE.scala 74:60]
  assign io_out_6 = connect_result[55:48]; // @[SE.scala 74:60]
  assign io_out_7 = connect_result[63:56]; // @[SE.scala 74:60]
  assign io_out_8 = connect_result[71:64]; // @[SE.scala 74:60]
  assign io_out_9 = connect_result[79:72]; // @[SE.scala 74:60]
  assign io_out_10 = connect_result[87:80]; // @[SE.scala 74:60]
  assign io_out_11 = connect_result[95:88]; // @[SE.scala 74:60]
  assign io_out_12 = connect_result[103:96]; // @[SE.scala 74:60]
  assign io_out_13 = connect_result[111:104]; // @[SE.scala 74:60]
  assign io_out_14 = connect_result[119:112]; // @[SE.scala 74:60]
  assign io_out_15 = connect_result[127:120]; // @[SE.scala 74:60]
endmodule
module Hash_Compare(
  input  [59:0] io_hash_orig,
  input  [59:0] io_hash_regenerated,
  input         io_valid_in,
  output        io_valid_out,
  output        io_compare_result
);
  assign io_valid_out = io_valid_in; // @[SE.scala 96:47]
  assign io_compare_result = io_hash_orig == io_hash_regenerated; // @[SE.scala 97:49]
endmodule
module Version_ID_Generator(
  input         io_pub_priv_opA,
  input         io_pub_priv_opB,
  input  [15:0] io_version_id_opA,
  input  [15:0] io_version_id_opB,
  input         io_valid_in,
  output        io_valid_out,
  output [15:0] io_version_id_out,
  output        io_pub_priv_out
);
  wire  _T_1 = ~io_pub_priv_opB; // @[SE.scala 124:38]
  wire [15:0] _GEN_0 = io_version_id_opA != io_version_id_opB ? 16'hffff : io_version_id_opA; // @[SE.scala 126:71 127:47 129:47]
  wire [15:0] _GEN_1 = ~io_pub_priv_opB ? _GEN_0 : io_version_id_opA; // @[SE.scala 124:51 133:39]
  wire [15:0] _GEN_2 = _T_1 ? io_version_id_opB : 16'h0; // @[SE.scala 136:51 138:39 141:39]
  assign io_valid_out = io_valid_in; // @[SE.scala 121:39]
  assign io_version_id_out = ~io_pub_priv_opA ? _GEN_1 : _GEN_2; // @[SE.scala 123:43]
  assign io_pub_priv_out = io_pub_priv_opA & io_pub_priv_opB; // @[SE.scala 147:38]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  input   io_increment,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19,
  output  io_out_20,
  output  io_out_21,
  output  io_out_22,
  output  io_out_23,
  output  io_out_24,
  output  io_out_25,
  output  io_out_26,
  output  io_out_27,
  output  io_out_28,
  output  io_out_29,
  output  io_out_30,
  output  io_out_31,
  output  io_out_32,
  output  io_out_33,
  output  io_out_34,
  output  io_out_35,
  output  io_out_36,
  output  io_out_37,
  output  io_out_38,
  output  io_out_39,
  output  io_out_40,
  output  io_out_41,
  output  io_out_42,
  output  io_out_43,
  output  io_out_44,
  output  io_out_45,
  output  io_out_46,
  output  io_out_47,
  output  io_out_48,
  output  io_out_49,
  output  io_out_50,
  output  io_out_51,
  output  io_out_52,
  output  io_out_53,
  output  io_out_54,
  output  io_out_55,
  output  io_out_56,
  output  io_out_57,
  output  io_out_58,
  output  io_out_59,
  output  io_out_60,
  output  io_out_61,
  output  io_out_62,
  output  io_out_63
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  reg  state_16; // @[PRNG.scala 55:49]
  reg  state_17; // @[PRNG.scala 55:49]
  reg  state_18; // @[PRNG.scala 55:49]
  reg  state_19; // @[PRNG.scala 55:49]
  reg  state_20; // @[PRNG.scala 55:49]
  reg  state_21; // @[PRNG.scala 55:49]
  reg  state_22; // @[PRNG.scala 55:49]
  reg  state_23; // @[PRNG.scala 55:49]
  reg  state_24; // @[PRNG.scala 55:49]
  reg  state_25; // @[PRNG.scala 55:49]
  reg  state_26; // @[PRNG.scala 55:49]
  reg  state_27; // @[PRNG.scala 55:49]
  reg  state_28; // @[PRNG.scala 55:49]
  reg  state_29; // @[PRNG.scala 55:49]
  reg  state_30; // @[PRNG.scala 55:49]
  reg  state_31; // @[PRNG.scala 55:49]
  reg  state_32; // @[PRNG.scala 55:49]
  reg  state_33; // @[PRNG.scala 55:49]
  reg  state_34; // @[PRNG.scala 55:49]
  reg  state_35; // @[PRNG.scala 55:49]
  reg  state_36; // @[PRNG.scala 55:49]
  reg  state_37; // @[PRNG.scala 55:49]
  reg  state_38; // @[PRNG.scala 55:49]
  reg  state_39; // @[PRNG.scala 55:49]
  reg  state_40; // @[PRNG.scala 55:49]
  reg  state_41; // @[PRNG.scala 55:49]
  reg  state_42; // @[PRNG.scala 55:49]
  reg  state_43; // @[PRNG.scala 55:49]
  reg  state_44; // @[PRNG.scala 55:49]
  reg  state_45; // @[PRNG.scala 55:49]
  reg  state_46; // @[PRNG.scala 55:49]
  reg  state_47; // @[PRNG.scala 55:49]
  reg  state_48; // @[PRNG.scala 55:49]
  reg  state_49; // @[PRNG.scala 55:49]
  reg  state_50; // @[PRNG.scala 55:49]
  reg  state_51; // @[PRNG.scala 55:49]
  reg  state_52; // @[PRNG.scala 55:49]
  reg  state_53; // @[PRNG.scala 55:49]
  reg  state_54; // @[PRNG.scala 55:49]
  reg  state_55; // @[PRNG.scala 55:49]
  reg  state_56; // @[PRNG.scala 55:49]
  reg  state_57; // @[PRNG.scala 55:49]
  reg  state_58; // @[PRNG.scala 55:49]
  reg  state_59; // @[PRNG.scala 55:49]
  reg  state_60; // @[PRNG.scala 55:49]
  reg  state_61; // @[PRNG.scala 55:49]
  reg  state_62; // @[PRNG.scala 55:49]
  reg  state_63; // @[PRNG.scala 55:49]
  wire  _T_2 = state_63 ^ state_62 ^ state_60 ^ state_59; // @[LFSR.scala 15:41]
  wire  _GEN_0 = io_increment ? _T_2 : state_0; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_1 = io_increment ? state_0 : state_1; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_2 = io_increment ? state_1 : state_2; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_3 = io_increment ? state_2 : state_3; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_5 = io_increment ? state_4 : state_5; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_6 = io_increment ? state_5 : state_6; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_7 = io_increment ? state_6 : state_7; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_9 = io_increment ? state_8 : state_9; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_10 = io_increment ? state_9 : state_10; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_11 = io_increment ? state_10 : state_11; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_12 = io_increment ? state_11 : state_12; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_13 = io_increment ? state_12 : state_13; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_15 = io_increment ? state_14 : state_15; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_16 = io_increment ? state_15 : state_16; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_18 = io_increment ? state_17 : state_18; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_19 = io_increment ? state_18 : state_19; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_21 = io_increment ? state_20 : state_21; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_23 = io_increment ? state_22 : state_23; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_25 = io_increment ? state_24 : state_25; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_26 = io_increment ? state_25 : state_26; // @[PRNG.scala 69:22 70:11 55:49]
  wire  _GEN_27 = io_increment ? state_26 : state_27; // @[PRNG.scala 69:22 70:11 55:49]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  assign io_out_16 = state_16; // @[PRNG.scala 78:10]
  assign io_out_17 = state_17; // @[PRNG.scala 78:10]
  assign io_out_18 = state_18; // @[PRNG.scala 78:10]
  assign io_out_19 = state_19; // @[PRNG.scala 78:10]
  assign io_out_20 = state_20; // @[PRNG.scala 78:10]
  assign io_out_21 = state_21; // @[PRNG.scala 78:10]
  assign io_out_22 = state_22; // @[PRNG.scala 78:10]
  assign io_out_23 = state_23; // @[PRNG.scala 78:10]
  assign io_out_24 = state_24; // @[PRNG.scala 78:10]
  assign io_out_25 = state_25; // @[PRNG.scala 78:10]
  assign io_out_26 = state_26; // @[PRNG.scala 78:10]
  assign io_out_27 = state_27; // @[PRNG.scala 78:10]
  assign io_out_28 = state_28; // @[PRNG.scala 78:10]
  assign io_out_29 = state_29; // @[PRNG.scala 78:10]
  assign io_out_30 = state_30; // @[PRNG.scala 78:10]
  assign io_out_31 = state_31; // @[PRNG.scala 78:10]
  assign io_out_32 = state_32; // @[PRNG.scala 78:10]
  assign io_out_33 = state_33; // @[PRNG.scala 78:10]
  assign io_out_34 = state_34; // @[PRNG.scala 78:10]
  assign io_out_35 = state_35; // @[PRNG.scala 78:10]
  assign io_out_36 = state_36; // @[PRNG.scala 78:10]
  assign io_out_37 = state_37; // @[PRNG.scala 78:10]
  assign io_out_38 = state_38; // @[PRNG.scala 78:10]
  assign io_out_39 = state_39; // @[PRNG.scala 78:10]
  assign io_out_40 = state_40; // @[PRNG.scala 78:10]
  assign io_out_41 = state_41; // @[PRNG.scala 78:10]
  assign io_out_42 = state_42; // @[PRNG.scala 78:10]
  assign io_out_43 = state_43; // @[PRNG.scala 78:10]
  assign io_out_44 = state_44; // @[PRNG.scala 78:10]
  assign io_out_45 = state_45; // @[PRNG.scala 78:10]
  assign io_out_46 = state_46; // @[PRNG.scala 78:10]
  assign io_out_47 = state_47; // @[PRNG.scala 78:10]
  assign io_out_48 = state_48; // @[PRNG.scala 78:10]
  assign io_out_49 = state_49; // @[PRNG.scala 78:10]
  assign io_out_50 = state_50; // @[PRNG.scala 78:10]
  assign io_out_51 = state_51; // @[PRNG.scala 78:10]
  assign io_out_52 = state_52; // @[PRNG.scala 78:10]
  assign io_out_53 = state_53; // @[PRNG.scala 78:10]
  assign io_out_54 = state_54; // @[PRNG.scala 78:10]
  assign io_out_55 = state_55; // @[PRNG.scala 78:10]
  assign io_out_56 = state_56; // @[PRNG.scala 78:10]
  assign io_out_57 = state_57; // @[PRNG.scala 78:10]
  assign io_out_58 = state_58; // @[PRNG.scala 78:10]
  assign io_out_59 = state_59; // @[PRNG.scala 78:10]
  assign io_out_60 = state_60; // @[PRNG.scala 78:10]
  assign io_out_61 = state_61; // @[PRNG.scala 78:10]
  assign io_out_62 = state_62; // @[PRNG.scala 78:10]
  assign io_out_63 = state_63; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _GEN_0; // @[PRNG.scala 55:{49,49}]
    state_1 <= reset | _GEN_1; // @[PRNG.scala 55:{49,49}]
    state_2 <= reset | _GEN_2; // @[PRNG.scala 55:{49,49}]
    state_3 <= reset | _GEN_3; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_4 <= state_3; // @[PRNG.scala 70:11]
    end
    state_5 <= reset | _GEN_5; // @[PRNG.scala 55:{49,49}]
    state_6 <= reset | _GEN_6; // @[PRNG.scala 55:{49,49}]
    state_7 <= reset | _GEN_7; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_8 <= state_7; // @[PRNG.scala 70:11]
    end
    state_9 <= reset | _GEN_9; // @[PRNG.scala 55:{49,49}]
    state_10 <= reset | _GEN_10; // @[PRNG.scala 55:{49,49}]
    state_11 <= reset | _GEN_11; // @[PRNG.scala 55:{49,49}]
    state_12 <= reset | _GEN_12; // @[PRNG.scala 55:{49,49}]
    state_13 <= reset | _GEN_13; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_14 <= state_13; // @[PRNG.scala 70:11]
    end
    state_15 <= reset | _GEN_15; // @[PRNG.scala 55:{49,49}]
    state_16 <= reset | _GEN_16; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_17 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_17 <= state_16; // @[PRNG.scala 70:11]
    end
    state_18 <= reset | _GEN_18; // @[PRNG.scala 55:{49,49}]
    state_19 <= reset | _GEN_19; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_20 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_20 <= state_19; // @[PRNG.scala 70:11]
    end
    state_21 <= reset | _GEN_21; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_22 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_22 <= state_21; // @[PRNG.scala 70:11]
    end
    state_23 <= reset | _GEN_23; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_24 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_24 <= state_23; // @[PRNG.scala 70:11]
    end
    state_25 <= reset | _GEN_25; // @[PRNG.scala 55:{49,49}]
    state_26 <= reset | _GEN_26; // @[PRNG.scala 55:{49,49}]
    state_27 <= reset | _GEN_27; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_28 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_28 <= state_27; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_29 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_29 <= state_28; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_30 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_30 <= state_29; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_31 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_31 <= state_30; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_32 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_32 <= state_31; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_33 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_33 <= state_32; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_34 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_34 <= state_33; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_35 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_35 <= state_34; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_36 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_36 <= state_35; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_37 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_37 <= state_36; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_38 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_38 <= state_37; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_39 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_39 <= state_38; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_40 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_40 <= state_39; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_41 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_41 <= state_40; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_42 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_42 <= state_41; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_43 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_43 <= state_42; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_44 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_44 <= state_43; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_45 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_45 <= state_44; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_46 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_46 <= state_45; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_47 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_47 <= state_46; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_48 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_48 <= state_47; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_49 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_49 <= state_48; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_50 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_50 <= state_49; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_51 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_51 <= state_50; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_52 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_52 <= state_51; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_53 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_53 <= state_52; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_54 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_54 <= state_53; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_55 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_55 <= state_54; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_56 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_56 <= state_55; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_57 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_57 <= state_56; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_58 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_58 <= state_57; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_59 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_59 <= state_58; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_60 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_60 <= state_59; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_61 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_61 <= state_60; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_62 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_62 <= state_61; // @[PRNG.scala 70:11]
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_63 <= 1'h0; // @[PRNG.scala 55:49]
    end else if (io_increment) begin // @[PRNG.scala 69:22]
      state_63 <= state_62; // @[PRNG.scala 70:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  state_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  state_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  state_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  state_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  state_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  state_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  state_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  state_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  state_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  state_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  state_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  state_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  state_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  state_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  state_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  state_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  state_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  state_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  state_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  state_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  state_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  state_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  state_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  state_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  state_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  state_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  state_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  state_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  state_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  state_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  state_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  state_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  state_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  state_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  state_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  state_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  state_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  state_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  state_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  state_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  state_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  state_63 = _RAND_63[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module moduled_prng(
  input         clock,
  input         reset,
  input         io_increment,
  output [63:0] io_PUB_VAR_HASH_LFSR
);
  wire  io_PUB_VAR_HASH_LFSR_prng_clock; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_reset; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_increment; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_20; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_21; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_22; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_23; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_24; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_25; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_26; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_27; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_28; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_29; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_30; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_31; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_32; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_33; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_34; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_35; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_36; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_37; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_38; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_39; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_40; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_41; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_42; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_43; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_44; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_45; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_46; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_47; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_48; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_49; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_50; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_51; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_52; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_53; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_54; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_55; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_56; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_57; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_58; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_59; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_60; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_61; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_62; // @[PRNG.scala 91:22]
  wire  io_PUB_VAR_HASH_LFSR_prng_io_out_63; // @[PRNG.scala 91:22]
  wire [7:0] io_PUB_VAR_HASH_LFSR_lo_lo_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_7,io_PUB_VAR_HASH_LFSR_prng_io_out_6,
    io_PUB_VAR_HASH_LFSR_prng_io_out_5,io_PUB_VAR_HASH_LFSR_prng_io_out_4,io_PUB_VAR_HASH_LFSR_prng_io_out_3,
    io_PUB_VAR_HASH_LFSR_prng_io_out_2,io_PUB_VAR_HASH_LFSR_prng_io_out_1,io_PUB_VAR_HASH_LFSR_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [15:0] io_PUB_VAR_HASH_LFSR_lo_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_15,io_PUB_VAR_HASH_LFSR_prng_io_out_14,
    io_PUB_VAR_HASH_LFSR_prng_io_out_13,io_PUB_VAR_HASH_LFSR_prng_io_out_12,io_PUB_VAR_HASH_LFSR_prng_io_out_11,
    io_PUB_VAR_HASH_LFSR_prng_io_out_10,io_PUB_VAR_HASH_LFSR_prng_io_out_9,io_PUB_VAR_HASH_LFSR_prng_io_out_8,
    io_PUB_VAR_HASH_LFSR_lo_lo_lo}; // @[PRNG.scala 95:17]
  wire [7:0] io_PUB_VAR_HASH_LFSR_lo_hi_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_23,io_PUB_VAR_HASH_LFSR_prng_io_out_22,
    io_PUB_VAR_HASH_LFSR_prng_io_out_21,io_PUB_VAR_HASH_LFSR_prng_io_out_20,io_PUB_VAR_HASH_LFSR_prng_io_out_19,
    io_PUB_VAR_HASH_LFSR_prng_io_out_18,io_PUB_VAR_HASH_LFSR_prng_io_out_17,io_PUB_VAR_HASH_LFSR_prng_io_out_16}; // @[PRNG.scala 95:17]
  wire [31:0] io_PUB_VAR_HASH_LFSR_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_31,io_PUB_VAR_HASH_LFSR_prng_io_out_30,
    io_PUB_VAR_HASH_LFSR_prng_io_out_29,io_PUB_VAR_HASH_LFSR_prng_io_out_28,io_PUB_VAR_HASH_LFSR_prng_io_out_27,
    io_PUB_VAR_HASH_LFSR_prng_io_out_26,io_PUB_VAR_HASH_LFSR_prng_io_out_25,io_PUB_VAR_HASH_LFSR_prng_io_out_24,
    io_PUB_VAR_HASH_LFSR_lo_hi_lo,io_PUB_VAR_HASH_LFSR_lo_lo}; // @[PRNG.scala 95:17]
  wire [7:0] io_PUB_VAR_HASH_LFSR_hi_lo_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_39,io_PUB_VAR_HASH_LFSR_prng_io_out_38,
    io_PUB_VAR_HASH_LFSR_prng_io_out_37,io_PUB_VAR_HASH_LFSR_prng_io_out_36,io_PUB_VAR_HASH_LFSR_prng_io_out_35,
    io_PUB_VAR_HASH_LFSR_prng_io_out_34,io_PUB_VAR_HASH_LFSR_prng_io_out_33,io_PUB_VAR_HASH_LFSR_prng_io_out_32}; // @[PRNG.scala 95:17]
  wire [15:0] io_PUB_VAR_HASH_LFSR_hi_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_47,io_PUB_VAR_HASH_LFSR_prng_io_out_46,
    io_PUB_VAR_HASH_LFSR_prng_io_out_45,io_PUB_VAR_HASH_LFSR_prng_io_out_44,io_PUB_VAR_HASH_LFSR_prng_io_out_43,
    io_PUB_VAR_HASH_LFSR_prng_io_out_42,io_PUB_VAR_HASH_LFSR_prng_io_out_41,io_PUB_VAR_HASH_LFSR_prng_io_out_40,
    io_PUB_VAR_HASH_LFSR_hi_lo_lo}; // @[PRNG.scala 95:17]
  wire [7:0] io_PUB_VAR_HASH_LFSR_hi_hi_lo = {io_PUB_VAR_HASH_LFSR_prng_io_out_55,io_PUB_VAR_HASH_LFSR_prng_io_out_54,
    io_PUB_VAR_HASH_LFSR_prng_io_out_53,io_PUB_VAR_HASH_LFSR_prng_io_out_52,io_PUB_VAR_HASH_LFSR_prng_io_out_51,
    io_PUB_VAR_HASH_LFSR_prng_io_out_50,io_PUB_VAR_HASH_LFSR_prng_io_out_49,io_PUB_VAR_HASH_LFSR_prng_io_out_48}; // @[PRNG.scala 95:17]
  wire [31:0] io_PUB_VAR_HASH_LFSR_hi = {io_PUB_VAR_HASH_LFSR_prng_io_out_63,io_PUB_VAR_HASH_LFSR_prng_io_out_62,
    io_PUB_VAR_HASH_LFSR_prng_io_out_61,io_PUB_VAR_HASH_LFSR_prng_io_out_60,io_PUB_VAR_HASH_LFSR_prng_io_out_59,
    io_PUB_VAR_HASH_LFSR_prng_io_out_58,io_PUB_VAR_HASH_LFSR_prng_io_out_57,io_PUB_VAR_HASH_LFSR_prng_io_out_56,
    io_PUB_VAR_HASH_LFSR_hi_hi_lo,io_PUB_VAR_HASH_LFSR_hi_lo}; // @[PRNG.scala 95:17]
  MaxPeriodFibonacciLFSR io_PUB_VAR_HASH_LFSR_prng ( // @[PRNG.scala 91:22]
    .clock(io_PUB_VAR_HASH_LFSR_prng_clock),
    .reset(io_PUB_VAR_HASH_LFSR_prng_reset),
    .io_increment(io_PUB_VAR_HASH_LFSR_prng_io_increment),
    .io_out_0(io_PUB_VAR_HASH_LFSR_prng_io_out_0),
    .io_out_1(io_PUB_VAR_HASH_LFSR_prng_io_out_1),
    .io_out_2(io_PUB_VAR_HASH_LFSR_prng_io_out_2),
    .io_out_3(io_PUB_VAR_HASH_LFSR_prng_io_out_3),
    .io_out_4(io_PUB_VAR_HASH_LFSR_prng_io_out_4),
    .io_out_5(io_PUB_VAR_HASH_LFSR_prng_io_out_5),
    .io_out_6(io_PUB_VAR_HASH_LFSR_prng_io_out_6),
    .io_out_7(io_PUB_VAR_HASH_LFSR_prng_io_out_7),
    .io_out_8(io_PUB_VAR_HASH_LFSR_prng_io_out_8),
    .io_out_9(io_PUB_VAR_HASH_LFSR_prng_io_out_9),
    .io_out_10(io_PUB_VAR_HASH_LFSR_prng_io_out_10),
    .io_out_11(io_PUB_VAR_HASH_LFSR_prng_io_out_11),
    .io_out_12(io_PUB_VAR_HASH_LFSR_prng_io_out_12),
    .io_out_13(io_PUB_VAR_HASH_LFSR_prng_io_out_13),
    .io_out_14(io_PUB_VAR_HASH_LFSR_prng_io_out_14),
    .io_out_15(io_PUB_VAR_HASH_LFSR_prng_io_out_15),
    .io_out_16(io_PUB_VAR_HASH_LFSR_prng_io_out_16),
    .io_out_17(io_PUB_VAR_HASH_LFSR_prng_io_out_17),
    .io_out_18(io_PUB_VAR_HASH_LFSR_prng_io_out_18),
    .io_out_19(io_PUB_VAR_HASH_LFSR_prng_io_out_19),
    .io_out_20(io_PUB_VAR_HASH_LFSR_prng_io_out_20),
    .io_out_21(io_PUB_VAR_HASH_LFSR_prng_io_out_21),
    .io_out_22(io_PUB_VAR_HASH_LFSR_prng_io_out_22),
    .io_out_23(io_PUB_VAR_HASH_LFSR_prng_io_out_23),
    .io_out_24(io_PUB_VAR_HASH_LFSR_prng_io_out_24),
    .io_out_25(io_PUB_VAR_HASH_LFSR_prng_io_out_25),
    .io_out_26(io_PUB_VAR_HASH_LFSR_prng_io_out_26),
    .io_out_27(io_PUB_VAR_HASH_LFSR_prng_io_out_27),
    .io_out_28(io_PUB_VAR_HASH_LFSR_prng_io_out_28),
    .io_out_29(io_PUB_VAR_HASH_LFSR_prng_io_out_29),
    .io_out_30(io_PUB_VAR_HASH_LFSR_prng_io_out_30),
    .io_out_31(io_PUB_VAR_HASH_LFSR_prng_io_out_31),
    .io_out_32(io_PUB_VAR_HASH_LFSR_prng_io_out_32),
    .io_out_33(io_PUB_VAR_HASH_LFSR_prng_io_out_33),
    .io_out_34(io_PUB_VAR_HASH_LFSR_prng_io_out_34),
    .io_out_35(io_PUB_VAR_HASH_LFSR_prng_io_out_35),
    .io_out_36(io_PUB_VAR_HASH_LFSR_prng_io_out_36),
    .io_out_37(io_PUB_VAR_HASH_LFSR_prng_io_out_37),
    .io_out_38(io_PUB_VAR_HASH_LFSR_prng_io_out_38),
    .io_out_39(io_PUB_VAR_HASH_LFSR_prng_io_out_39),
    .io_out_40(io_PUB_VAR_HASH_LFSR_prng_io_out_40),
    .io_out_41(io_PUB_VAR_HASH_LFSR_prng_io_out_41),
    .io_out_42(io_PUB_VAR_HASH_LFSR_prng_io_out_42),
    .io_out_43(io_PUB_VAR_HASH_LFSR_prng_io_out_43),
    .io_out_44(io_PUB_VAR_HASH_LFSR_prng_io_out_44),
    .io_out_45(io_PUB_VAR_HASH_LFSR_prng_io_out_45),
    .io_out_46(io_PUB_VAR_HASH_LFSR_prng_io_out_46),
    .io_out_47(io_PUB_VAR_HASH_LFSR_prng_io_out_47),
    .io_out_48(io_PUB_VAR_HASH_LFSR_prng_io_out_48),
    .io_out_49(io_PUB_VAR_HASH_LFSR_prng_io_out_49),
    .io_out_50(io_PUB_VAR_HASH_LFSR_prng_io_out_50),
    .io_out_51(io_PUB_VAR_HASH_LFSR_prng_io_out_51),
    .io_out_52(io_PUB_VAR_HASH_LFSR_prng_io_out_52),
    .io_out_53(io_PUB_VAR_HASH_LFSR_prng_io_out_53),
    .io_out_54(io_PUB_VAR_HASH_LFSR_prng_io_out_54),
    .io_out_55(io_PUB_VAR_HASH_LFSR_prng_io_out_55),
    .io_out_56(io_PUB_VAR_HASH_LFSR_prng_io_out_56),
    .io_out_57(io_PUB_VAR_HASH_LFSR_prng_io_out_57),
    .io_out_58(io_PUB_VAR_HASH_LFSR_prng_io_out_58),
    .io_out_59(io_PUB_VAR_HASH_LFSR_prng_io_out_59),
    .io_out_60(io_PUB_VAR_HASH_LFSR_prng_io_out_60),
    .io_out_61(io_PUB_VAR_HASH_LFSR_prng_io_out_61),
    .io_out_62(io_PUB_VAR_HASH_LFSR_prng_io_out_62),
    .io_out_63(io_PUB_VAR_HASH_LFSR_prng_io_out_63)
  );
  assign io_PUB_VAR_HASH_LFSR = {io_PUB_VAR_HASH_LFSR_hi,io_PUB_VAR_HASH_LFSR_lo}; // @[PRNG.scala 95:17]
  assign io_PUB_VAR_HASH_LFSR_prng_clock = clock;
  assign io_PUB_VAR_HASH_LFSR_prng_reset = reset;
  assign io_PUB_VAR_HASH_LFSR_prng_io_increment = io_increment; // @[PRNG.scala 94:23]
endmodule
module MaxPeriodFibonacciLFSR_1(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19,
  output  io_out_20,
  output  io_out_21,
  output  io_out_22,
  output  io_out_23,
  output  io_out_24,
  output  io_out_25,
  output  io_out_26,
  output  io_out_27,
  output  io_out_28,
  output  io_out_29,
  output  io_out_30,
  output  io_out_31,
  output  io_out_32,
  output  io_out_33,
  output  io_out_34,
  output  io_out_35,
  output  io_out_36,
  output  io_out_37,
  output  io_out_38,
  output  io_out_39,
  output  io_out_40,
  output  io_out_41,
  output  io_out_42,
  output  io_out_43,
  output  io_out_44,
  output  io_out_45,
  output  io_out_46
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  reg  state_16; // @[PRNG.scala 55:49]
  reg  state_17; // @[PRNG.scala 55:49]
  reg  state_18; // @[PRNG.scala 55:49]
  reg  state_19; // @[PRNG.scala 55:49]
  reg  state_20; // @[PRNG.scala 55:49]
  reg  state_21; // @[PRNG.scala 55:49]
  reg  state_22; // @[PRNG.scala 55:49]
  reg  state_23; // @[PRNG.scala 55:49]
  reg  state_24; // @[PRNG.scala 55:49]
  reg  state_25; // @[PRNG.scala 55:49]
  reg  state_26; // @[PRNG.scala 55:49]
  reg  state_27; // @[PRNG.scala 55:49]
  reg  state_28; // @[PRNG.scala 55:49]
  reg  state_29; // @[PRNG.scala 55:49]
  reg  state_30; // @[PRNG.scala 55:49]
  reg  state_31; // @[PRNG.scala 55:49]
  reg  state_32; // @[PRNG.scala 55:49]
  reg  state_33; // @[PRNG.scala 55:49]
  reg  state_34; // @[PRNG.scala 55:49]
  reg  state_35; // @[PRNG.scala 55:49]
  reg  state_36; // @[PRNG.scala 55:49]
  reg  state_37; // @[PRNG.scala 55:49]
  reg  state_38; // @[PRNG.scala 55:49]
  reg  state_39; // @[PRNG.scala 55:49]
  reg  state_40; // @[PRNG.scala 55:49]
  reg  state_41; // @[PRNG.scala 55:49]
  reg  state_42; // @[PRNG.scala 55:49]
  reg  state_43; // @[PRNG.scala 55:49]
  reg  state_44; // @[PRNG.scala 55:49]
  reg  state_45; // @[PRNG.scala 55:49]
  reg  state_46; // @[PRNG.scala 55:49]
  wire  _T = state_46 ^ state_41; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  assign io_out_16 = state_16; // @[PRNG.scala 78:10]
  assign io_out_17 = state_17; // @[PRNG.scala 78:10]
  assign io_out_18 = state_18; // @[PRNG.scala 78:10]
  assign io_out_19 = state_19; // @[PRNG.scala 78:10]
  assign io_out_20 = state_20; // @[PRNG.scala 78:10]
  assign io_out_21 = state_21; // @[PRNG.scala 78:10]
  assign io_out_22 = state_22; // @[PRNG.scala 78:10]
  assign io_out_23 = state_23; // @[PRNG.scala 78:10]
  assign io_out_24 = state_24; // @[PRNG.scala 78:10]
  assign io_out_25 = state_25; // @[PRNG.scala 78:10]
  assign io_out_26 = state_26; // @[PRNG.scala 78:10]
  assign io_out_27 = state_27; // @[PRNG.scala 78:10]
  assign io_out_28 = state_28; // @[PRNG.scala 78:10]
  assign io_out_29 = state_29; // @[PRNG.scala 78:10]
  assign io_out_30 = state_30; // @[PRNG.scala 78:10]
  assign io_out_31 = state_31; // @[PRNG.scala 78:10]
  assign io_out_32 = state_32; // @[PRNG.scala 78:10]
  assign io_out_33 = state_33; // @[PRNG.scala 78:10]
  assign io_out_34 = state_34; // @[PRNG.scala 78:10]
  assign io_out_35 = state_35; // @[PRNG.scala 78:10]
  assign io_out_36 = state_36; // @[PRNG.scala 78:10]
  assign io_out_37 = state_37; // @[PRNG.scala 78:10]
  assign io_out_38 = state_38; // @[PRNG.scala 78:10]
  assign io_out_39 = state_39; // @[PRNG.scala 78:10]
  assign io_out_40 = state_40; // @[PRNG.scala 78:10]
  assign io_out_41 = state_41; // @[PRNG.scala 78:10]
  assign io_out_42 = state_42; // @[PRNG.scala 78:10]
  assign io_out_43 = state_43; // @[PRNG.scala 78:10]
  assign io_out_44 = state_44; // @[PRNG.scala 78:10]
  assign io_out_45 = state_45; // @[PRNG.scala 78:10]
  assign io_out_46 = state_46; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    state_2 <= reset | state_1; // @[PRNG.scala 55:{49,49}]
    state_3 <= reset | state_2; // @[PRNG.scala 55:{49,49}]
    state_4 <= reset | state_3; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    state_6 <= reset | state_5; // @[PRNG.scala 55:{49,49}]
    state_7 <= reset | state_6; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    state_9 <= reset | state_8; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    state_11 <= reset | state_10; // @[PRNG.scala 55:{49,49}]
    state_12 <= reset | state_11; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    state_14 <= reset | state_13; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
    state_16 <= reset | state_15; // @[PRNG.scala 55:{49,49}]
    state_17 <= reset | state_16; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_18 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_18 <= state_17;
    end
    state_19 <= reset | state_18; // @[PRNG.scala 55:{49,49}]
    state_20 <= reset | state_19; // @[PRNG.scala 55:{49,49}]
    state_21 <= reset | state_20; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_22 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_22 <= state_21;
    end
    state_23 <= reset | state_22; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_24 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_24 <= state_23;
    end
    state_25 <= reset | state_24; // @[PRNG.scala 55:{49,49}]
    state_26 <= reset | state_25; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_27 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_27 <= state_26;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_28 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_28 <= state_27;
    end
    state_29 <= reset | state_28; // @[PRNG.scala 55:{49,49}]
    state_30 <= reset | state_29; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_31 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_31 <= state_30;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_32 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_32 <= state_31;
    end
    state_33 <= reset | state_32; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_34 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_34 <= state_33;
    end
    state_35 <= reset | state_34; // @[PRNG.scala 55:{49,49}]
    state_36 <= reset | state_35; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_37 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_37 <= state_36;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_38 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_38 <= state_37;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_39 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_39 <= state_38;
    end
    state_40 <= reset | state_39; // @[PRNG.scala 55:{49,49}]
    state_41 <= reset | state_40; // @[PRNG.scala 55:{49,49}]
    state_42 <= reset | state_41; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_43 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_43 <= state_42;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_44 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_44 <= state_43;
    end
    state_45 <= reset | state_44; // @[PRNG.scala 55:{49,49}]
    state_46 <= reset | state_45; // @[PRNG.scala 55:{49,49}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  state_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  state_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  state_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  state_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  state_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  state_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  state_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  state_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  state_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  state_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  state_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  state_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  state_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  state_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  state_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  state_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  state_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  state_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  state_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  state_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  state_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  state_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  state_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  state_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  state_46 = _RAND_46[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SE(
  input          clock,
  input          reset,
  input  [7:0]   io_in_inst,
  input  [315:0] io_in_op1,
  input  [315:0] io_in_op2,
  input          io_in_valid,
  output         io_in_ready,
  input          io_out_ready,
  output [315:0] io_out_result,
  output         io_out_valid,
  output         io_out_op1_hash_compare,
  output         io_out_op2_hash_compare
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [319:0] _RAND_1;
  reg [319:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [319:0] _RAND_16;
  reg [319:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [255:0] _RAND_52;
  reg [319:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] seoperation_io_inst; // @[SE.scala 166:33]
  wire  seoperation_io_in_valid; // @[SE.scala 166:33]
  wire [63:0] seoperation_io_op1_input; // @[SE.scala 166:33]
  wire [63:0] seoperation_io_op2_input; // @[SE.scala 166:33]
  wire [63:0] seoperation_io_result; // @[SE.scala 166:33]
  wire  seoperation_io_out_valid; // @[SE.scala 166:33]
  wire  aes_invcipher_op1_clock; // @[SE.scala 174:39]
  wire  aes_invcipher_op1_reset; // @[SE.scala 174:39]
  wire  aes_invcipher_op1_io_input_valid; // @[SE.scala 174:39]
  wire [255:0] aes_invcipher_op1_io_input_text; // @[SE.scala 174:39]
  wire [255:0] aes_invcipher_op1_io_output_text; // @[SE.scala 174:39]
  wire  aes_invcipher_op1_io_output_valid; // @[SE.scala 174:39]
  wire  aes_invcipher_op2_clock; // @[SE.scala 175:39]
  wire  aes_invcipher_op2_reset; // @[SE.scala 175:39]
  wire  aes_invcipher_op2_io_input_valid; // @[SE.scala 175:39]
  wire [255:0] aes_invcipher_op2_io_input_text; // @[SE.scala 175:39]
  wire [255:0] aes_invcipher_op2_io_output_text; // @[SE.scala 175:39]
  wire  aes_invcipher_op2_io_output_valid; // @[SE.scala 175:39]
  wire  aes_cipher_clock; // @[SE.scala 182:57]
  wire  aes_cipher_reset; // @[SE.scala 182:57]
  wire  aes_cipher_io_input_valid; // @[SE.scala 182:57]
  wire [127:0] aes_cipher_io_input_op1; // @[SE.scala 182:57]
  wire [127:0] aes_cipher_io_input_op2; // @[SE.scala 182:57]
  wire [255:0] aes_cipher_io_output_text; // @[SE.scala 182:57]
  wire  aes_cipher_io_output_valid; // @[SE.scala 182:57]
  wire  aes_cipher_for_hash_C_clock; // @[SE.scala 185:49]
  wire  aes_cipher_for_hash_C_reset; // @[SE.scala 185:49]
  wire  aes_cipher_for_hash_C_io_input_valid; // @[SE.scala 185:49]
  wire [127:0] aes_cipher_for_hash_C_io_input_text; // @[SE.scala 185:49]
  wire [127:0] aes_cipher_for_hash_C_io_output_text; // @[SE.scala 185:49]
  wire  aes_cipher_for_hash_C_io_output_valid; // @[SE.scala 185:49]
  wire  aes_cipher_for_op1_clock; // @[SE.scala 186:49]
  wire  aes_cipher_for_op1_reset; // @[SE.scala 186:49]
  wire  aes_cipher_for_op1_io_input_valid; // @[SE.scala 186:49]
  wire [127:0] aes_cipher_for_op1_io_input_text; // @[SE.scala 186:49]
  wire [127:0] aes_cipher_for_op1_io_output_text; // @[SE.scala 186:49]
  wire  aes_cipher_for_op1_io_output_valid; // @[SE.scala 186:49]
  wire  aes_cipher_for_op2_clock; // @[SE.scala 187:49]
  wire  aes_cipher_for_op2_reset; // @[SE.scala 187:49]
  wire  aes_cipher_for_op2_io_input_valid; // @[SE.scala 187:49]
  wire [127:0] aes_cipher_for_op2_io_input_text; // @[SE.scala 187:49]
  wire [127:0] aes_cipher_for_op2_io_output_text; // @[SE.scala 187:49]
  wire  aes_cipher_for_op2_io_output_valid; // @[SE.scala 187:49]
  wire  aes_cipher_for_pub_var_clock; // @[SE.scala 188:44]
  wire  aes_cipher_for_pub_var_reset; // @[SE.scala 188:44]
  wire  aes_cipher_for_pub_var_io_input_valid; // @[SE.scala 188:44]
  wire [127:0] aes_cipher_for_pub_var_io_input_text; // @[SE.scala 188:44]
  wire [127:0] aes_cipher_for_pub_var_io_output_text; // @[SE.scala 188:44]
  wire  aes_cipher_for_pub_var_io_output_valid; // @[SE.scala 188:44]
  wire [315:0] PRC_0_io_op1; // @[SE.scala 211:23]
  wire [315:0] PRC_0_io_op2; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_inst; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_0; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_1; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_2; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_3; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_4; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_5; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_6; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_7; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_8; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_9; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_10; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_11; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_12; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_13; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_14; // @[SE.scala 211:23]
  wire [7:0] PRC_0_io_out_15; // @[SE.scala 211:23]
  wire [59:0] HC_op1_io_hash_orig; // @[SE.scala 214:28]
  wire [59:0] HC_op1_io_hash_regenerated; // @[SE.scala 214:28]
  wire  HC_op1_io_valid_in; // @[SE.scala 214:28]
  wire  HC_op1_io_valid_out; // @[SE.scala 214:28]
  wire  HC_op1_io_compare_result; // @[SE.scala 214:28]
  wire [59:0] HC_op2_io_hash_orig; // @[SE.scala 215:28]
  wire [59:0] HC_op2_io_hash_regenerated; // @[SE.scala 215:28]
  wire  HC_op2_io_valid_in; // @[SE.scala 215:28]
  wire  HC_op2_io_valid_out; // @[SE.scala 215:28]
  wire  HC_op2_io_compare_result; // @[SE.scala 215:28]
  wire  VID_0_io_pub_priv_opA; // @[SE.scala 219:27]
  wire  VID_0_io_pub_priv_opB; // @[SE.scala 219:27]
  wire [15:0] VID_0_io_version_id_opA; // @[SE.scala 219:27]
  wire [15:0] VID_0_io_version_id_opB; // @[SE.scala 219:27]
  wire  VID_0_io_valid_in; // @[SE.scala 219:27]
  wire  VID_0_io_valid_out; // @[SE.scala 219:27]
  wire [15:0] VID_0_io_version_id_out; // @[SE.scala 219:27]
  wire  VID_0_io_pub_priv_out; // @[SE.scala 219:27]
  wire  moduled_prng_pub_var_clock; // @[SE.scala 246:42]
  wire  moduled_prng_pub_var_reset; // @[SE.scala 246:42]
  wire  moduled_prng_pub_var_io_increment; // @[SE.scala 246:42]
  wire [63:0] moduled_prng_pub_var_io_PUB_VAR_HASH_LFSR; // @[SE.scala 246:42]
  wire  bit47_randnum_prng_clock; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_reset; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_20; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_21; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_22; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_23; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_24; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_25; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_26; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_27; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_28; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_29; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_30; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_31; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_32; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_33; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_34; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_35; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_36; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_37; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_38; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_39; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_40; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_41; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_42; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_43; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_44; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_45; // @[PRNG.scala 91:22]
  wire  bit47_randnum_prng_io_out_46; // @[PRNG.scala 91:22]
  reg [7:0] inst_buffer; // @[Reg.scala 16:16]
  reg [315:0] op1_buffer; // @[Reg.scala 16:16]
  reg [315:0] op2_buffer; // @[Reg.scala 16:16]
  reg  ready_for_input; // @[SE.scala 225:38]
  reg  lv1ok_buffer; // @[SE.scala 232:42]
  reg  lv2ok_buffer; // @[SE.scala 233:42]
  reg  lv3ok_buffer; // @[SE.scala 234:42]
  reg  lv4ok_buffer; // @[SE.scala 235:42]
  wire  is_enc_const = 8'hb0 == inst_buffer; // @[SE.scala 239:41]
  wire  is_enc_var = 8'ha0 == inst_buffer; // @[SE.scala 240:40]
  wire  is_enc_var_hash = 8'hb8 == inst_buffer; // @[SE.scala 241:44]
  wire  is_enc_inst = is_enc_const & is_enc_var & is_enc_var_hash; // @[SE.scala 242:53]
  reg [63:0] pub_var_hash_register; // @[SE.scala 251:40]
  reg  output_valid; // @[SE.scala 272:35]
  wire  _next_ready_for_input_T = io_in_valid & io_in_ready; // @[SE.scala 281:61]
  wire  _next_ready_for_input_T_1 = io_out_valid & io_out_ready; // @[SE.scala 281:105]
  reg  ready_for_input_REG; // @[SE.scala 282:59]
  wire  _next_lv1ok_buffer_T_1 = output_valid ? 1'h0 : lv1ok_buffer; // @[SE.scala 286:81]
  reg  lv1ok_buffer_REG; // @[SE.scala 287:51]
  wire  _T_3 = ~lv3ok_buffer; // @[SE.scala 290:47]
  wire  _T_5 = ~lv4ok_buffer; // @[SE.scala 290:64]
  wire  _T_6 = lv1ok_buffer & ~lv2ok_buffer & ~lv3ok_buffer & ~lv4ok_buffer; // @[SE.scala 290:61]
  wire  _T_8 = ~reset; // @[SE.scala 291:23]
  wire [255:0] ciph_op1 = op1_buffer[255:0]; // @[SE.scala 309:53]
  wire [127:0] ciph_op1_val = ciph_op1[127:0]; // @[SE.scala 310:51]
  wire [127:0] ciph_op1_hash = ciph_op1[255:128]; // @[SE.scala 311:51]
  wire [255:0] ciph_op2 = op2_buffer[255:0]; // @[SE.scala 312:53]
  wire [127:0] ciph_op2_val = ciph_op2[127:0]; // @[SE.scala 313:51]
  wire [127:0] ciph_op2_hash = ciph_op2[255:128]; // @[SE.scala 314:51]
  reg  lv2_AES_valid; // @[SE.scala 315:42]
  reg  tmp_1; // @[SE.scala 316:58]
  wire  _next_tmp_1_T_2 = output_valid ? 1'h0 : tmp_1; // @[SE.scala 324:101]
  reg  lv2_AES_valid_REG; // @[SE.scala 325:51]
  reg  tmp_1_REG; // @[SE.scala 326:59]
  wire [7:0] connected_reversed_plaintext_buffer_1 = PRC_0_io_out_1; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_0 = PRC_0_io_out_0; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_3 = PRC_0_io_out_3; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_2 = PRC_0_io_out_2; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_5 = PRC_0_io_out_5; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_4 = PRC_0_io_out_4; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_7 = PRC_0_io_out_7; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_6 = PRC_0_io_out_6; // @[SE.scala 305:51 306:49]
  wire [63:0] aes_cipher_for_hash_C_io_input_text_lo = {connected_reversed_plaintext_buffer_7,
    connected_reversed_plaintext_buffer_6,connected_reversed_plaintext_buffer_5,connected_reversed_plaintext_buffer_4,
    connected_reversed_plaintext_buffer_3,connected_reversed_plaintext_buffer_2,connected_reversed_plaintext_buffer_1,
    connected_reversed_plaintext_buffer_0}; // @[SE.scala 335:96]
  wire [7:0] connected_reversed_plaintext_buffer_9 = PRC_0_io_out_9; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_8 = PRC_0_io_out_8; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_11 = PRC_0_io_out_11; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_10 = PRC_0_io_out_10; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_13 = PRC_0_io_out_13; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_12 = PRC_0_io_out_12; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_15 = PRC_0_io_out_15; // @[SE.scala 305:51 306:49]
  wire [7:0] connected_reversed_plaintext_buffer_14 = PRC_0_io_out_14; // @[SE.scala 305:51 306:49]
  wire [63:0] aes_cipher_for_hash_C_io_input_text_hi = {connected_reversed_plaintext_buffer_15,
    connected_reversed_plaintext_buffer_14,connected_reversed_plaintext_buffer_13,connected_reversed_plaintext_buffer_12
    ,connected_reversed_plaintext_buffer_11,connected_reversed_plaintext_buffer_10,connected_reversed_plaintext_buffer_9
    ,connected_reversed_plaintext_buffer_8}; // @[SE.scala 335:96]
  reg [315:0] lv2_op1_buffer; // @[Reg.scala 16:16]
  reg [315:0] lv2_op2_buffer; // @[Reg.scala 16:16]
  reg [127:0] hash_C_original_buffer; // @[Reg.scala 16:16]
  reg  hash_C_original_buffer_valid; // @[SE.scala 348:66]
  reg [127:0] decrypted_op1_val_buffer; // @[Reg.scala 16:16]
  reg [127:0] decrypted_op1_hash_buffer; // @[Reg.scala 16:16]
  reg [127:0] decrypted_op2_val_buffer; // @[Reg.scala 16:16]
  reg [127:0] decrypted_op2_hash_buffer; // @[Reg.scala 16:16]
  reg  lv3_AES_valid; // @[SE.scala 359:42]
  reg  tmp_2; // @[SE.scala 360:58]
  wire  _next_hash_C_original_buffer_valid_T = output_valid ? 1'h0 : hash_C_original_buffer_valid; // @[SE.scala 364:102]
  reg  hash_C_original_buffer_valid_REG; // @[SE.scala 365:59]
  wire  lv2_bypass = lv1ok_buffer & is_enc_inst; // @[SE.scala 383:39]
  wire  _next_lv2ok_buffer_T_3 = output_valid ? 1'h0 : lv2ok_buffer; // @[SE.scala 384:180]
  reg  lv2ok_buffer_REG; // @[SE.scala 385:51]
  wire  _next_tmp_2_T_2 = output_valid ? 1'h0 : tmp_2; // @[SE.scala 392:101]
  reg  lv3_AES_valid_REG; // @[SE.scala 393:51]
  reg  tmp_2_REG; // @[SE.scala 394:59]
  wire  _T_22 = lv2ok_buffer & _T_3 & _T_5; // @[SE.scala 397:44]
  wire [63:0] _op1_plaintext_64_T_3 = is_enc_var | is_enc_const ? op1_buffer[255:192] : decrypted_op1_val_buffer[127:64]
    ; // @[SE.scala 439:132]
  wire  opA_pub_priv = decrypted_op1_val_buffer[16]; // @[SE.scala 448:35]
  wire  opB_pub_priv = decrypted_op2_val_buffer[16]; // @[SE.scala 449:35]
  reg [15:0] verID_C; // @[Reg.scala 16:16]
  reg  verID_C_valid; // @[SE.scala 458:36]
  wire  _next_verID_C_valid_T = output_valid ? 1'h0 : verID_C_valid; // @[SE.scala 460:79]
  reg  verID_C_valid_REG; // @[SE.scala 461:51]
  reg  pub_prv_bit; // @[Reg.scala 16:16]
  wire [4:0] bit47_randnum_lo_lo_lo = {bit47_randnum_prng_io_out_4,bit47_randnum_prng_io_out_3,
    bit47_randnum_prng_io_out_2,bit47_randnum_prng_io_out_1,bit47_randnum_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [10:0] bit47_randnum_lo_lo = {bit47_randnum_prng_io_out_10,bit47_randnum_prng_io_out_9,
    bit47_randnum_prng_io_out_8,bit47_randnum_prng_io_out_7,bit47_randnum_prng_io_out_6,bit47_randnum_prng_io_out_5,
    bit47_randnum_lo_lo_lo}; // @[PRNG.scala 95:17]
  wire [5:0] bit47_randnum_lo_hi_lo = {bit47_randnum_prng_io_out_16,bit47_randnum_prng_io_out_15,
    bit47_randnum_prng_io_out_14,bit47_randnum_prng_io_out_13,bit47_randnum_prng_io_out_12,bit47_randnum_prng_io_out_11}
    ; // @[PRNG.scala 95:17]
  wire [22:0] bit47_randnum_lo = {bit47_randnum_prng_io_out_22,bit47_randnum_prng_io_out_21,bit47_randnum_prng_io_out_20
    ,bit47_randnum_prng_io_out_19,bit47_randnum_prng_io_out_18,bit47_randnum_prng_io_out_17,bit47_randnum_lo_hi_lo,
    bit47_randnum_lo_lo}; // @[PRNG.scala 95:17]
  wire [5:0] bit47_randnum_hi_lo_lo = {bit47_randnum_prng_io_out_28,bit47_randnum_prng_io_out_27,
    bit47_randnum_prng_io_out_26,bit47_randnum_prng_io_out_25,bit47_randnum_prng_io_out_24,bit47_randnum_prng_io_out_23}
    ; // @[PRNG.scala 95:17]
  wire [11:0] bit47_randnum_hi_lo = {bit47_randnum_prng_io_out_34,bit47_randnum_prng_io_out_33,
    bit47_randnum_prng_io_out_32,bit47_randnum_prng_io_out_31,bit47_randnum_prng_io_out_30,bit47_randnum_prng_io_out_29,
    bit47_randnum_hi_lo_lo}; // @[PRNG.scala 95:17]
  wire [5:0] bit47_randnum_hi_hi_lo = {bit47_randnum_prng_io_out_40,bit47_randnum_prng_io_out_39,
    bit47_randnum_prng_io_out_38,bit47_randnum_prng_io_out_37,bit47_randnum_prng_io_out_36,bit47_randnum_prng_io_out_35}
    ; // @[PRNG.scala 95:17]
  wire [46:0] bit47_randnum = {bit47_randnum_prng_io_out_46,bit47_randnum_prng_io_out_45,bit47_randnum_prng_io_out_44,
    bit47_randnum_prng_io_out_43,bit47_randnum_prng_io_out_42,bit47_randnum_prng_io_out_41,bit47_randnum_hi_hi_lo,
    bit47_randnum_hi_lo,bit47_randnum_lo}; // @[PRNG.scala 95:17]
  wire [110:0] non_enc_padded_result_hi_hi = {seoperation_io_result,bit47_randnum_prng_io_out_46,
    bit47_randnum_prng_io_out_45,bit47_randnum_prng_io_out_44,bit47_randnum_prng_io_out_43,bit47_randnum_prng_io_out_42,
    bit47_randnum_prng_io_out_41,bit47_randnum_hi_hi_lo,bit47_randnum_hi_lo,bit47_randnum_lo}; // @[Cat.scala 31:58]
  wire [255:0] non_enc_padded_result = {non_enc_padded_result_hi_hi,pub_prv_bit,verID_C,lv2_op1_buffer[315:256],
    lv2_op2_buffer[315:256],inst_buffer}; // @[Cat.scala 31:58]
  wire [59:0] enc_datahash = is_enc_var ? seoperation_io_result[59:0] : moduled_prng_pub_var_io_PUB_VAR_HASH_LFSR[59:0]; // @[SE.scala 471:25]
  wire [255:0] enc_padded_result = {non_enc_padded_result_hi_hi,pub_prv_bit,verID_C,enc_datahash,60'h0,inst_buffer}; // @[Cat.scala 31:58]
  wire  _result_buffer_T = seoperation_io_out_valid & verID_C_valid; // @[SE.scala 483:117]
  reg [255:0] result_buffer; // @[Reg.scala 16:16]
  reg  result_valid_buffer; // @[SE.scala 484:66]
  reg  hash_C_buffer_valid; // @[SE.scala 486:66]
  reg [59:0] hash_C_buffer; // @[Reg.scala 16:16]
  reg  op1_rehash_result_buffer_valid; // @[SE.scala 488:58]
  reg [127:0] op1_rehash_result_bit; // @[Reg.scala 16:16]
  reg  op2_rehash_result_buffer_valid; // @[SE.scala 490:58]
  reg [127:0] op2_rehash_result_bit; // @[Reg.scala 16:16]
  wire  _next_op1_rehash_result_buffer_valid_T = output_valid ? 1'h0 : op1_rehash_result_buffer_valid; // @[SE.scala 501:111]
  wire  _next_op2_rehash_result_buffer_valid_T = output_valid ? 1'h0 : op2_rehash_result_buffer_valid; // @[SE.scala 502:111]
  reg  op1_rehash_result_buffer_valid_REG; // @[SE.scala 503:75]
  reg  op2_rehash_result_buffer_valid_REG; // @[SE.scala 504:75]
  wire  _next_hash_C_buffer_valid_T = output_valid ? 1'h0 : hash_C_buffer_valid; // @[SE.scala 508:88]
  reg  hash_C_buffer_valid_REG; // @[SE.scala 509:50]
  wire  _n_result_valid_buffer_T = output_valid ? 1'h0 : result_valid_buffer; // @[SE.scala 513:60]
  reg  result_valid_buffer_REG; // @[SE.scala 514:39]
  wire  _next_lv3ok_buffer_T_3 = output_valid ? 1'h0 : lv3ok_buffer; // @[SE.scala 518:165]
  reg  lv3ok_buffer_REG; // @[SE.scala 519:51]
  wire  _T_224 = lv3ok_buffer & _T_5; // @[SE.scala 522:27]
  wire [7:0] result_buffer_vectorized_0 = result_buffer[7:0]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_1 = result_buffer[15:8]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_2 = result_buffer[23:16]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_3 = result_buffer[31:24]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_4 = result_buffer[39:32]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_5 = result_buffer[47:40]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_6 = result_buffer[55:48]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_7 = result_buffer[63:56]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_8 = result_buffer[71:64]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_9 = result_buffer[79:72]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_10 = result_buffer[87:80]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_11 = result_buffer[95:88]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_12 = result_buffer[103:96]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_13 = result_buffer[111:104]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_14 = result_buffer[119:112]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_15 = result_buffer[127:120]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_16 = result_buffer[135:128]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_17 = result_buffer[143:136]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_18 = result_buffer[151:144]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_19 = result_buffer[159:152]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_20 = result_buffer[167:160]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_21 = result_buffer[175:168]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_22 = result_buffer[183:176]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_23 = result_buffer[191:184]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_24 = result_buffer[199:192]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_25 = result_buffer[207:200]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_26 = result_buffer[215:208]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_27 = result_buffer[223:216]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_28 = result_buffer[231:224]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_29 = result_buffer[239:232]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_30 = result_buffer[247:240]; // @[SE.scala 542:110]
  wire [7:0] result_buffer_vectorized_31 = result_buffer[255:248]; // @[SE.scala 542:110]
  wire [63:0] aes_input_reverse_bit_lo_lo = {result_buffer_vectorized_24,result_buffer_vectorized_25,
    result_buffer_vectorized_26,result_buffer_vectorized_27,result_buffer_vectorized_28,result_buffer_vectorized_29,
    result_buffer_vectorized_30,result_buffer_vectorized_31}; // @[Cat.scala 31:58]
  wire [127:0] aes_input_reverse_bit_lo = {result_buffer_vectorized_16,result_buffer_vectorized_17,
    result_buffer_vectorized_18,result_buffer_vectorized_19,result_buffer_vectorized_20,result_buffer_vectorized_21,
    result_buffer_vectorized_22,result_buffer_vectorized_23,aes_input_reverse_bit_lo_lo}; // @[Cat.scala 31:58]
  wire [63:0] aes_input_reverse_bit_hi_lo = {result_buffer_vectorized_8,result_buffer_vectorized_9,
    result_buffer_vectorized_10,result_buffer_vectorized_11,result_buffer_vectorized_12,result_buffer_vectorized_13,
    result_buffer_vectorized_14,result_buffer_vectorized_15}; // @[Cat.scala 31:58]
  wire [255:0] aes_input_reverse_bit = {result_buffer_vectorized_0,result_buffer_vectorized_1,result_buffer_vectorized_2
    ,result_buffer_vectorized_3,result_buffer_vectorized_4,result_buffer_vectorized_5,result_buffer_vectorized_6,
    result_buffer_vectorized_7,aes_input_reverse_bit_hi_lo,aes_input_reverse_bit_lo}; // @[Cat.scala 31:58]
  reg  lv4_AES_valid; // @[SE.scala 548:42]
  reg  tmp_3; // @[SE.scala 549:58]
  wire  _next_tmp_3_T_2 = output_valid ? 1'h0 : tmp_3; // @[SE.scala 556:101]
  reg  lv4_AES_valid_REG; // @[SE.scala 557:51]
  reg  tmp_3_REG; // @[SE.scala 558:59]
  reg  output_buffer_enc_valid; // @[SE.scala 584:66]
  reg [255:0] output_buffer_enc; // @[Reg.scala 16:16]
  reg [315:0] output_buffer; // @[SE.scala 586:74]
  wire  _hash_compare_result_op1_T = ~is_enc_var_hash; // @[SE.scala 587:90]
  wire  _hash_compare_result_op1_T_1 = HC_op1_io_compare_result | ~is_enc_var_hash; // @[SE.scala 587:86]
  reg  hash_compare_result_op1; // @[Reg.scala 16:16]
  reg  hash_compare_result_op1_valid; // @[SE.scala 588:58]
  wire  _hash_compare_result_op2_T_1 = HC_op2_io_compare_result | _hash_compare_result_op1_T; // @[SE.scala 589:86]
  reg  hash_compare_result_op2; // @[Reg.scala 16:16]
  reg  hash_compare_result_op2_valid; // @[SE.scala 590:58]
  wire  _next_output_buffer_enc_valid_T = output_valid ? 1'h0 : output_buffer_enc_valid; // @[SE.scala 594:94]
  reg  output_buffer_enc_valid_REG; // @[SE.scala 595:67]
  wire  _next_lv4ok_buffer_T_2 = output_valid ? 1'h0 : lv4ok_buffer; // @[SE.scala 598:143]
  reg  lv4ok_buffer_REG; // @[SE.scala 599:51]
  wire  _GEN_196 = _next_ready_for_input_T_1 ? 1'h0 : output_valid; // @[SE.scala 603:50 604:30 272:35]
  wire  _GEN_197 = lv4ok_buffer | _GEN_196; // @[SE.scala 601:28 602:30]
  wire  _next_hash_compare_result_op1_valid_T = output_valid ? 1'h0 : hash_compare_result_op1_valid; // @[SE.scala 610:96]
  wire  _next_hash_compare_result_op2_valid_T = output_valid ? 1'h0 : hash_compare_result_op2_valid; // @[SE.scala 611:96]
  reg  hash_compare_result_op1_valid_REG; // @[SE.scala 612:67]
  reg  hash_compare_result_op2_valid_REG; // @[SE.scala 613:67]
  wire [315:0] output_connect = {hash_C_buffer,output_buffer_enc}; // @[Cat.scala 31:58]
  wire  compare_hash_total = hash_compare_result_op1 & hash_compare_result_op1_valid & hash_compare_result_op2 &
    hash_compare_result_op2_valid; // @[SE.scala 621:128]
  SEOperation seoperation ( // @[SE.scala 166:33]
    .io_inst(seoperation_io_inst),
    .io_in_valid(seoperation_io_in_valid),
    .io_op1_input(seoperation_io_op1_input),
    .io_op2_input(seoperation_io_op2_input),
    .io_result(seoperation_io_result),
    .io_out_valid(seoperation_io_out_valid)
  );
  AESDecrypt aes_invcipher_op1 ( // @[SE.scala 174:39]
    .clock(aes_invcipher_op1_clock),
    .reset(aes_invcipher_op1_reset),
    .io_input_valid(aes_invcipher_op1_io_input_valid),
    .io_input_text(aes_invcipher_op1_io_input_text),
    .io_output_text(aes_invcipher_op1_io_output_text),
    .io_output_valid(aes_invcipher_op1_io_output_valid)
  );
  AESDecrypt_1 aes_invcipher_op2 ( // @[SE.scala 175:39]
    .clock(aes_invcipher_op2_clock),
    .reset(aes_invcipher_op2_reset),
    .io_input_valid(aes_invcipher_op2_io_input_valid),
    .io_input_text(aes_invcipher_op2_io_input_text),
    .io_output_text(aes_invcipher_op2_io_output_text),
    .io_output_valid(aes_invcipher_op2_io_output_valid)
  );
  AESEncrypt256 aes_cipher ( // @[SE.scala 182:57]
    .clock(aes_cipher_clock),
    .reset(aes_cipher_reset),
    .io_input_valid(aes_cipher_io_input_valid),
    .io_input_op1(aes_cipher_io_input_op1),
    .io_input_op2(aes_cipher_io_input_op2),
    .io_output_text(aes_cipher_io_output_text),
    .io_output_valid(aes_cipher_io_output_valid)
  );
  AESEncrypt aes_cipher_for_hash_C ( // @[SE.scala 185:49]
    .clock(aes_cipher_for_hash_C_clock),
    .reset(aes_cipher_for_hash_C_reset),
    .io_input_valid(aes_cipher_for_hash_C_io_input_valid),
    .io_input_text(aes_cipher_for_hash_C_io_input_text),
    .io_output_text(aes_cipher_for_hash_C_io_output_text),
    .io_output_valid(aes_cipher_for_hash_C_io_output_valid)
  );
  AESEncrypt aes_cipher_for_op1 ( // @[SE.scala 186:49]
    .clock(aes_cipher_for_op1_clock),
    .reset(aes_cipher_for_op1_reset),
    .io_input_valid(aes_cipher_for_op1_io_input_valid),
    .io_input_text(aes_cipher_for_op1_io_input_text),
    .io_output_text(aes_cipher_for_op1_io_output_text),
    .io_output_valid(aes_cipher_for_op1_io_output_valid)
  );
  AESEncrypt aes_cipher_for_op2 ( // @[SE.scala 187:49]
    .clock(aes_cipher_for_op2_clock),
    .reset(aes_cipher_for_op2_reset),
    .io_input_valid(aes_cipher_for_op2_io_input_valid),
    .io_input_text(aes_cipher_for_op2_io_input_text),
    .io_output_text(aes_cipher_for_op2_io_output_text),
    .io_output_valid(aes_cipher_for_op2_io_output_valid)
  );
  AESEncrypt aes_cipher_for_pub_var ( // @[SE.scala 188:44]
    .clock(aes_cipher_for_pub_var_clock),
    .reset(aes_cipher_for_pub_var_reset),
    .io_input_valid(aes_cipher_for_pub_var_io_input_valid),
    .io_input_text(aes_cipher_for_pub_var_io_input_text),
    .io_output_text(aes_cipher_for_pub_var_io_output_text),
    .io_output_valid(aes_cipher_for_pub_var_io_output_valid)
  );
  Plaintext_Reverse_Connector PRC_0 ( // @[SE.scala 211:23]
    .io_op1(PRC_0_io_op1),
    .io_op2(PRC_0_io_op2),
    .io_inst(PRC_0_io_inst),
    .io_out_0(PRC_0_io_out_0),
    .io_out_1(PRC_0_io_out_1),
    .io_out_2(PRC_0_io_out_2),
    .io_out_3(PRC_0_io_out_3),
    .io_out_4(PRC_0_io_out_4),
    .io_out_5(PRC_0_io_out_5),
    .io_out_6(PRC_0_io_out_6),
    .io_out_7(PRC_0_io_out_7),
    .io_out_8(PRC_0_io_out_8),
    .io_out_9(PRC_0_io_out_9),
    .io_out_10(PRC_0_io_out_10),
    .io_out_11(PRC_0_io_out_11),
    .io_out_12(PRC_0_io_out_12),
    .io_out_13(PRC_0_io_out_13),
    .io_out_14(PRC_0_io_out_14),
    .io_out_15(PRC_0_io_out_15)
  );
  Hash_Compare HC_op1 ( // @[SE.scala 214:28]
    .io_hash_orig(HC_op1_io_hash_orig),
    .io_hash_regenerated(HC_op1_io_hash_regenerated),
    .io_valid_in(HC_op1_io_valid_in),
    .io_valid_out(HC_op1_io_valid_out),
    .io_compare_result(HC_op1_io_compare_result)
  );
  Hash_Compare HC_op2 ( // @[SE.scala 215:28]
    .io_hash_orig(HC_op2_io_hash_orig),
    .io_hash_regenerated(HC_op2_io_hash_regenerated),
    .io_valid_in(HC_op2_io_valid_in),
    .io_valid_out(HC_op2_io_valid_out),
    .io_compare_result(HC_op2_io_compare_result)
  );
  Version_ID_Generator VID_0 ( // @[SE.scala 219:27]
    .io_pub_priv_opA(VID_0_io_pub_priv_opA),
    .io_pub_priv_opB(VID_0_io_pub_priv_opB),
    .io_version_id_opA(VID_0_io_version_id_opA),
    .io_version_id_opB(VID_0_io_version_id_opB),
    .io_valid_in(VID_0_io_valid_in),
    .io_valid_out(VID_0_io_valid_out),
    .io_version_id_out(VID_0_io_version_id_out),
    .io_pub_priv_out(VID_0_io_pub_priv_out)
  );
  moduled_prng g ( // @[SE.scala 246:42]
    .clock(moduled_prng_pub_var_clock),
    .reset(moduled_prng_pub_var_reset),
    .io_increment(moduled_prng_pub_var_io_increment),
    .io_PUB_VAR_HASH_LFSR(moduled_prng_pub_var_io_PUB_VAR_HASH_LFSR)
  );
  MaxPeriodFibonacciLFSR_1 bit47_randnum_prng ( // @[PRNG.scala 91:22]
    .clock(bit47_randnum_prng_clock),
    .reset(bit47_randnum_prng_reset),
    .io_out_0(bit47_randnum_prng_io_out_0),
    .io_out_1(bit47_randnum_prng_io_out_1),
    .io_out_2(bit47_randnum_prng_io_out_2),
    .io_out_3(bit47_randnum_prng_io_out_3),
    .io_out_4(bit47_randnum_prng_io_out_4),
    .io_out_5(bit47_randnum_prng_io_out_5),
    .io_out_6(bit47_randnum_prng_io_out_6),
    .io_out_7(bit47_randnum_prng_io_out_7),
    .io_out_8(bit47_randnum_prng_io_out_8),
    .io_out_9(bit47_randnum_prng_io_out_9),
    .io_out_10(bit47_randnum_prng_io_out_10),
    .io_out_11(bit47_randnum_prng_io_out_11),
    .io_out_12(bit47_randnum_prng_io_out_12),
    .io_out_13(bit47_randnum_prng_io_out_13),
    .io_out_14(bit47_randnum_prng_io_out_14),
    .io_out_15(bit47_randnum_prng_io_out_15),
    .io_out_16(bit47_randnum_prng_io_out_16),
    .io_out_17(bit47_randnum_prng_io_out_17),
    .io_out_18(bit47_randnum_prng_io_out_18),
    .io_out_19(bit47_randnum_prng_io_out_19),
    .io_out_20(bit47_randnum_prng_io_out_20),
    .io_out_21(bit47_randnum_prng_io_out_21),
    .io_out_22(bit47_randnum_prng_io_out_22),
    .io_out_23(bit47_randnum_prng_io_out_23),
    .io_out_24(bit47_randnum_prng_io_out_24),
    .io_out_25(bit47_randnum_prng_io_out_25),
    .io_out_26(bit47_randnum_prng_io_out_26),
    .io_out_27(bit47_randnum_prng_io_out_27),
    .io_out_28(bit47_randnum_prng_io_out_28),
    .io_out_29(bit47_randnum_prng_io_out_29),
    .io_out_30(bit47_randnum_prng_io_out_30),
    .io_out_31(bit47_randnum_prng_io_out_31),
    .io_out_32(bit47_randnum_prng_io_out_32),
    .io_out_33(bit47_randnum_prng_io_out_33),
    .io_out_34(bit47_randnum_prng_io_out_34),
    .io_out_35(bit47_randnum_prng_io_out_35),
    .io_out_36(bit47_randnum_prng_io_out_36),
    .io_out_37(bit47_randnum_prng_io_out_37),
    .io_out_38(bit47_randnum_prng_io_out_38),
    .io_out_39(bit47_randnum_prng_io_out_39),
    .io_out_40(bit47_randnum_prng_io_out_40),
    .io_out_41(bit47_randnum_prng_io_out_41),
    .io_out_42(bit47_randnum_prng_io_out_42),
    .io_out_43(bit47_randnum_prng_io_out_43),
    .io_out_44(bit47_randnum_prng_io_out_44),
    .io_out_45(bit47_randnum_prng_io_out_45),
    .io_out_46(bit47_randnum_prng_io_out_46)
  );
  assign io_in_ready = ready_for_input; // @[SE.scala 277:21]
  assign io_out_result = output_buffer; // @[SE.scala 645:41]
  assign io_out_valid = output_valid; // @[SE.scala 643:41]
  assign io_out_op1_hash_compare = hash_compare_result_op1; // @[SE.scala 646:33]
  assign io_out_op2_hash_compare = hash_compare_result_op2; // @[SE.scala 647:33]
  assign seoperation_io_inst = inst_buffer; // @[SE.scala 433:33]
  assign seoperation_io_in_valid = lv2ok_buffer; // @[SE.scala 435:41]
  assign seoperation_io_op1_input = is_enc_var_hash ? pub_var_hash_register : _op1_plaintext_64_T_3; // @[SE.scala 438:46]
  assign seoperation_io_op2_input = decrypted_op2_val_buffer[127:64]; // @[SE.scala 440:50]
  assign aes_invcipher_op1_clock = clock;
  assign aes_invcipher_op1_reset = reset;
  assign aes_invcipher_op1_io_input_valid = lv2_AES_valid; // @[SE.scala 331:57]
  assign aes_invcipher_op1_io_input_text = {ciph_op1_val,ciph_op1_hash}; // @[Cat.scala 31:58]
  assign aes_invcipher_op2_clock = clock;
  assign aes_invcipher_op2_reset = reset;
  assign aes_invcipher_op2_io_input_valid = lv2_AES_valid; // @[SE.scala 334:57]
  assign aes_invcipher_op2_io_input_text = {ciph_op2_val,ciph_op2_hash}; // @[Cat.scala 31:58]
  assign aes_cipher_clock = clock;
  assign aes_cipher_reset = reset;
  assign aes_cipher_io_input_valid = lv4_AES_valid; // @[SE.scala 562:49]
  assign aes_cipher_io_input_op1 = aes_input_reverse_bit[127:0]; // @[SE.scala 544:80]
  assign aes_cipher_io_input_op2 = aes_input_reverse_bit[255:128]; // @[SE.scala 545:80]
  assign aes_cipher_for_hash_C_clock = clock;
  assign aes_cipher_for_hash_C_reset = reset;
  assign aes_cipher_for_hash_C_io_input_valid = lv2_AES_valid; // @[SE.scala 336:57]
  assign aes_cipher_for_hash_C_io_input_text = {aes_cipher_for_hash_C_io_input_text_hi,
    aes_cipher_for_hash_C_io_input_text_lo}; // @[SE.scala 335:96]
  assign aes_cipher_for_op1_clock = clock;
  assign aes_cipher_for_op1_reset = reset;
  assign aes_cipher_for_op1_io_input_valid = lv3_AES_valid; // @[SE.scala 476:57]
  assign aes_cipher_for_op1_io_input_text = decrypted_op1_hash_buffer; // @[SE.scala 475:57]
  assign aes_cipher_for_op2_clock = clock;
  assign aes_cipher_for_op2_reset = reset;
  assign aes_cipher_for_op2_io_input_valid = lv3_AES_valid; // @[SE.scala 479:57]
  assign aes_cipher_for_op2_io_input_text = decrypted_op2_hash_buffer; // @[SE.scala 478:57]
  assign aes_cipher_for_pub_var_clock = clock;
  assign aes_cipher_for_pub_var_reset = reset;
  assign aes_cipher_for_pub_var_io_input_valid = lv1ok_buffer & is_enc_var; // @[SE.scala 243:41]
  assign aes_cipher_for_pub_var_io_input_text = {pub_var_hash_register,op1_buffer[255:192]}; // @[Cat.scala 31:58]
  assign PRC_0_io_op1 = op1_buffer; // @[SE.scala 302:41]
  assign PRC_0_io_op2 = op2_buffer; // @[SE.scala 303:49]
  assign PRC_0_io_inst = inst_buffer; // @[SE.scala 304:47]
  assign HC_op1_io_hash_orig = lv2_op1_buffer[315:256]; // @[SE.scala 569:58]
  assign HC_op1_io_hash_regenerated = opA_pub_priv ? decrypted_op1_hash_buffer[127:68] : op1_rehash_result_bit[127:68]; // @[SE.scala 570:47]
  assign HC_op1_io_valid_in = lv3ok_buffer; // @[SE.scala 571:49]
  assign HC_op2_io_hash_orig = lv2_op2_buffer[315:256]; // @[SE.scala 572:58]
  assign HC_op2_io_hash_regenerated = opB_pub_priv ? decrypted_op2_hash_buffer[127:68] : op2_rehash_result_bit[127:68]; // @[SE.scala 573:47]
  assign HC_op2_io_valid_in = lv3ok_buffer; // @[SE.scala 574:49]
  assign VID_0_io_pub_priv_opA = is_enc_inst | opA_pub_priv; // @[SE.scala 451:39]
  assign VID_0_io_pub_priv_opB = is_enc_inst | opB_pub_priv; // @[SE.scala 452:39]
  assign VID_0_io_version_id_opA = decrypted_op1_val_buffer[15:0]; // @[SE.scala 453:43]
  assign VID_0_io_version_id_opB = decrypted_op2_val_buffer[15:0]; // @[SE.scala 454:43]
  assign VID_0_io_valid_in = lv2ok_buffer; // @[SE.scala 455:41]
  assign moduled_prng_pub_var_clock = clock;
  assign moduled_prng_pub_var_reset = reset;
  assign moduled_prng_pub_var_io_increment = lv1ok_buffer & is_enc_var; // @[SE.scala 243:41]
  assign bit47_randnum_prng_clock = clock;
  assign bit47_randnum_prng_reset = reset;
  always @(posedge clock) begin
    if (io_in_valid) begin // @[Reg.scala 17:18]
      inst_buffer <= io_in_inst; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      op1_buffer <= io_in_op1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      op2_buffer <= io_in_op2; // @[Reg.scala 17:22]
    end
    ready_for_input <= reset | ready_for_input_REG; // @[SE.scala 225:{38,38} 282:49]
    if (reset) begin // @[SE.scala 232:42]
      lv1ok_buffer <= 1'h0; // @[SE.scala 232:42]
    end else begin
      lv1ok_buffer <= lv1ok_buffer_REG; // @[SE.scala 287:41]
    end
    if (reset) begin // @[SE.scala 233:42]
      lv2ok_buffer <= 1'h0; // @[SE.scala 233:42]
    end else begin
      lv2ok_buffer <= lv2ok_buffer_REG; // @[SE.scala 385:41]
    end
    if (reset) begin // @[SE.scala 234:42]
      lv3ok_buffer <= 1'h0; // @[SE.scala 234:42]
    end else begin
      lv3ok_buffer <= lv3ok_buffer_REG; // @[SE.scala 519:41]
    end
    if (reset) begin // @[SE.scala 235:42]
      lv4ok_buffer <= 1'h0; // @[SE.scala 235:42]
    end else begin
      lv4ok_buffer <= lv4ok_buffer_REG; // @[SE.scala 599:41]
    end
    if (aes_cipher_for_pub_var_io_output_valid) begin // @[SE.scala 252:53]
      pub_var_hash_register <= aes_cipher_for_pub_var_io_output_text[127:64]; // @[SE.scala 253:39]
    end
    if (reset) begin // @[SE.scala 272:35]
      output_valid <= 1'h0; // @[SE.scala 272:35]
    end else begin
      output_valid <= _GEN_197;
    end
    if (io_in_valid & io_in_ready) begin // @[SE.scala 281:47]
      ready_for_input_REG <= 1'h0;
    end else begin
      ready_for_input_REG <= io_out_valid & io_out_ready | ready_for_input;
    end
    lv1ok_buffer_REG <= _next_ready_for_input_T | _next_lv1ok_buffer_T_1; // @[SE.scala 286:39]
    if (reset) begin // @[SE.scala 315:42]
      lv2_AES_valid <= 1'h0; // @[SE.scala 315:42]
    end else begin
      lv2_AES_valid <= lv2_AES_valid_REG; // @[SE.scala 325:41]
    end
    if (reset) begin // @[SE.scala 316:58]
      tmp_1 <= 1'h0; // @[SE.scala 316:58]
    end else begin
      tmp_1 <= tmp_1_REG; // @[SE.scala 326:49]
    end
    lv2_AES_valid_REG <= lv1ok_buffer & ~tmp_1 & ~is_enc_inst; // @[SE.scala 323:72]
    tmp_1_REG <= lv1ok_buffer & ~lv2_AES_valid | _next_tmp_1_T_2; // @[SE.scala 324:55]
    if (aes_invcipher_op1_io_output_valid) begin // @[Reg.scala 17:18]
      lv2_op1_buffer <= op1_buffer; // @[Reg.scala 17:22]
    end
    if (aes_invcipher_op1_io_output_valid) begin // @[Reg.scala 17:18]
      lv2_op2_buffer <= op2_buffer; // @[Reg.scala 17:22]
    end
    if (aes_cipher_for_hash_C_io_output_valid) begin // @[Reg.scala 17:18]
      hash_C_original_buffer <= aes_cipher_for_hash_C_io_output_text; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 348:66]
      hash_C_original_buffer_valid <= 1'h0; // @[SE.scala 348:66]
    end else begin
      hash_C_original_buffer_valid <= hash_C_original_buffer_valid_REG; // @[SE.scala 365:49]
    end
    if (aes_invcipher_op1_io_output_valid) begin // @[Reg.scala 17:18]
      decrypted_op1_val_buffer <= aes_invcipher_op1_io_output_text[255:128]; // @[Reg.scala 17:22]
    end
    if (aes_invcipher_op1_io_output_valid) begin // @[Reg.scala 17:18]
      decrypted_op1_hash_buffer <= aes_invcipher_op1_io_output_text[127:0]; // @[Reg.scala 17:22]
    end
    if (aes_invcipher_op2_io_output_valid) begin // @[Reg.scala 17:18]
      decrypted_op2_val_buffer <= aes_invcipher_op2_io_output_text[255:128]; // @[Reg.scala 17:22]
    end
    if (aes_invcipher_op2_io_output_valid) begin // @[Reg.scala 17:18]
      decrypted_op2_hash_buffer <= aes_invcipher_op2_io_output_text[127:0]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 359:42]
      lv3_AES_valid <= 1'h0; // @[SE.scala 359:42]
    end else begin
      lv3_AES_valid <= lv3_AES_valid_REG; // @[SE.scala 393:41]
    end
    if (reset) begin // @[SE.scala 360:58]
      tmp_2 <= 1'h0; // @[SE.scala 360:58]
    end else begin
      tmp_2 <= tmp_2_REG; // @[SE.scala 394:49]
    end
    hash_C_original_buffer_valid_REG <= aes_cipher_for_hash_C_io_output_valid | _next_hash_C_original_buffer_valid_T; // @[SE.scala 364:51]
    lv2ok_buffer_REG <= lv2_bypass | aes_invcipher_op1_io_output_valid & aes_invcipher_op2_io_output_valid &
      aes_cipher_for_hash_C_io_output_valid | _next_lv2ok_buffer_T_3; // @[SE.scala 384:39]
    lv3_AES_valid_REG <= lv2ok_buffer & ~tmp_2; // @[SE.scala 391:62]
    tmp_2_REG <= lv2ok_buffer & ~lv3_AES_valid | _next_tmp_2_T_2; // @[SE.scala 392:55]
    if (VID_0_io_valid_out) begin // @[Reg.scala 17:18]
      verID_C <= VID_0_io_version_id_out; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 458:36]
      verID_C_valid <= 1'h0; // @[SE.scala 458:36]
    end else begin
      verID_C_valid <= verID_C_valid_REG; // @[SE.scala 461:41]
    end
    verID_C_valid_REG <= VID_0_io_valid_out | _next_verID_C_valid_T; // @[SE.scala 460:47]
    if (VID_0_io_valid_out) begin // @[Reg.scala 17:18]
      pub_prv_bit <= VID_0_io_pub_priv_out; // @[Reg.scala 17:22]
    end
    if (_result_buffer_T) begin // @[Reg.scala 17:18]
      if (is_enc_inst) begin // @[SE.scala 473:32]
        result_buffer <= enc_padded_result;
      end else begin
        result_buffer <= non_enc_padded_result;
      end
    end
    if (reset) begin // @[SE.scala 484:66]
      result_valid_buffer <= 1'h0; // @[SE.scala 484:66]
    end else begin
      result_valid_buffer <= result_valid_buffer_REG; // @[SE.scala 514:29]
    end
    if (reset) begin // @[SE.scala 486:66]
      hash_C_buffer_valid <= 1'h0; // @[SE.scala 486:66]
    end else begin
      hash_C_buffer_valid <= hash_C_buffer_valid_REG; // @[SE.scala 509:40]
    end
    if (hash_C_buffer_valid) begin // @[Reg.scala 17:18]
      if (is_enc_inst) begin // @[SE.scala 487:81]
        if (is_enc_var) begin // @[SE.scala 471:25]
          hash_C_buffer <= seoperation_io_result[59:0];
        end else begin
          hash_C_buffer <= moduled_prng_pub_var_io_PUB_VAR_HASH_LFSR[59:0];
        end
      end else begin
        hash_C_buffer <= hash_C_original_buffer[125:66];
      end
    end
    if (reset) begin // @[SE.scala 488:58]
      op1_rehash_result_buffer_valid <= 1'h0; // @[SE.scala 488:58]
    end else begin
      op1_rehash_result_buffer_valid <= op1_rehash_result_buffer_valid_REG; // @[SE.scala 503:65]
    end
    if (aes_cipher_for_op1_io_output_valid) begin // @[Reg.scala 17:18]
      op1_rehash_result_bit <= aes_cipher_for_op1_io_output_text; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 490:58]
      op2_rehash_result_buffer_valid <= 1'h0; // @[SE.scala 490:58]
    end else begin
      op2_rehash_result_buffer_valid <= op2_rehash_result_buffer_valid_REG; // @[SE.scala 504:65]
    end
    if (aes_cipher_for_op2_io_output_valid) begin // @[Reg.scala 17:18]
      op2_rehash_result_bit <= aes_cipher_for_op2_io_output_text; // @[Reg.scala 17:22]
    end
    op1_rehash_result_buffer_valid_REG <= aes_cipher_for_op1_io_output_valid | _next_op1_rehash_result_buffer_valid_T; // @[SE.scala 501:63]
    op2_rehash_result_buffer_valid_REG <= aes_cipher_for_op2_io_output_valid | _next_op2_rehash_result_buffer_valid_T; // @[SE.scala 502:63]
    hash_C_buffer_valid_REG <= hash_C_original_buffer_valid | _next_hash_C_buffer_valid_T; // @[SE.scala 508:46]
    result_valid_buffer_REG <= lv2ok_buffer | _n_result_valid_buffer_T; // @[SE.scala 513:37]
    lv3ok_buffer_REG <= result_valid_buffer & hash_C_buffer_valid & op1_rehash_result_buffer_valid &
      op2_rehash_result_buffer_valid | _next_lv3ok_buffer_T_3; // @[SE.scala 518:39]
    if (reset) begin // @[SE.scala 548:42]
      lv4_AES_valid <= 1'h0; // @[SE.scala 548:42]
    end else begin
      lv4_AES_valid <= lv4_AES_valid_REG; // @[SE.scala 557:41]
    end
    if (reset) begin // @[SE.scala 549:58]
      tmp_3 <= 1'h0; // @[SE.scala 549:58]
    end else begin
      tmp_3 <= tmp_3_REG; // @[SE.scala 558:49]
    end
    lv4_AES_valid_REG <= lv3ok_buffer & ~tmp_3; // @[SE.scala 555:62]
    tmp_3_REG <= lv3ok_buffer & ~lv4_AES_valid | _next_tmp_3_T_2; // @[SE.scala 556:55]
    if (reset) begin // @[SE.scala 584:66]
      output_buffer_enc_valid <= 1'h0; // @[SE.scala 584:66]
    end else begin
      output_buffer_enc_valid <= output_buffer_enc_valid_REG; // @[SE.scala 595:57]
    end
    if (aes_cipher_io_output_valid) begin // @[Reg.scala 17:18]
      output_buffer_enc <= aes_cipher_io_output_text; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 586:74]
      output_buffer <= 316'h0; // @[SE.scala 586:74]
    end else if (compare_hash_total) begin // @[SE.scala 622:34]
      output_buffer <= output_connect; // @[SE.scala 623:31]
    end else begin
      output_buffer <= 316'h0; // @[SE.scala 625:31]
    end
    if (HC_op1_io_valid_out) begin // @[Reg.scala 17:18]
      hash_compare_result_op1 <= _hash_compare_result_op1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 588:58]
      hash_compare_result_op1_valid <= 1'h0; // @[SE.scala 588:58]
    end else begin
      hash_compare_result_op1_valid <= hash_compare_result_op1_valid_REG; // @[SE.scala 612:57]
    end
    if (HC_op2_io_valid_out) begin // @[Reg.scala 17:18]
      hash_compare_result_op2 <= _hash_compare_result_op2_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[SE.scala 590:58]
      hash_compare_result_op2_valid <= 1'h0; // @[SE.scala 590:58]
    end else begin
      hash_compare_result_op2_valid <= hash_compare_result_op2_valid_REG; // @[SE.scala 613:57]
    end
    output_buffer_enc_valid_REG <= aes_cipher_io_output_valid | _next_output_buffer_enc_valid_T; // @[SE.scala 594:54]
    lv4ok_buffer_REG <= output_buffer_enc_valid & hash_compare_result_op1_valid & hash_compare_result_op2_valid |
      _next_lv4ok_buffer_T_2; // @[SE.scala 598:38]
    hash_compare_result_op1_valid_REG <= HC_op1_io_valid_out | _next_hash_compare_result_op1_valid_T; // @[SE.scala 610:63]
    hash_compare_result_op2_valid_REG <= HC_op2_io_valid_out | _next_hash_compare_result_op2_valid_T; // @[SE.scala 611:63]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & ~reset) begin
          $fwrite(32'h80000002,"\tinst_buffer: %x\n",inst_buffer); // @[SE.scala 291:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & _T_8) begin
          $fwrite(32'h80000002,"\top1_buffer: %x\n",op1_buffer); // @[SE.scala 292:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & _T_8) begin
          $fwrite(32'h80000002,"\top2_buffer: %x\n",op2_buffer); // @[SE.scala 293:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & _T_8) begin
          $fwrite(32'h80000002,"\tready_for_input: %x\n",ready_for_input); // @[SE.scala 294:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & _T_8) begin
          $fwrite(32'h80000002,"\tlv1ok_buffer: %x\n",lv1ok_buffer); // @[SE.scala 295:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8) begin
          $fwrite(32'h80000002,"[Stage: Level_1 Buffer -> Level_2 Buffer]\n"); // @[SE.scala 299:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\tconnected_reversed_plaintext_buffer: "); // @[SE.scala 398:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_0); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_1); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_2); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_3); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_4); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_5); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_6); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_7); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_8); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_9); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_10); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_11); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_12); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_13); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_14); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",connected_reversed_plaintext_buffer_15); // @[SE.scala 400:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\n"); // @[SE.scala 402:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\thash_C_original_buffer: %x\n",hash_C_original_buffer); // @[SE.scala 403:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\tdecrypted_op1_val_buffer: %x\n",decrypted_op1_val_buffer); // @[SE.scala 408:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\tdecrypted_op1_hash_buffer: "); // @[SE.scala 409:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[0]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[1]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[2]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[3]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[4]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[5]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[6]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[7]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[8]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[9]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[10]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[11]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[12]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[13]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[14]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op1_hash_buffer[15]); // @[SE.scala 411:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\n"); // @[SE.scala 413:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\tdecrypted_op2_val_buffer: "); // @[SE.scala 414:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[0]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[1]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[2]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[3]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[4]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[5]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[6]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[7]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[8]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[9]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[10]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[11]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[12]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[13]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[14]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_val_buffer[15]); // @[SE.scala 416:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\n"); // @[SE.scala 418:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\tdecrypted_op2_hash_buffer: "); // @[SE.scala 419:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[0]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[1]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[2]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[3]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[4]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[5]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[6]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[7]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[8]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[9]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[10]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[11]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[12]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[13]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[14]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"%x",decrypted_op2_hash_buffer[15]); // @[SE.scala 421:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\n"); // @[SE.scala 423:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22 & _T_8) begin
          $fwrite(32'h80000002,"\tlv2ok_buffer: %x\n",lv2ok_buffer); // @[SE.scala 424:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8) begin
          $fwrite(32'h80000002,"[Stage: Level_2 Buffer -> Level_3 Buffer]\n"); // @[SE.scala 428:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\tresult_buffer: %x %x (<- RdNum, ignore) %x\n",result_buffer[255:192],result_buffer[191
            :128],result_buffer[127:0]); // @[SE.scala 523:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\thash_C_buffer: %x\n",hash_C_buffer); // @[SE.scala 524:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\top1_bit: %x\n",decrypted_op1_val_buffer); // @[SE.scala 525:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\top2_bit: %x\n",decrypted_op2_val_buffer); // @[SE.scala 526:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\tseoperation.io.op1_input: %x\n",seoperation_io_op1_input); // @[SE.scala 527:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\tseoperation.io.op2_input: %x\n",seoperation_io_op2_input); // @[SE.scala 528:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\tSE Computation Result: %x\n",seoperation_io_result); // @[SE.scala 529:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\tRdNum: %x\n",bit47_randnum); // @[SE.scala 530:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\top1_rehash_result_buffer: %x\n",op1_rehash_result_bit); // @[SE.scala 531:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\top2_rehash_result_buffer: %x\n",op2_rehash_result_bit); // @[SE.scala 532:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_224 & _T_8) begin
          $fwrite(32'h80000002,"\tlv3ok_buffer: %x\n",lv3ok_buffer); // @[SE.scala 533:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8) begin
          $fwrite(32'h80000002,"[Stage: Level_3 Buffer -> Level_4 Buffer]\n"); // @[SE.scala 537:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\taes_input_reverse_bit: %x\n",aes_input_reverse_bit); // @[SE.scala 630:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\tcompare_hash_total: %x\n",compare_hash_total); // @[SE.scala 635:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\toutput_connect: %x\n",output_connect); // @[SE.scala 636:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\toutput_buffer: %x\n",output_buffer); // @[SE.scala 637:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\thash_compare_result_op1: %x\n",hash_compare_result_op1); // @[SE.scala 638:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\thash_compare_result_op2: %x\n",hash_compare_result_op2); // @[SE.scala 639:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (lv4ok_buffer & _T_8) begin
          $fwrite(32'h80000002,"\tlv4ok_buffer: %x\n",lv4ok_buffer); // @[SE.scala 640:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_buffer = _RAND_0[7:0];
  _RAND_1 = {10{`RANDOM}};
  op1_buffer = _RAND_1[315:0];
  _RAND_2 = {10{`RANDOM}};
  op2_buffer = _RAND_2[315:0];
  _RAND_3 = {1{`RANDOM}};
  ready_for_input = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lv1ok_buffer = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lv2ok_buffer = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lv3ok_buffer = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lv4ok_buffer = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  pub_var_hash_register = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  output_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ready_for_input_REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lv1ok_buffer_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lv2_AES_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  tmp_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lv2_AES_valid_REG = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  tmp_1_REG = _RAND_15[0:0];
  _RAND_16 = {10{`RANDOM}};
  lv2_op1_buffer = _RAND_16[315:0];
  _RAND_17 = {10{`RANDOM}};
  lv2_op2_buffer = _RAND_17[315:0];
  _RAND_18 = {4{`RANDOM}};
  hash_C_original_buffer = _RAND_18[127:0];
  _RAND_19 = {1{`RANDOM}};
  hash_C_original_buffer_valid = _RAND_19[0:0];
  _RAND_20 = {4{`RANDOM}};
  decrypted_op1_val_buffer = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  decrypted_op1_hash_buffer = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  decrypted_op2_val_buffer = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  decrypted_op2_hash_buffer = _RAND_23[127:0];
  _RAND_24 = {1{`RANDOM}};
  lv3_AES_valid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tmp_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  hash_C_original_buffer_valid_REG = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lv2ok_buffer_REG = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lv3_AES_valid_REG = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  tmp_2_REG = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  verID_C = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  verID_C_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  verID_C_valid_REG = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  pub_prv_bit = _RAND_33[0:0];
  _RAND_34 = {8{`RANDOM}};
  result_buffer = _RAND_34[255:0];
  _RAND_35 = {1{`RANDOM}};
  result_valid_buffer = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  hash_C_buffer_valid = _RAND_36[0:0];
  _RAND_37 = {2{`RANDOM}};
  hash_C_buffer = _RAND_37[59:0];
  _RAND_38 = {1{`RANDOM}};
  op1_rehash_result_buffer_valid = _RAND_38[0:0];
  _RAND_39 = {4{`RANDOM}};
  op1_rehash_result_bit = _RAND_39[127:0];
  _RAND_40 = {1{`RANDOM}};
  op2_rehash_result_buffer_valid = _RAND_40[0:0];
  _RAND_41 = {4{`RANDOM}};
  op2_rehash_result_bit = _RAND_41[127:0];
  _RAND_42 = {1{`RANDOM}};
  op1_rehash_result_buffer_valid_REG = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  op2_rehash_result_buffer_valid_REG = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  hash_C_buffer_valid_REG = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  result_valid_buffer_REG = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lv3ok_buffer_REG = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lv4_AES_valid = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  tmp_3 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lv4_AES_valid_REG = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  tmp_3_REG = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  output_buffer_enc_valid = _RAND_51[0:0];
  _RAND_52 = {8{`RANDOM}};
  output_buffer_enc = _RAND_52[255:0];
  _RAND_53 = {10{`RANDOM}};
  output_buffer = _RAND_53[315:0];
  _RAND_54 = {1{`RANDOM}};
  hash_compare_result_op1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  hash_compare_result_op1_valid = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  hash_compare_result_op2 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  hash_compare_result_op2_valid = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  output_buffer_enc_valid_REG = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lv4ok_buffer_REG = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  hash_compare_result_op1_valid_REG = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  hash_compare_result_op2_valid_REG = _RAND_61[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
