module FU(
  input   io_A,
  input   io_B,
  output  io_out
);
  wire  _T_2 = io_B; // @[FU.scala 48:29]
  wire  _T_7 = io_A; // @[FU.scala 54:25]
  wire  _T_8 = io_A; // @[FU.scala 54:36]
  wire  _T_11 = _T_8 & _T_2; // @[FU.scala 54:56]
  wire  _T_12 = _T_7 & _T_11; // @[Cat.scala 30:58]
  wire  _GEN_0 = io_A & _T_2 & _T_12; // @[FU.scala 49:41 51:14 54:14]
  wire  _GEN_1 = io_A & _T_2 & _GEN_0; // @[FU.scala 46:35 48:14]
  wire  _T_15 = io_B; // @[FU.scala 59:39]
  wire  _GEN_2 = io_A & io_B & (io_A & io_B); // @[FU.scala 64:43 66:16 69:16]
  wire  _GEN_3 = io_A & io_B & _GEN_2; // @[FU.scala 61:37 63:16]
  wire  _GEN_4 = _T_8 & _T_15 & _GEN_3; // @[FU.scala 57:20 59:16]
  wire  _GEN_5 = io_A & io_B & (io_A & io_B); // @[FU.scala 76:44 78:16 81:16]
  wire  _GEN_6 = io_A & io_B & _GEN_5; // @[FU.scala 73:39 75:16]
  wire  _GEN_7 = _T_8 & _T_15 & (io_A & io_B); // @[FU.scala 84:20 86:14 89:14]
  wire  _GEN_8 = io_A & io_B; // @[FU.scala 92:26 94:14 97:14]
  wire  _GEN_9 = _GEN_8 & io_A; // @[FU.scala 101:14 91:37]
  wire  _GEN_10 = _GEN_7 & _GEN_9; // @[FU.scala 83:35]
  wire  _GEN_11 = _GEN_6 & _GEN_10; // @[FU.scala 72:38]
  wire  _GEN_12 = _GEN_4 & _GEN_11; // @[FU.scala 56:36]
  wire  _GEN_13 = _GEN_1 & _GEN_12; // @[FU.scala 45:30]
  assign io_out = _GEN_13; // @[FU.scala 43:20]
endmodule
module SEOperation(
  input   io_op1_input,
  input   io_op2_input,
  output  io_result
);
  wire  fu_io_A; // @[SEOperation.scala 32:24]
  wire  fu_io_B; // @[SEOperation.scala 32:24]
  wire  fu_io_out; // @[SEOperation.scala 32:24]
  FU fu ( // @[SEOperation.scala 32:24]
    .io_A(fu_io_A),
    .io_B(fu_io_B),
    .io_out(fu_io_out)
  );
  assign io_result = fu_io_out; // @[SEOperation.scala 47:19]
  assign fu_io_A = io_op1_input; // @[SEOperation.scala 41:11]
  assign fu_io_B = io_op2_input; // @[SEOperation.scala 42:11]
endmodule
module AddRoundKey(
  input   io_state_in_0,
  input   io_state_in_1,
  input   io_state_in_2,
  input   io_state_in_3,
  input   io_state_in_4,
  input   io_state_in_5,
  input   io_state_in_6,
  input   io_state_in_7,
  input   io_state_in_8,
  input   io_state_in_9,
  input   io_state_in_10,
  input   io_state_in_11,
  input   io_state_in_12,
  input   io_state_in_13,
  input   io_state_in_14,
  input   io_state_in_15,
  input   io_roundKey_0,
  input   io_roundKey_1,
  input   io_roundKey_2,
  input   io_roundKey_3,
  input   io_roundKey_4,
  input   io_roundKey_5,
  input   io_roundKey_6,
  input   io_roundKey_7,
  input   io_roundKey_8,
  input   io_roundKey_9,
  input   io_roundKey_10,
  input   io_roundKey_11,
  input   io_roundKey_12,
  input   io_roundKey_13,
  input   io_roundKey_14,
  input   io_roundKey_15,
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15
);
  assign io_state_out_0 = io_state_in_0 & io_roundKey_0; // @[AddRoundKey.scala 19:41]
  assign io_state_out_1 = io_state_in_1 & io_roundKey_1; // @[AddRoundKey.scala 19:41]
  assign io_state_out_2 = io_state_in_2 & io_roundKey_2; // @[AddRoundKey.scala 19:41]
  assign io_state_out_3 = io_state_in_3 & io_roundKey_3; // @[AddRoundKey.scala 19:41]
  assign io_state_out_4 = io_state_in_4 & io_roundKey_4; // @[AddRoundKey.scala 19:41]
  assign io_state_out_5 = io_state_in_5 & io_roundKey_5; // @[AddRoundKey.scala 19:41]
  assign io_state_out_6 = io_state_in_6 & io_roundKey_6; // @[AddRoundKey.scala 19:41]
  assign io_state_out_7 = io_state_in_7 & io_roundKey_7; // @[AddRoundKey.scala 19:41]
  assign io_state_out_8 = io_state_in_8 & io_roundKey_8; // @[AddRoundKey.scala 19:41]
  assign io_state_out_9 = io_state_in_9 & io_roundKey_9; // @[AddRoundKey.scala 19:41]
  assign io_state_out_10 = io_state_in_10 & io_roundKey_10; // @[AddRoundKey.scala 19:41]
  assign io_state_out_11 = io_state_in_11 & io_roundKey_11; // @[AddRoundKey.scala 19:41]
  assign io_state_out_12 = io_state_in_12 & io_roundKey_12; // @[AddRoundKey.scala 19:41]
  assign io_state_out_13 = io_state_in_13 & io_roundKey_13; // @[AddRoundKey.scala 19:41]
  assign io_state_out_14 = io_state_in_14 & io_roundKey_14; // @[AddRoundKey.scala 19:41]
  assign io_state_out_15 = io_state_in_15 & io_roundKey_15; // @[AddRoundKey.scala 19:41]
endmodule
module InvCipherRound(
  input   clock,
  input   io_input_valid,
  input   io_state_in_0,
  input   io_state_in_1,
  input   io_state_in_2,
  input   io_state_in_3,
  input   io_state_in_4,
  input   io_state_in_5,
  input   io_state_in_6,
  input   io_state_in_7,
  input   io_state_in_8,
  input   io_state_in_9,
  input   io_state_in_10,
  input   io_state_in_11,
  input   io_state_in_12,
  input   io_state_in_13,
  input   io_state_in_14,
  input   io_state_in_15,
  input   io_roundKey_0,
  input   io_roundKey_1,
  input   io_roundKey_2,
  input   io_roundKey_3,
  input   io_roundKey_4,
  input   io_roundKey_5,
  input   io_roundKey_6,
  input   io_roundKey_7,
  input   io_roundKey_8,
  input   io_roundKey_9,
  input   io_roundKey_10,
  input   io_roundKey_11,
  input   io_roundKey_12,
  input   io_roundKey_13,
  input   io_roundKey_14,
  input   io_roundKey_15,
  output  io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  AddRoundKey_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_15; // @[AddRoundKey.scala 25:62]
  reg  r_1; // @[Reg.scala 15:16]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKey_io_state_in_0),
    .io_state_in_1(AddRoundKey_io_state_in_1),
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_state_in_3(AddRoundKey_io_state_in_3),
    .io_state_in_4(AddRoundKey_io_state_in_4),
    .io_state_in_5(AddRoundKey_io_state_in_5),
    .io_state_in_6(AddRoundKey_io_state_in_6),
    .io_state_in_7(AddRoundKey_io_state_in_7),
    .io_state_in_8(AddRoundKey_io_state_in_8),
    .io_state_in_9(AddRoundKey_io_state_in_9),
    .io_state_in_10(AddRoundKey_io_state_in_10),
    .io_state_in_11(AddRoundKey_io_state_in_11),
    .io_state_in_12(AddRoundKey_io_state_in_12),
    .io_state_in_13(AddRoundKey_io_state_in_13),
    .io_state_in_14(AddRoundKey_io_state_in_14),
    .io_state_in_15(AddRoundKey_io_state_in_15),
    .io_roundKey_0(AddRoundKey_io_roundKey_0),
    .io_roundKey_1(AddRoundKey_io_roundKey_1),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_roundKey_3(AddRoundKey_io_roundKey_3),
    .io_roundKey_4(AddRoundKey_io_roundKey_4),
    .io_roundKey_5(AddRoundKey_io_roundKey_5),
    .io_roundKey_6(AddRoundKey_io_roundKey_6),
    .io_roundKey_7(AddRoundKey_io_roundKey_7),
    .io_roundKey_8(AddRoundKey_io_roundKey_8),
    .io_roundKey_9(AddRoundKey_io_roundKey_9),
    .io_roundKey_10(AddRoundKey_io_roundKey_10),
    .io_roundKey_11(AddRoundKey_io_roundKey_11),
    .io_roundKey_12(AddRoundKey_io_roundKey_12),
    .io_roundKey_13(AddRoundKey_io_roundKey_13),
    .io_roundKey_14(AddRoundKey_io_roundKey_14),
    .io_roundKey_15(AddRoundKey_io_roundKey_15),
    .io_state_out_0(AddRoundKey_io_state_out_0),
    .io_state_out_1(AddRoundKey_io_state_out_1),
    .io_state_out_2(AddRoundKey_io_state_out_2),
    .io_state_out_3(AddRoundKey_io_state_out_3),
    .io_state_out_4(AddRoundKey_io_state_out_4),
    .io_state_out_5(AddRoundKey_io_state_out_5),
    .io_state_out_6(AddRoundKey_io_state_out_6),
    .io_state_out_7(AddRoundKey_io_state_out_7),
    .io_state_out_8(AddRoundKey_io_state_out_8),
    .io_state_out_9(AddRoundKey_io_state_out_9),
    .io_state_out_10(AddRoundKey_io_state_out_10),
    .io_state_out_11(AddRoundKey_io_state_out_11),
    .io_state_out_12(AddRoundKey_io_state_out_12),
    .io_state_out_13(AddRoundKey_io_state_out_13),
    .io_state_out_14(AddRoundKey_io_state_out_14),
    .io_state_out_15(AddRoundKey_io_state_out_15)
  );
  assign io_output_valid = r_1; // @[InvCipherRound.scala 38:21]
  assign AddRoundKey_io_state_in_0 = io_state_in_0 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_1 = io_state_in_1 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_2 = io_state_in_2 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_3 = io_state_in_3 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_4 = io_state_in_4 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_5 = io_state_in_5 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_6 = io_state_in_6 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_7 = io_state_in_7 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_8 = io_state_in_8 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_9 = io_state_in_9 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_10 = io_state_in_10 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_11 = io_state_in_11 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_12 = io_state_in_12 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_13 = io_state_in_13 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_14 = io_state_in_14 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_state_in_15 = io_state_in_15 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_roundKey_0 = io_roundKey_0 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_1 = io_roundKey_1 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_2 = io_roundKey_2 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_3 = io_roundKey_3 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_4 = io_roundKey_4 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_5 = io_roundKey_5 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_6 = io_roundKey_6 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_7 = io_roundKey_7 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_8 = io_roundKey_8 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_9 = io_roundKey_9 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_10 = io_roundKey_10 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_11 = io_roundKey_11 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_12 = io_roundKey_12 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_13 = io_roundKey_13 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_14 = io_roundKey_14 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  assign AddRoundKey_io_roundKey_15 = io_roundKey_15 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
  always @(posedge clock) begin
    r_1 <= io_input_valid; // @[Reg.scala 15:16 16:{19,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_1 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InvSubBytes(
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15
);
  wire  _GEN_30 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_60 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_30))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_90 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_60))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_120 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_90))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_150 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_120))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_180 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_150))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_210 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_180))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_240 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_210))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_286 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_316 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_286))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_346 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_316))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_376 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_346))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_406 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_376))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_436 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_406))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_466 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_436))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_496 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_466))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_542 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_572 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_542))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_602 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_572))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_632 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_602))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_662 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_632))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_692 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_662))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_722 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_692))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_752 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_722))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_798 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_828 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_798))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_858 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_828))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_888 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_858))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_918 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_888))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_948 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_918))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_978 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_948))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1008 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_978))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1054 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1084 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1054))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1114 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1084))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1144 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1114))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1174 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1144))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1204 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1174))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1234 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1204))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1264 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1234))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1310 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1340 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1310))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1370 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1340))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1400 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1370))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1430 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1400))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1460 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1430))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1490 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1460))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1520 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1490))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1566 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1596 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1566))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1626 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1596))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1656 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1626))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1686 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1656))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1716 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1686))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1746 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1716))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1776 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1746))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1822 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1852 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1822))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1882 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1852))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1912 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1882))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1942 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1912))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_1972 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1942))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2002 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1972))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2032 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2002))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2078 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2108 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2078))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2138 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2108))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2168 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2138))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2198 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2168))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2228 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2198))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2258 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2228))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2288 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2258))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2334 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2364 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2334))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2394 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2364))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2424 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2394))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2454 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2424))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2484 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2454))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2514 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2484))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2544 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2514))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2590 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2620 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2590))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2650 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2620))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2680 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2650))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2710 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2680))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2740 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2710))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2770 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2740))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2800 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2770))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2846 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2876 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2846))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2906 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2876))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2936 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2906))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2966 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2936))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_2996 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2966))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3026 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2996))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3056 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3026))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3102 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3132 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3102))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3162 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3132))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3192 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3162))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3222 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3192))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3252 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3222))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3282 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3252))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3312 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3282))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3358 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3388 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3358))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3418 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3388))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3448 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3418))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3478 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3448))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3508 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3478))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3538 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3508))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3568 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3538))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3614 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3644 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3614))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3674 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3644))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3704 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3674))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3734 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3704))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3764 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3734))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3794 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3764))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3824 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3794))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3870 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3900 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3870))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3930 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3900))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3960 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3930))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_3990 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3960))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_4020 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3990))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_4050 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4020))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_4080 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4050))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_0 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_240)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_1 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_496)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_2 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_752)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_3 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1008)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_4 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1264)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_5 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1520)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_6 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1776)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_7 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2032)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_8 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2288)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_9 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2544)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_10 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2800)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_11 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3056)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_12 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3312)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_13 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3568)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_14 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3824)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_15 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_4080)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
endmodule
module InvCipherRound_3(
  input   clock,
  input   io_input_valid,
  input   io_roundKey_0,
  input   io_roundKey_1,
  input   io_roundKey_2,
  input   io_roundKey_3,
  input   io_roundKey_4,
  input   io_roundKey_5,
  input   io_roundKey_6,
  input   io_roundKey_7,
  input   io_roundKey_8,
  input   io_roundKey_9,
  input   io_roundKey_10,
  input   io_roundKey_11,
  input   io_roundKey_12,
  input   io_roundKey_13,
  input   io_roundKey_14,
  input   io_roundKey_15,
  output  io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  AddRoundKey_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire  InvSubBytes_io_state_out_0; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_1; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_2; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_3; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_4; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_5; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_6; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_7; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_8; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_9; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_10; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_11; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_12; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_13; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_14; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_15; // @[InvSubBytes.scala 43:84]
  reg  r_1; // @[Reg.scala 15:16]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKey_io_state_in_0),
    .io_state_in_1(AddRoundKey_io_state_in_1),
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_state_in_3(AddRoundKey_io_state_in_3),
    .io_state_in_4(AddRoundKey_io_state_in_4),
    .io_state_in_5(AddRoundKey_io_state_in_5),
    .io_state_in_6(AddRoundKey_io_state_in_6),
    .io_state_in_7(AddRoundKey_io_state_in_7),
    .io_state_in_8(AddRoundKey_io_state_in_8),
    .io_state_in_9(AddRoundKey_io_state_in_9),
    .io_state_in_10(AddRoundKey_io_state_in_10),
    .io_state_in_11(AddRoundKey_io_state_in_11),
    .io_state_in_12(AddRoundKey_io_state_in_12),
    .io_state_in_13(AddRoundKey_io_state_in_13),
    .io_state_in_14(AddRoundKey_io_state_in_14),
    .io_state_in_15(AddRoundKey_io_state_in_15),
    .io_roundKey_0(AddRoundKey_io_roundKey_0),
    .io_roundKey_1(AddRoundKey_io_roundKey_1),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_roundKey_3(AddRoundKey_io_roundKey_3),
    .io_roundKey_4(AddRoundKey_io_roundKey_4),
    .io_roundKey_5(AddRoundKey_io_roundKey_5),
    .io_roundKey_6(AddRoundKey_io_roundKey_6),
    .io_roundKey_7(AddRoundKey_io_roundKey_7),
    .io_roundKey_8(AddRoundKey_io_roundKey_8),
    .io_roundKey_9(AddRoundKey_io_roundKey_9),
    .io_roundKey_10(AddRoundKey_io_roundKey_10),
    .io_roundKey_11(AddRoundKey_io_roundKey_11),
    .io_roundKey_12(AddRoundKey_io_roundKey_12),
    .io_roundKey_13(AddRoundKey_io_roundKey_13),
    .io_roundKey_14(AddRoundKey_io_roundKey_14),
    .io_roundKey_15(AddRoundKey_io_roundKey_15),
    .io_state_out_0(AddRoundKey_io_state_out_0),
    .io_state_out_1(AddRoundKey_io_state_out_1),
    .io_state_out_2(AddRoundKey_io_state_out_2),
    .io_state_out_3(AddRoundKey_io_state_out_3),
    .io_state_out_4(AddRoundKey_io_state_out_4),
    .io_state_out_5(AddRoundKey_io_state_out_5),
    .io_state_out_6(AddRoundKey_io_state_out_6),
    .io_state_out_7(AddRoundKey_io_state_out_7),
    .io_state_out_8(AddRoundKey_io_state_out_8),
    .io_state_out_9(AddRoundKey_io_state_out_9),
    .io_state_out_10(AddRoundKey_io_state_out_10),
    .io_state_out_11(AddRoundKey_io_state_out_11),
    .io_state_out_12(AddRoundKey_io_state_out_12),
    .io_state_out_13(AddRoundKey_io_state_out_13),
    .io_state_out_14(AddRoundKey_io_state_out_14),
    .io_state_out_15(AddRoundKey_io_state_out_15)
  );
  InvSubBytes InvSubBytes ( // @[InvSubBytes.scala 43:84]
    .io_state_out_0(InvSubBytes_io_state_out_0),
    .io_state_out_1(InvSubBytes_io_state_out_1),
    .io_state_out_2(InvSubBytes_io_state_out_2),
    .io_state_out_3(InvSubBytes_io_state_out_3),
    .io_state_out_4(InvSubBytes_io_state_out_4),
    .io_state_out_5(InvSubBytes_io_state_out_5),
    .io_state_out_6(InvSubBytes_io_state_out_6),
    .io_state_out_7(InvSubBytes_io_state_out_7),
    .io_state_out_8(InvSubBytes_io_state_out_8),
    .io_state_out_9(InvSubBytes_io_state_out_9),
    .io_state_out_10(InvSubBytes_io_state_out_10),
    .io_state_out_11(InvSubBytes_io_state_out_11),
    .io_state_out_12(InvSubBytes_io_state_out_12),
    .io_state_out_13(InvSubBytes_io_state_out_13),
    .io_state_out_14(InvSubBytes_io_state_out_14),
    .io_state_out_15(InvSubBytes_io_state_out_15)
  );
  assign io_output_valid = r_1; // @[InvCipherRound.scala 89:21]
  assign AddRoundKey_io_state_in_0 = InvSubBytes_io_state_out_0; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_1 = InvSubBytes_io_state_out_1; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_2 = InvSubBytes_io_state_out_2; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_3 = InvSubBytes_io_state_out_3; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_4 = InvSubBytes_io_state_out_4; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_5 = InvSubBytes_io_state_out_5; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_6 = InvSubBytes_io_state_out_6; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_7 = InvSubBytes_io_state_out_7; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_8 = InvSubBytes_io_state_out_8; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_9 = InvSubBytes_io_state_out_9; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_10 = InvSubBytes_io_state_out_10; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_11 = InvSubBytes_io_state_out_11; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_12 = InvSubBytes_io_state_out_12; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_13 = InvSubBytes_io_state_out_13; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_14 = InvSubBytes_io_state_out_14; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_state_in_15 = InvSubBytes_io_state_out_15; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_roundKey_0 = io_roundKey_0 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_1 = io_roundKey_1 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_2 = io_roundKey_2 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_3 = io_roundKey_3 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_4 = io_roundKey_4 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_5 = io_roundKey_5 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_6 = io_roundKey_6 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_7 = io_roundKey_7 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_8 = io_roundKey_8 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_9 = io_roundKey_9 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_10 = io_roundKey_10 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_11 = io_roundKey_11 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_12 = io_roundKey_12 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_13 = io_roundKey_13 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_14 = io_roundKey_14 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_15 = io_roundKey_15 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
  always @(posedge clock) begin
    r_1 <= io_input_valid; // @[Reg.scala 15:16 16:{19,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_1 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InvCipherRound_30(
  input   clock,
  input   io_input_valid,
  output  io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  AddRoundKey_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire  InvSubBytes_io_state_out_0; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_1; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_2; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_3; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_4; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_5; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_6; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_7; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_8; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_9; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_10; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_11; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_12; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_13; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_14; // @[InvSubBytes.scala 43:84]
  wire  InvSubBytes_io_state_out_15; // @[InvSubBytes.scala 43:84]
  reg  r_1; // @[Reg.scala 15:16]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKey_io_state_in_0),
    .io_state_in_1(AddRoundKey_io_state_in_1),
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_state_in_3(AddRoundKey_io_state_in_3),
    .io_state_in_4(AddRoundKey_io_state_in_4),
    .io_state_in_5(AddRoundKey_io_state_in_5),
    .io_state_in_6(AddRoundKey_io_state_in_6),
    .io_state_in_7(AddRoundKey_io_state_in_7),
    .io_state_in_8(AddRoundKey_io_state_in_8),
    .io_state_in_9(AddRoundKey_io_state_in_9),
    .io_state_in_10(AddRoundKey_io_state_in_10),
    .io_state_in_11(AddRoundKey_io_state_in_11),
    .io_state_in_12(AddRoundKey_io_state_in_12),
    .io_state_in_13(AddRoundKey_io_state_in_13),
    .io_state_in_14(AddRoundKey_io_state_in_14),
    .io_state_in_15(AddRoundKey_io_state_in_15),
    .io_roundKey_0(AddRoundKey_io_roundKey_0),
    .io_roundKey_1(AddRoundKey_io_roundKey_1),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_roundKey_3(AddRoundKey_io_roundKey_3),
    .io_roundKey_4(AddRoundKey_io_roundKey_4),
    .io_roundKey_5(AddRoundKey_io_roundKey_5),
    .io_roundKey_6(AddRoundKey_io_roundKey_6),
    .io_roundKey_7(AddRoundKey_io_roundKey_7),
    .io_roundKey_8(AddRoundKey_io_roundKey_8),
    .io_roundKey_9(AddRoundKey_io_roundKey_9),
    .io_roundKey_10(AddRoundKey_io_roundKey_10),
    .io_roundKey_11(AddRoundKey_io_roundKey_11),
    .io_roundKey_12(AddRoundKey_io_roundKey_12),
    .io_roundKey_13(AddRoundKey_io_roundKey_13),
    .io_roundKey_14(AddRoundKey_io_roundKey_14),
    .io_roundKey_15(AddRoundKey_io_roundKey_15),
    .io_state_out_0(AddRoundKey_io_state_out_0),
    .io_state_out_1(AddRoundKey_io_state_out_1),
    .io_state_out_2(AddRoundKey_io_state_out_2),
    .io_state_out_3(AddRoundKey_io_state_out_3),
    .io_state_out_4(AddRoundKey_io_state_out_4),
    .io_state_out_5(AddRoundKey_io_state_out_5),
    .io_state_out_6(AddRoundKey_io_state_out_6),
    .io_state_out_7(AddRoundKey_io_state_out_7),
    .io_state_out_8(AddRoundKey_io_state_out_8),
    .io_state_out_9(AddRoundKey_io_state_out_9),
    .io_state_out_10(AddRoundKey_io_state_out_10),
    .io_state_out_11(AddRoundKey_io_state_out_11),
    .io_state_out_12(AddRoundKey_io_state_out_12),
    .io_state_out_13(AddRoundKey_io_state_out_13),
    .io_state_out_14(AddRoundKey_io_state_out_14),
    .io_state_out_15(AddRoundKey_io_state_out_15)
  );
  InvSubBytes InvSubBytes ( // @[InvSubBytes.scala 43:84]
    .io_state_out_0(InvSubBytes_io_state_out_0),
    .io_state_out_1(InvSubBytes_io_state_out_1),
    .io_state_out_2(InvSubBytes_io_state_out_2),
    .io_state_out_3(InvSubBytes_io_state_out_3),
    .io_state_out_4(InvSubBytes_io_state_out_4),
    .io_state_out_5(InvSubBytes_io_state_out_5),
    .io_state_out_6(InvSubBytes_io_state_out_6),
    .io_state_out_7(InvSubBytes_io_state_out_7),
    .io_state_out_8(InvSubBytes_io_state_out_8),
    .io_state_out_9(InvSubBytes_io_state_out_9),
    .io_state_out_10(InvSubBytes_io_state_out_10),
    .io_state_out_11(InvSubBytes_io_state_out_11),
    .io_state_out_12(InvSubBytes_io_state_out_12),
    .io_state_out_13(InvSubBytes_io_state_out_13),
    .io_state_out_14(InvSubBytes_io_state_out_14),
    .io_state_out_15(InvSubBytes_io_state_out_15)
  );
  assign io_output_valid = r_1; // @[InvCipherRound.scala 62:21]
  assign AddRoundKey_io_state_in_0 = InvSubBytes_io_state_out_0; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_1 = InvSubBytes_io_state_out_1; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_2 = InvSubBytes_io_state_out_2; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_3 = InvSubBytes_io_state_out_3; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_4 = InvSubBytes_io_state_out_4; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_5 = InvSubBytes_io_state_out_5; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_6 = InvSubBytes_io_state_out_6; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_7 = InvSubBytes_io_state_out_7; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_8 = InvSubBytes_io_state_out_8; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_9 = InvSubBytes_io_state_out_9; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_10 = InvSubBytes_io_state_out_10; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_11 = InvSubBytes_io_state_out_11; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_12 = InvSubBytes_io_state_out_12; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_13 = InvSubBytes_io_state_out_13; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_14 = InvSubBytes_io_state_out_14; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_15 = InvSubBytes_io_state_out_15; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_roundKey_0 = 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_1 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_2 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_3 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_4 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_5 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_6 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_7 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_8 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_9 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_10 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_11 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_12 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_13 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_14 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_15 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
  always @(posedge clock) begin
    r_1 <= io_input_valid; // @[Reg.scala 15:16 16:{19,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_1 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AESDecrypt(
  input   clock,
  input   io_input_valid,
  input   io_input_op1_0,
  input   io_input_op1_1,
  input   io_input_op1_2,
  input   io_input_op1_3,
  input   io_input_op1_4,
  input   io_input_op1_5,
  input   io_input_op1_6,
  input   io_input_op1_7,
  input   io_input_op1_8,
  input   io_input_op1_9,
  input   io_input_op1_10,
  input   io_input_op1_11,
  input   io_input_op1_12,
  input   io_input_op1_13,
  input   io_input_op1_14,
  input   io_input_op1_15,
  input   io_input_op2_0,
  input   io_input_op2_1,
  input   io_input_op2_2,
  input   io_input_op2_3,
  input   io_input_op2_4,
  input   io_input_op2_5,
  input   io_input_op2_6,
  input   io_input_op2_7,
  input   io_input_op2_8,
  input   io_input_op2_9,
  input   io_input_op2_10,
  input   io_input_op2_11,
  input   io_input_op2_12,
  input   io_input_op2_13,
  input   io_input_op2_14,
  input   io_input_op2_15,
  input   io_input_cond_0,
  input   io_input_cond_1,
  input   io_input_cond_2,
  input   io_input_cond_3,
  input   io_input_cond_4,
  input   io_input_cond_5,
  input   io_input_cond_6,
  input   io_input_cond_7,
  input   io_input_cond_8,
  input   io_input_cond_9,
  input   io_input_cond_10,
  input   io_input_cond_11,
  input   io_input_cond_12,
  input   io_input_cond_13,
  input   io_input_cond_14,
  input   io_input_cond_15,
  output  io_output_op1_0,
  output  io_output_op1_1,
  output  io_output_op1_2,
  output  io_output_op1_3,
  output  io_output_op1_4,
  output  io_output_op1_5,
  output  io_output_op1_6,
  output  io_output_op1_7,
  output  io_output_op1_8,
  output  io_output_op1_9,
  output  io_output_op1_10,
  output  io_output_op1_11,
  output  io_output_op1_12,
  output  io_output_op1_13,
  output  io_output_op1_14,
  output  io_output_op1_15,
  output  io_output_op2_0,
  output  io_output_op2_1,
  output  io_output_op2_2,
  output  io_output_op2_3,
  output  io_output_op2_4,
  output  io_output_op2_5,
  output  io_output_op2_6,
  output  io_output_op2_7,
  output  io_output_op2_8,
  output  io_output_op2_9,
  output  io_output_op2_10,
  output  io_output_op2_11,
  output  io_output_op2_12,
  output  io_output_op2_13,
  output  io_output_op2_14,
  output  io_output_op2_15,
  output  io_output_valid
);
  wire  InvCipherRound_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_state_in_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_0; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_1; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_3; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_4; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_5; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_6; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_7; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_8; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_9; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_10; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_11; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_12; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_13; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_14; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_15; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_30_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_30_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_30_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_31_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_31_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_31_io_output_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_32_clock; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_32_io_input_valid; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_32_io_output_valid; // @[InvCipherRound.scala 96:79]
  InvCipherRound InvCipherRound ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_clock),
    .io_input_valid(InvCipherRound_io_input_valid),
    .io_state_in_0(InvCipherRound_io_state_in_0),
    .io_state_in_1(InvCipherRound_io_state_in_1),
    .io_state_in_2(InvCipherRound_io_state_in_2),
    .io_state_in_3(InvCipherRound_io_state_in_3),
    .io_state_in_4(InvCipherRound_io_state_in_4),
    .io_state_in_5(InvCipherRound_io_state_in_5),
    .io_state_in_6(InvCipherRound_io_state_in_6),
    .io_state_in_7(InvCipherRound_io_state_in_7),
    .io_state_in_8(InvCipherRound_io_state_in_8),
    .io_state_in_9(InvCipherRound_io_state_in_9),
    .io_state_in_10(InvCipherRound_io_state_in_10),
    .io_state_in_11(InvCipherRound_io_state_in_11),
    .io_state_in_12(InvCipherRound_io_state_in_12),
    .io_state_in_13(InvCipherRound_io_state_in_13),
    .io_state_in_14(InvCipherRound_io_state_in_14),
    .io_state_in_15(InvCipherRound_io_state_in_15),
    .io_roundKey_0(InvCipherRound_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_io_roundKey_15),
    .io_output_valid(InvCipherRound_io_output_valid)
  );
  InvCipherRound InvCipherRound_1 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_1_clock),
    .io_input_valid(InvCipherRound_1_io_input_valid),
    .io_state_in_0(InvCipherRound_1_io_state_in_0),
    .io_state_in_1(InvCipherRound_1_io_state_in_1),
    .io_state_in_2(InvCipherRound_1_io_state_in_2),
    .io_state_in_3(InvCipherRound_1_io_state_in_3),
    .io_state_in_4(InvCipherRound_1_io_state_in_4),
    .io_state_in_5(InvCipherRound_1_io_state_in_5),
    .io_state_in_6(InvCipherRound_1_io_state_in_6),
    .io_state_in_7(InvCipherRound_1_io_state_in_7),
    .io_state_in_8(InvCipherRound_1_io_state_in_8),
    .io_state_in_9(InvCipherRound_1_io_state_in_9),
    .io_state_in_10(InvCipherRound_1_io_state_in_10),
    .io_state_in_11(InvCipherRound_1_io_state_in_11),
    .io_state_in_12(InvCipherRound_1_io_state_in_12),
    .io_state_in_13(InvCipherRound_1_io_state_in_13),
    .io_state_in_14(InvCipherRound_1_io_state_in_14),
    .io_state_in_15(InvCipherRound_1_io_state_in_15),
    .io_roundKey_0(InvCipherRound_1_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_1_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_1_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_1_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_1_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_1_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_1_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_1_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_1_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_1_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_1_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_1_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_1_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_1_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_1_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_1_io_roundKey_15),
    .io_output_valid(InvCipherRound_1_io_output_valid)
  );
  InvCipherRound InvCipherRound_2 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_2_clock),
    .io_input_valid(InvCipherRound_2_io_input_valid),
    .io_state_in_0(InvCipherRound_2_io_state_in_0),
    .io_state_in_1(InvCipherRound_2_io_state_in_1),
    .io_state_in_2(InvCipherRound_2_io_state_in_2),
    .io_state_in_3(InvCipherRound_2_io_state_in_3),
    .io_state_in_4(InvCipherRound_2_io_state_in_4),
    .io_state_in_5(InvCipherRound_2_io_state_in_5),
    .io_state_in_6(InvCipherRound_2_io_state_in_6),
    .io_state_in_7(InvCipherRound_2_io_state_in_7),
    .io_state_in_8(InvCipherRound_2_io_state_in_8),
    .io_state_in_9(InvCipherRound_2_io_state_in_9),
    .io_state_in_10(InvCipherRound_2_io_state_in_10),
    .io_state_in_11(InvCipherRound_2_io_state_in_11),
    .io_state_in_12(InvCipherRound_2_io_state_in_12),
    .io_state_in_13(InvCipherRound_2_io_state_in_13),
    .io_state_in_14(InvCipherRound_2_io_state_in_14),
    .io_state_in_15(InvCipherRound_2_io_state_in_15),
    .io_roundKey_0(InvCipherRound_2_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_2_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_2_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_2_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_2_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_2_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_2_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_2_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_2_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_2_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_2_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_2_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_2_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_2_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_2_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_2_io_roundKey_15),
    .io_output_valid(InvCipherRound_2_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_3 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_3_clock),
    .io_input_valid(InvCipherRound_3_io_input_valid),
    .io_roundKey_0(InvCipherRound_3_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_3_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_3_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_3_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_3_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_3_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_3_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_3_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_3_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_3_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_3_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_3_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_3_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_3_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_3_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_3_io_roundKey_15),
    .io_output_valid(InvCipherRound_3_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_4 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_4_clock),
    .io_input_valid(InvCipherRound_4_io_input_valid),
    .io_roundKey_0(InvCipherRound_4_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_4_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_4_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_4_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_4_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_4_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_4_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_4_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_4_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_4_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_4_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_4_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_4_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_4_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_4_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_4_io_roundKey_15),
    .io_output_valid(InvCipherRound_4_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_5 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_5_clock),
    .io_input_valid(InvCipherRound_5_io_input_valid),
    .io_roundKey_0(InvCipherRound_5_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_5_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_5_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_5_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_5_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_5_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_5_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_5_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_5_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_5_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_5_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_5_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_5_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_5_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_5_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_5_io_roundKey_15),
    .io_output_valid(InvCipherRound_5_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_6 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_6_clock),
    .io_input_valid(InvCipherRound_6_io_input_valid),
    .io_roundKey_0(InvCipherRound_6_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_6_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_6_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_6_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_6_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_6_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_6_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_6_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_6_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_6_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_6_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_6_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_6_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_6_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_6_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_6_io_roundKey_15),
    .io_output_valid(InvCipherRound_6_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_7 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_7_clock),
    .io_input_valid(InvCipherRound_7_io_input_valid),
    .io_roundKey_0(InvCipherRound_7_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_7_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_7_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_7_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_7_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_7_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_7_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_7_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_7_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_7_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_7_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_7_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_7_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_7_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_7_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_7_io_roundKey_15),
    .io_output_valid(InvCipherRound_7_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_8 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_8_clock),
    .io_input_valid(InvCipherRound_8_io_input_valid),
    .io_roundKey_0(InvCipherRound_8_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_8_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_8_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_8_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_8_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_8_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_8_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_8_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_8_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_8_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_8_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_8_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_8_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_8_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_8_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_8_io_roundKey_15),
    .io_output_valid(InvCipherRound_8_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_9 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_9_clock),
    .io_input_valid(InvCipherRound_9_io_input_valid),
    .io_roundKey_0(InvCipherRound_9_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_9_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_9_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_9_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_9_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_9_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_9_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_9_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_9_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_9_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_9_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_9_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_9_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_9_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_9_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_9_io_roundKey_15),
    .io_output_valid(InvCipherRound_9_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_10 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_10_clock),
    .io_input_valid(InvCipherRound_10_io_input_valid),
    .io_roundKey_0(InvCipherRound_10_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_10_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_10_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_10_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_10_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_10_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_10_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_10_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_10_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_10_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_10_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_10_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_10_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_10_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_10_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_10_io_roundKey_15),
    .io_output_valid(InvCipherRound_10_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_11 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_11_clock),
    .io_input_valid(InvCipherRound_11_io_input_valid),
    .io_roundKey_0(InvCipherRound_11_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_11_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_11_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_11_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_11_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_11_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_11_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_11_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_11_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_11_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_11_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_11_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_11_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_11_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_11_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_11_io_roundKey_15),
    .io_output_valid(InvCipherRound_11_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_12 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_12_clock),
    .io_input_valid(InvCipherRound_12_io_input_valid),
    .io_roundKey_0(InvCipherRound_12_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_12_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_12_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_12_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_12_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_12_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_12_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_12_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_12_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_12_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_12_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_12_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_12_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_12_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_12_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_12_io_roundKey_15),
    .io_output_valid(InvCipherRound_12_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_13 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_13_clock),
    .io_input_valid(InvCipherRound_13_io_input_valid),
    .io_roundKey_0(InvCipherRound_13_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_13_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_13_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_13_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_13_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_13_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_13_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_13_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_13_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_13_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_13_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_13_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_13_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_13_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_13_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_13_io_roundKey_15),
    .io_output_valid(InvCipherRound_13_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_14 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_14_clock),
    .io_input_valid(InvCipherRound_14_io_input_valid),
    .io_roundKey_0(InvCipherRound_14_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_14_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_14_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_14_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_14_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_14_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_14_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_14_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_14_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_14_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_14_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_14_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_14_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_14_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_14_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_14_io_roundKey_15),
    .io_output_valid(InvCipherRound_14_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_15 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_15_clock),
    .io_input_valid(InvCipherRound_15_io_input_valid),
    .io_roundKey_0(InvCipherRound_15_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_15_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_15_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_15_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_15_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_15_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_15_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_15_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_15_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_15_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_15_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_15_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_15_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_15_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_15_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_15_io_roundKey_15),
    .io_output_valid(InvCipherRound_15_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_16 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_16_clock),
    .io_input_valid(InvCipherRound_16_io_input_valid),
    .io_roundKey_0(InvCipherRound_16_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_16_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_16_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_16_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_16_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_16_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_16_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_16_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_16_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_16_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_16_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_16_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_16_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_16_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_16_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_16_io_roundKey_15),
    .io_output_valid(InvCipherRound_16_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_17 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_17_clock),
    .io_input_valid(InvCipherRound_17_io_input_valid),
    .io_roundKey_0(InvCipherRound_17_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_17_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_17_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_17_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_17_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_17_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_17_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_17_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_17_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_17_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_17_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_17_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_17_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_17_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_17_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_17_io_roundKey_15),
    .io_output_valid(InvCipherRound_17_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_18 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_18_clock),
    .io_input_valid(InvCipherRound_18_io_input_valid),
    .io_roundKey_0(InvCipherRound_18_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_18_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_18_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_18_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_18_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_18_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_18_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_18_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_18_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_18_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_18_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_18_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_18_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_18_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_18_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_18_io_roundKey_15),
    .io_output_valid(InvCipherRound_18_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_19 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_19_clock),
    .io_input_valid(InvCipherRound_19_io_input_valid),
    .io_roundKey_0(InvCipherRound_19_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_19_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_19_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_19_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_19_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_19_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_19_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_19_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_19_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_19_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_19_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_19_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_19_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_19_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_19_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_19_io_roundKey_15),
    .io_output_valid(InvCipherRound_19_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_20 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_20_clock),
    .io_input_valid(InvCipherRound_20_io_input_valid),
    .io_roundKey_0(InvCipherRound_20_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_20_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_20_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_20_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_20_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_20_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_20_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_20_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_20_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_20_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_20_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_20_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_20_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_20_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_20_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_20_io_roundKey_15),
    .io_output_valid(InvCipherRound_20_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_21 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_21_clock),
    .io_input_valid(InvCipherRound_21_io_input_valid),
    .io_roundKey_0(InvCipherRound_21_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_21_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_21_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_21_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_21_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_21_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_21_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_21_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_21_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_21_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_21_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_21_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_21_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_21_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_21_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_21_io_roundKey_15),
    .io_output_valid(InvCipherRound_21_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_22 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_22_clock),
    .io_input_valid(InvCipherRound_22_io_input_valid),
    .io_roundKey_0(InvCipherRound_22_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_22_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_22_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_22_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_22_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_22_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_22_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_22_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_22_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_22_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_22_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_22_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_22_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_22_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_22_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_22_io_roundKey_15),
    .io_output_valid(InvCipherRound_22_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_23 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_23_clock),
    .io_input_valid(InvCipherRound_23_io_input_valid),
    .io_roundKey_0(InvCipherRound_23_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_23_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_23_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_23_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_23_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_23_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_23_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_23_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_23_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_23_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_23_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_23_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_23_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_23_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_23_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_23_io_roundKey_15),
    .io_output_valid(InvCipherRound_23_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_24 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_24_clock),
    .io_input_valid(InvCipherRound_24_io_input_valid),
    .io_roundKey_0(InvCipherRound_24_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_24_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_24_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_24_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_24_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_24_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_24_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_24_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_24_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_24_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_24_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_24_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_24_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_24_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_24_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_24_io_roundKey_15),
    .io_output_valid(InvCipherRound_24_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_25 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_25_clock),
    .io_input_valid(InvCipherRound_25_io_input_valid),
    .io_roundKey_0(InvCipherRound_25_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_25_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_25_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_25_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_25_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_25_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_25_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_25_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_25_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_25_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_25_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_25_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_25_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_25_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_25_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_25_io_roundKey_15),
    .io_output_valid(InvCipherRound_25_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_26 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_26_clock),
    .io_input_valid(InvCipherRound_26_io_input_valid),
    .io_roundKey_0(InvCipherRound_26_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_26_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_26_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_26_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_26_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_26_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_26_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_26_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_26_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_26_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_26_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_26_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_26_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_26_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_26_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_26_io_roundKey_15),
    .io_output_valid(InvCipherRound_26_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_27 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_27_clock),
    .io_input_valid(InvCipherRound_27_io_input_valid),
    .io_roundKey_0(InvCipherRound_27_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_27_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_27_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_27_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_27_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_27_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_27_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_27_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_27_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_27_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_27_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_27_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_27_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_27_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_27_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_27_io_roundKey_15),
    .io_output_valid(InvCipherRound_27_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_28 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_28_clock),
    .io_input_valid(InvCipherRound_28_io_input_valid),
    .io_roundKey_0(InvCipherRound_28_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_28_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_28_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_28_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_28_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_28_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_28_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_28_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_28_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_28_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_28_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_28_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_28_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_28_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_28_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_28_io_roundKey_15),
    .io_output_valid(InvCipherRound_28_io_output_valid)
  );
  InvCipherRound_3 InvCipherRound_29 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_29_clock),
    .io_input_valid(InvCipherRound_29_io_input_valid),
    .io_roundKey_0(InvCipherRound_29_io_roundKey_0),
    .io_roundKey_1(InvCipherRound_29_io_roundKey_1),
    .io_roundKey_2(InvCipherRound_29_io_roundKey_2),
    .io_roundKey_3(InvCipherRound_29_io_roundKey_3),
    .io_roundKey_4(InvCipherRound_29_io_roundKey_4),
    .io_roundKey_5(InvCipherRound_29_io_roundKey_5),
    .io_roundKey_6(InvCipherRound_29_io_roundKey_6),
    .io_roundKey_7(InvCipherRound_29_io_roundKey_7),
    .io_roundKey_8(InvCipherRound_29_io_roundKey_8),
    .io_roundKey_9(InvCipherRound_29_io_roundKey_9),
    .io_roundKey_10(InvCipherRound_29_io_roundKey_10),
    .io_roundKey_11(InvCipherRound_29_io_roundKey_11),
    .io_roundKey_12(InvCipherRound_29_io_roundKey_12),
    .io_roundKey_13(InvCipherRound_29_io_roundKey_13),
    .io_roundKey_14(InvCipherRound_29_io_roundKey_14),
    .io_roundKey_15(InvCipherRound_29_io_roundKey_15),
    .io_output_valid(InvCipherRound_29_io_output_valid)
  );
  InvCipherRound_30 InvCipherRound_30 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_30_clock),
    .io_input_valid(InvCipherRound_30_io_input_valid),
    .io_output_valid(InvCipherRound_30_io_output_valid)
  );
  InvCipherRound_30 InvCipherRound_31 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_31_clock),
    .io_input_valid(InvCipherRound_31_io_input_valid),
    .io_output_valid(InvCipherRound_31_io_output_valid)
  );
  InvCipherRound_30 InvCipherRound_32 ( // @[InvCipherRound.scala 96:79]
    .clock(InvCipherRound_32_clock),
    .io_input_valid(InvCipherRound_32_io_input_valid),
    .io_output_valid(InvCipherRound_32_io_output_valid)
  );
  assign io_output_op1_0 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_1 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_2 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_3 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_4 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_5 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_6 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_7 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_8 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_9 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_10 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_11 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_12 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_13 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_14 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_15 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op2_0 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_1 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_2 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_3 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_4 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_5 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_6 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_7 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_8 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_9 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_10 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_11 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_12 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_13 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_14 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_15 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_valid = InvCipherRound_30_io_output_valid & InvCipherRound_31_io_output_valid &
    InvCipherRound_32_io_output_valid; // @[AESDecrypt.scala 77:99]
  assign InvCipherRound_clock = clock;
  assign InvCipherRound_io_input_valid = io_input_valid; // @[AESDecrypt.scala 42:39]
  assign InvCipherRound_io_state_in_0 = io_input_op1_0; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_1 = io_input_op1_1; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_2 = io_input_op1_2; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_3 = io_input_op1_3; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_4 = io_input_op1_4; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_5 = io_input_op1_5; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_6 = io_input_op1_6; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_7 = io_input_op1_7; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_8 = io_input_op1_8; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_9 = io_input_op1_9; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_10 = io_input_op1_10; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_11 = io_input_op1_11; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_12 = io_input_op1_12; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_13 = io_input_op1_13; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_14 = io_input_op1_14; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_state_in_15 = io_input_op1_15; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_1_clock = clock;
  assign InvCipherRound_1_io_input_valid = io_input_valid; // @[AESDecrypt.scala 46:39]
  assign InvCipherRound_1_io_state_in_0 = io_input_op2_0; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_1 = io_input_op2_1; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_2 = io_input_op2_2; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_3 = io_input_op2_3; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_4 = io_input_op2_4; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_5 = io_input_op2_5; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_6 = io_input_op2_6; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_7 = io_input_op2_7; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_8 = io_input_op2_8; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_9 = io_input_op2_9; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_10 = io_input_op2_10; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_11 = io_input_op2_11; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_12 = io_input_op2_12; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_13 = io_input_op2_13; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_14 = io_input_op2_14; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_state_in_15 = io_input_op2_15; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_1_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_2_clock = clock;
  assign InvCipherRound_2_io_input_valid = io_input_valid; // @[AESDecrypt.scala 50:39]
  assign InvCipherRound_2_io_state_in_0 = io_input_cond_0; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_1 = io_input_cond_1; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_2 = io_input_cond_2; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_3 = io_input_cond_3; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_4 = io_input_cond_4; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_5 = io_input_cond_5; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_6 = io_input_cond_6; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_7 = io_input_cond_7; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_8 = io_input_cond_8; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_9 = io_input_cond_9; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_10 = io_input_cond_10; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_11 = io_input_cond_11; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_12 = io_input_cond_12; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_13 = io_input_cond_13; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_14 = io_input_cond_14; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_state_in_15 = io_input_cond_15; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_2_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_3_clock = clock;
  assign InvCipherRound_3_io_input_valid = InvCipherRound_io_output_valid; // @[AESDecrypt.scala 57:46]
  assign InvCipherRound_3_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_3_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_clock = clock;
  assign InvCipherRound_4_io_input_valid = InvCipherRound_3_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_4_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_clock = clock;
  assign InvCipherRound_5_io_input_valid = InvCipherRound_4_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_5_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_clock = clock;
  assign InvCipherRound_6_io_input_valid = InvCipherRound_5_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_6_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_clock = clock;
  assign InvCipherRound_7_io_input_valid = InvCipherRound_6_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_7_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_clock = clock;
  assign InvCipherRound_8_io_input_valid = InvCipherRound_7_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_8_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_clock = clock;
  assign InvCipherRound_9_io_input_valid = InvCipherRound_8_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_9_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_clock = clock;
  assign InvCipherRound_10_io_input_valid = InvCipherRound_9_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_10_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_clock = clock;
  assign InvCipherRound_11_io_input_valid = InvCipherRound_10_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_11_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_clock = clock;
  assign InvCipherRound_12_io_input_valid = InvCipherRound_1_io_output_valid; // @[AESDecrypt.scala 57:46]
  assign InvCipherRound_12_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_clock = clock;
  assign InvCipherRound_13_io_input_valid = InvCipherRound_12_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_13_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_clock = clock;
  assign InvCipherRound_14_io_input_valid = InvCipherRound_13_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_14_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_clock = clock;
  assign InvCipherRound_15_io_input_valid = InvCipherRound_14_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_15_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_clock = clock;
  assign InvCipherRound_16_io_input_valid = InvCipherRound_15_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_16_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_clock = clock;
  assign InvCipherRound_17_io_input_valid = InvCipherRound_16_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_17_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_clock = clock;
  assign InvCipherRound_18_io_input_valid = InvCipherRound_17_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_18_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_clock = clock;
  assign InvCipherRound_19_io_input_valid = InvCipherRound_18_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_19_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_clock = clock;
  assign InvCipherRound_20_io_input_valid = InvCipherRound_19_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_20_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_clock = clock;
  assign InvCipherRound_21_io_input_valid = InvCipherRound_2_io_output_valid; // @[AESDecrypt.scala 57:46]
  assign InvCipherRound_21_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_clock = clock;
  assign InvCipherRound_22_io_input_valid = InvCipherRound_21_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_22_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_clock = clock;
  assign InvCipherRound_23_io_input_valid = InvCipherRound_22_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_23_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_clock = clock;
  assign InvCipherRound_24_io_input_valid = InvCipherRound_23_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_24_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_clock = clock;
  assign InvCipherRound_25_io_input_valid = InvCipherRound_24_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_25_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_clock = clock;
  assign InvCipherRound_26_io_input_valid = InvCipherRound_25_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_26_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_clock = clock;
  assign InvCipherRound_27_io_input_valid = InvCipherRound_26_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_27_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_clock = clock;
  assign InvCipherRound_28_io_input_valid = InvCipherRound_27_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_28_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_clock = clock;
  assign InvCipherRound_29_io_input_valid = InvCipherRound_28_io_output_valid; // @[AESDecrypt.scala 61:46]
  assign InvCipherRound_29_io_roundKey_0 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_1 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_3 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_4 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_5 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_6 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_7 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_8 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_9 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_10 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_11 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_12 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_13 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_14 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_15 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_30_clock = clock;
  assign InvCipherRound_30_io_input_valid = InvCipherRound_11_io_output_valid; // @[AESDecrypt.scala 69:41]
  assign InvCipherRound_31_clock = clock;
  assign InvCipherRound_31_io_input_valid = InvCipherRound_20_io_output_valid; // @[AESDecrypt.scala 69:41]
  assign InvCipherRound_32_clock = clock;
  assign InvCipherRound_32_io_input_valid = InvCipherRound_29_io_output_valid; // @[AESDecrypt.scala 69:41]
  assign io_output_valid = 1'h0;
endmodule
module SubBytes(
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15
);
  wire  _GEN_30 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_60 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_30))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_90 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_60))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_120 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_90))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_150 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_120))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_180 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_150))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_210 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_180))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_240 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_210))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_286 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_316 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_286))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_346 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_316))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_376 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_346))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_406 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_376))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_436 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_406))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_466 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_436))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_496 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_466))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_542 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_572 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_542))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_602 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_572))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_632 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_602))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_662 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_632))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_692 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_662))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_722 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_692))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_752 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_722))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_798 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_828 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_798))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_858 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_828))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_888 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_858))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_918 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_888))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_948 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_918))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_978 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_948))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1008 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_978))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1054 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1084 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1054))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1114 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1084))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1144 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1114))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1174 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1144))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1204 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1174))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1234 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1204))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1264 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1234))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1310 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1340 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1310))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1370 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1340))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1400 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1370))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1430 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1400))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1460 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1430))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1490 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1460))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1520 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1490))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1566 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1596 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1566))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1626 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1596))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1656 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1626))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1686 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1656))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1716 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1686))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1746 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1716))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1776 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1746))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1822 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1852 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1822))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1882 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1852))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1912 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1882))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1942 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1912))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1972 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1942))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2002 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1972))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2032 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2002))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2078 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2108 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2078))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2138 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2108))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2168 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2138))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2198 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2168))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2228 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2198))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2258 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2228))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2288 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2258))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2334 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2364 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2334))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2394 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2364))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2424 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2394))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2454 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2424))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2484 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2454))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2514 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2484))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2544 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2514))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2590 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2620 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2590))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2650 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2620))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2680 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2650))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2710 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2680))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2740 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2710))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2770 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2740))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2800 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2770))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2846 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2876 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2846))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2906 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2876))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2936 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2906))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2966 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2936))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2996 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2966))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3026 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2996))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3056 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3026))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3102 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3132 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3102))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3162 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3132))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3192 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3162))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3222 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3192))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3252 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3222))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3282 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3252))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3312 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3282))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3358 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3388 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3358))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3418 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3388))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3448 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3418))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3478 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3448))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3508 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3478))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3538 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3508))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3568 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3538))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3614 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3644 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3614))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3674 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3644))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3704 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3674))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3734 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3704))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3764 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3734))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3794 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3764))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3824 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3794))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3870 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3900 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3870))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3930 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3900))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3960 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3930))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_3990 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3960))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_4020 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3990))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_4050 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4020))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_4080 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4050))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_0 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_240)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_1 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_496)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_2 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_752)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_3 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1008)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_4 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1264)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_5 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1520)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_6 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1776)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_7 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2032)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_8 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2288)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_9 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2544)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_10 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2800)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_11 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3056)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_12 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3312)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_13 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3568)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_14 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3824)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_15 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_4080)))))))))))))); // @[SubBytes.scala 35:{23,23}]
endmodule
module ShiftRows(
  input   io_state_in_0,
  input   io_state_in_1,
  input   io_state_in_2,
  input   io_state_in_3,
  input   io_state_in_4,
  input   io_state_in_5,
  input   io_state_in_6,
  input   io_state_in_7,
  input   io_state_in_8,
  input   io_state_in_9,
  input   io_state_in_10,
  input   io_state_in_11,
  input   io_state_in_12,
  input   io_state_in_13,
  input   io_state_in_14,
  input   io_state_in_15,
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15
);
  assign io_state_out_0 = io_state_in_0; // @[ShiftRows.scala 13:19]
  assign io_state_out_1 = io_state_in_5; // @[ShiftRows.scala 14:19]
  assign io_state_out_2 = io_state_in_10; // @[ShiftRows.scala 15:19]
  assign io_state_out_3 = io_state_in_15; // @[ShiftRows.scala 16:19]
  assign io_state_out_4 = io_state_in_4; // @[ShiftRows.scala 18:19]
  assign io_state_out_5 = io_state_in_9; // @[ShiftRows.scala 19:19]
  assign io_state_out_6 = io_state_in_14; // @[ShiftRows.scala 20:19]
  assign io_state_out_7 = io_state_in_3; // @[ShiftRows.scala 21:19]
  assign io_state_out_8 = io_state_in_8; // @[ShiftRows.scala 23:19]
  assign io_state_out_9 = io_state_in_13; // @[ShiftRows.scala 24:19]
  assign io_state_out_10 = io_state_in_2; // @[ShiftRows.scala 25:20]
  assign io_state_out_11 = io_state_in_7; // @[ShiftRows.scala 26:20]
  assign io_state_out_12 = io_state_in_12; // @[ShiftRows.scala 28:20]
  assign io_state_out_13 = io_state_in_1; // @[ShiftRows.scala 29:20]
  assign io_state_out_14 = io_state_in_6; // @[ShiftRows.scala 30:20]
  assign io_state_out_15 = io_state_in_11; // @[ShiftRows.scala 31:20]
endmodule
module MixColumns(
  input   io_state_in_0,
  input   io_state_in_1,
  input   io_state_in_2,
  input   io_state_in_3,
  input   io_state_in_4,
  input   io_state_in_5,
  input   io_state_in_6,
  input   io_state_in_7,
  input   io_state_in_8,
  input   io_state_in_9,
  input   io_state_in_10,
  input   io_state_in_11,
  input   io_state_in_12,
  input   io_state_in_13,
  input   io_state_in_14,
  input   io_state_in_15,
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15
);
  wire  _GEN_30 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_60 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_30))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_90 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_60))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_120 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_90))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_150 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_120))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_180 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_150))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_210 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_180))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_240 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_210))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_286 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_316 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_286))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_346 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_316))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_376 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_346))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_406 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_376))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_436 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_406))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_466 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_436))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_496 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_466))))))))))))))))))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_511 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_496)))))))))))))); // @[MixColumns.scala 125:{41,41}]
  wire  _GEN_542 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_572 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_542))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_602 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_572))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_632 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_602))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_662 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_632))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_692 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_662))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_722 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_692))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_752 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_722))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{34,34}]
  wire  _GEN_798 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_828 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_798))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_858 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_828))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_888 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_858))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_918 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_888))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_948 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_918))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_978 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_948))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_1008 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_978))))))))))))))))))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_1023 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1008)))))))))))))); // @[MixColumns.scala 126:{58,58}]
  wire  _GEN_1054 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1084 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1054))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1114 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1084))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1144 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1114))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1174 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1144))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1204 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1174))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1234 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1204))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1264 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1234))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1310 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1340 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1310))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1370 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1340))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1400 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1370))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1430 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1400))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1460 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1430))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1490 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1460))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1520 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1490))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1535 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1520)))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1566 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1596 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1566))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1626 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1596))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1656 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1626))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1686 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1656))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1716 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1686))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1746 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1716))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1776 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1746))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{41,41}]
  wire  _GEN_1822 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_1852 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1822))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_1882 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1852))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_1912 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1882))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_1942 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1912))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_1972 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1942))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_2002 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1972))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_2032 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2002))))))))))))))))))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_2047 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2032)))))))))))))); // @[MixColumns.scala 128:{75,75}]
  wire  _GEN_2078 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2108 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2078))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2138 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2108))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2168 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2138))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2198 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2168))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2228 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2198))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2258 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2228))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2288 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2258))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2334 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2364 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2334))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2394 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2364))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2424 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2394))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2454 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2424))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2484 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2454))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2514 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2484))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2544 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2514))))))))))))))))))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2559 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2544)))))))))))))); // @[MixColumns.scala 130:{41,41}]
  wire  _GEN_2590 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2620 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2590))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2650 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2620))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2680 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2650))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2710 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2680))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2740 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2710))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2770 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2740))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2800 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2770))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{34,34}]
  wire  _GEN_2846 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_2876 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2846))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_2906 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2876))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_2936 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2906))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_2966 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2936))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_2996 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2966))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_3026 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2996))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_3056 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3026))))))))))))))))))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_3071 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3056)))))))))))))); // @[MixColumns.scala 131:{58,58}]
  wire  _GEN_3102 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3132 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3102))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3162 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3132))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3192 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3162))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3222 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3192))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3252 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3222))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3282 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3252))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3312 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3282))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{51,51}]
  wire  _GEN_3358 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3388 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3358))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3418 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3388))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3448 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3418))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3478 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3448))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3508 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3478))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3538 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3508))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3568 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3538))))))))))))))))))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3583 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3568)))))))))))))); // @[MixColumns.scala 132:{75,75}]
  wire  _GEN_3614 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3644 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3614))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3674 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3644))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3704 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3674))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3734 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3704))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3764 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3734))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3794 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3764))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3824 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3794))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{41,41}]
  wire  _GEN_3870 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_3900 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3870))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_3930 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3900))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_3960 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3930))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_3990 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3960))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_4020 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_3990))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_4050 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4020))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_4080 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4050))))))))))))))))))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_4095 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4080)))))))))))))); // @[MixColumns.scala 133:{75,75}]
  wire  _GEN_4126 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4156 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4126))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4186 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4156))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4216 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4186))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4246 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4216))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4276 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4246))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4306 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4276))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4336 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4306))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4382 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4412 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4382))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4442 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4412))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4472 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4442))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4502 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4472))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4532 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4502))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4562 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4532))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4592 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4562))))))))))))))))))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4607 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4592)))))))))))))); // @[MixColumns.scala 135:{41,41}]
  wire  _GEN_4638 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4668 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4638))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4698 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4668))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4728 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4698))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4758 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4728))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4788 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4758))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4818 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4788))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4848 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4818))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{34,34}]
  wire  _GEN_4894 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_4924 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4894))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_4954 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4924))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_4984 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4954))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_5014 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_4984))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_5044 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5014))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_5074 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5044))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_5104 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5074))))))))))))))))))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_5119 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5104)))))))))))))); // @[MixColumns.scala 136:{58,58}]
  wire  _GEN_5150 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5180 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5150))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5210 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5180))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5240 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5210))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5270 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5240))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5300 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5270))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5330 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5300))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5360 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5330))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{52,52}]
  wire  _GEN_5406 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5436 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5406))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5466 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5436))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5496 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5466))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5526 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5496))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5556 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5526))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5586 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5556))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5616 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5586))))))))))))))))))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5631 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5616)))))))))))))); // @[MixColumns.scala 137:{77,77}]
  wire  _GEN_5662 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5692 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5662))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5722 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5692))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5752 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5722))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5782 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5752))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5812 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5782))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5842 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5812))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5872 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5842))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{42,42}]
  wire  _GEN_5918 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_5948 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5918))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_5978 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5948))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6008 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_5978))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6038 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6008))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6068 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6038))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6098 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6068))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6128 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6098))))))))))))))))))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6143 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6128)))))))))))))); // @[MixColumns.scala 138:{77,77}]
  wire  _GEN_6174 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6204 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6174))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6234 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6204))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6264 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6234))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6294 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6264))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6324 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6294))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6354 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6324))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6384 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6354))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6430 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6460 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6430))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6490 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6460))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6520 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6490))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6550 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6520))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6580 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6550))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6610 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6580))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6640 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6610))))))))))))))))))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6655 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6640)))))))))))))); // @[MixColumns.scala 140:{43,43}]
  wire  _GEN_6686 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6716 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6686))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6746 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6716))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6776 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6746))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6806 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6776))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6836 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6806))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6866 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6836))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6896 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6866))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{36,36}]
  wire  _GEN_6942 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_6972 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6942))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7002 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_6972))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7032 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7002))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7062 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7032))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7092 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7062))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7122 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7092))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7152 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7122))))))))))))))))))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7167 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7152)))))))))))))); // @[MixColumns.scala 141:{61,61}]
  wire  _GEN_7198 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7228 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7198))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7258 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7228))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7288 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7258))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7318 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7288))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7348 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7318))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7378 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7348))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7408 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7378))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{54,54}]
  wire  _GEN_7454 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7484 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7454))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7514 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7484))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7544 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7514))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7574 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7544))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7604 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7574))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7634 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7604))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7664 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7634))))))))))))))))))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7679 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7664)))))))))))))); // @[MixColumns.scala 142:{79,79}]
  wire  _GEN_7710 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7740 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7710))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7770 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7740))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7800 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7770))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7830 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7800))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7860 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7830))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7890 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7860))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7920 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7890))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{43,43}]
  wire  _GEN_7966 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_7996 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7966))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8026 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_7996))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8056 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_8026))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8086 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_8056))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8116 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_8086))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8146 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_8116))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8176 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_8146))))))))))))))))))))))))))))); // @[MixColumns.scala 143:{79,79}]
  wire  _GEN_8191 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_8176)))))))))))))); // @[MixColumns.scala 143:{79,79}]
  assign io_state_out_0 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_240)))))))))))))) & _GEN_511 & io_state_in_2 & io_state_in_3; // @[MixColumns.scala 125:82]
  assign io_state_out_1 = io_state_in_0 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_752))))))))))))))) & _GEN_1023 & io_state_in_3; // @[MixColumns.scala 126:82]
  assign io_state_out_2 = io_state_in_0 & io_state_in_1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_1264))))))))))))))) & _GEN_1535; // @[MixColumns.scala 127:75]
  assign io_state_out_3 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1776)))))))))))))) & io_state_in_1 & io_state_in_2 & _GEN_2047; // @[MixColumns.scala 128:75]
  assign io_state_out_4 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2288)))))))))))))) & _GEN_2559 & io_state_in_6 & io_state_in_7; // @[MixColumns.scala 130:82]
  assign io_state_out_5 = io_state_in_4 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_2800))))))))))))))) & _GEN_3071 & io_state_in_7; // @[MixColumns.scala 131:82]
  assign io_state_out_6 = io_state_in_4 & io_state_in_5 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_3312))))))))))))))) & _GEN_3583; // @[MixColumns.scala 132:75]
  assign io_state_out_7 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_3824)))))))))))))) & io_state_in_5 & io_state_in_6 & _GEN_4095; // @[MixColumns.scala 133:75]
  assign io_state_out_8 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_4336)))))))))))))) & _GEN_4607 & io_state_in_10 & io_state_in_11; // @[MixColumns.scala 135:83]
  assign io_state_out_9 = io_state_in_8 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_4848))))))))))))))) & _GEN_5119 & io_state_in_11; // @[MixColumns.scala 136:83]
  assign io_state_out_10 = io_state_in_8 & io_state_in_9 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_5360))))))))))))))) & _GEN_5631; // @[MixColumns.scala 137:77]
  assign io_state_out_11 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_5872)))))))))))))) & io_state_in_9 & io_state_in_10 & _GEN_6143; // @[MixColumns.scala 138:77]
  assign io_state_out_12 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_6384)))))))))))))) & _GEN_6655 & io_state_in_14 & io_state_in_15; // @[MixColumns.scala 140:86]
  assign io_state_out_13 = io_state_in_12 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_6896))))))))))))))) & _GEN_7167 & io_state_in_15; // @[MixColumns.scala 141:86]
  assign io_state_out_14 = io_state_in_12 & io_state_in_13 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_7408))))))))))))))) & _GEN_7679; // @[MixColumns.scala 142:79]
  assign io_state_out_15 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_7920)))))))))))))) & io_state_in_13 & io_state_in_14 & _GEN_8191; // @[MixColumns.scala 143:79]
endmodule
module CipherRound_1(
  input   clock,
  input   io_input_valid,
  input   io_roundKey_0,
  input   io_roundKey_1,
  input   io_roundKey_2,
  input   io_roundKey_3,
  input   io_roundKey_4,
  input   io_roundKey_5,
  input   io_roundKey_6,
  input   io_roundKey_7,
  input   io_roundKey_8,
  input   io_roundKey_9,
  input   io_roundKey_10,
  input   io_roundKey_11,
  input   io_roundKey_12,
  input   io_roundKey_13,
  input   io_roundKey_14,
  input   io_roundKey_15,
  output  io_state_out_2,
  output  io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  AddRoundKey_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire  SubBytes_io_state_out_0; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_1; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_2; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_3; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_4; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_5; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_6; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_7; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_8; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_9; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_10; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_11; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_12; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_13; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_14; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_15; // @[SubBytes.scala 41:81]
  wire  ShiftRows_io_state_in_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_1; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_2; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_3; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_4; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_5; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_6; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_7; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_8; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_9; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_10; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_11; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_12; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_13; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_14; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_15; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_1; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_2; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_3; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_4; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_5; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_6; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_7; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_8; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_9; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_10; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_11; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_12; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_13; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_14; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_15; // @[ShiftRows.scala 35:34]
  wire  MixColumns_io_state_in_0; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_1; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_2; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_3; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_4; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_5; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_6; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_7; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_8; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_9; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_10; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_11; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_12; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_13; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_14; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_15; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_0; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_1; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_2; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_3; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_4; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_5; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_6; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_7; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_8; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_9; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_10; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_11; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_12; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_13; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_14; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_15; // @[MixColumns.scala 153:61]
  reg  r__2; // @[Reg.scala 15:16]
  reg  r_1; // @[Reg.scala 15:16]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKey_io_state_in_0),
    .io_state_in_1(AddRoundKey_io_state_in_1),
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_state_in_3(AddRoundKey_io_state_in_3),
    .io_state_in_4(AddRoundKey_io_state_in_4),
    .io_state_in_5(AddRoundKey_io_state_in_5),
    .io_state_in_6(AddRoundKey_io_state_in_6),
    .io_state_in_7(AddRoundKey_io_state_in_7),
    .io_state_in_8(AddRoundKey_io_state_in_8),
    .io_state_in_9(AddRoundKey_io_state_in_9),
    .io_state_in_10(AddRoundKey_io_state_in_10),
    .io_state_in_11(AddRoundKey_io_state_in_11),
    .io_state_in_12(AddRoundKey_io_state_in_12),
    .io_state_in_13(AddRoundKey_io_state_in_13),
    .io_state_in_14(AddRoundKey_io_state_in_14),
    .io_state_in_15(AddRoundKey_io_state_in_15),
    .io_roundKey_0(AddRoundKey_io_roundKey_0),
    .io_roundKey_1(AddRoundKey_io_roundKey_1),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_roundKey_3(AddRoundKey_io_roundKey_3),
    .io_roundKey_4(AddRoundKey_io_roundKey_4),
    .io_roundKey_5(AddRoundKey_io_roundKey_5),
    .io_roundKey_6(AddRoundKey_io_roundKey_6),
    .io_roundKey_7(AddRoundKey_io_roundKey_7),
    .io_roundKey_8(AddRoundKey_io_roundKey_8),
    .io_roundKey_9(AddRoundKey_io_roundKey_9),
    .io_roundKey_10(AddRoundKey_io_roundKey_10),
    .io_roundKey_11(AddRoundKey_io_roundKey_11),
    .io_roundKey_12(AddRoundKey_io_roundKey_12),
    .io_roundKey_13(AddRoundKey_io_roundKey_13),
    .io_roundKey_14(AddRoundKey_io_roundKey_14),
    .io_roundKey_15(AddRoundKey_io_roundKey_15),
    .io_state_out_0(AddRoundKey_io_state_out_0),
    .io_state_out_1(AddRoundKey_io_state_out_1),
    .io_state_out_2(AddRoundKey_io_state_out_2),
    .io_state_out_3(AddRoundKey_io_state_out_3),
    .io_state_out_4(AddRoundKey_io_state_out_4),
    .io_state_out_5(AddRoundKey_io_state_out_5),
    .io_state_out_6(AddRoundKey_io_state_out_6),
    .io_state_out_7(AddRoundKey_io_state_out_7),
    .io_state_out_8(AddRoundKey_io_state_out_8),
    .io_state_out_9(AddRoundKey_io_state_out_9),
    .io_state_out_10(AddRoundKey_io_state_out_10),
    .io_state_out_11(AddRoundKey_io_state_out_11),
    .io_state_out_12(AddRoundKey_io_state_out_12),
    .io_state_out_13(AddRoundKey_io_state_out_13),
    .io_state_out_14(AddRoundKey_io_state_out_14),
    .io_state_out_15(AddRoundKey_io_state_out_15)
  );
  SubBytes SubBytes ( // @[SubBytes.scala 41:81]
    .io_state_out_0(SubBytes_io_state_out_0),
    .io_state_out_1(SubBytes_io_state_out_1),
    .io_state_out_2(SubBytes_io_state_out_2),
    .io_state_out_3(SubBytes_io_state_out_3),
    .io_state_out_4(SubBytes_io_state_out_4),
    .io_state_out_5(SubBytes_io_state_out_5),
    .io_state_out_6(SubBytes_io_state_out_6),
    .io_state_out_7(SubBytes_io_state_out_7),
    .io_state_out_8(SubBytes_io_state_out_8),
    .io_state_out_9(SubBytes_io_state_out_9),
    .io_state_out_10(SubBytes_io_state_out_10),
    .io_state_out_11(SubBytes_io_state_out_11),
    .io_state_out_12(SubBytes_io_state_out_12),
    .io_state_out_13(SubBytes_io_state_out_13),
    .io_state_out_14(SubBytes_io_state_out_14),
    .io_state_out_15(SubBytes_io_state_out_15)
  );
  ShiftRows ShiftRows ( // @[ShiftRows.scala 35:34]
    .io_state_in_0(ShiftRows_io_state_in_0),
    .io_state_in_1(ShiftRows_io_state_in_1),
    .io_state_in_2(ShiftRows_io_state_in_2),
    .io_state_in_3(ShiftRows_io_state_in_3),
    .io_state_in_4(ShiftRows_io_state_in_4),
    .io_state_in_5(ShiftRows_io_state_in_5),
    .io_state_in_6(ShiftRows_io_state_in_6),
    .io_state_in_7(ShiftRows_io_state_in_7),
    .io_state_in_8(ShiftRows_io_state_in_8),
    .io_state_in_9(ShiftRows_io_state_in_9),
    .io_state_in_10(ShiftRows_io_state_in_10),
    .io_state_in_11(ShiftRows_io_state_in_11),
    .io_state_in_12(ShiftRows_io_state_in_12),
    .io_state_in_13(ShiftRows_io_state_in_13),
    .io_state_in_14(ShiftRows_io_state_in_14),
    .io_state_in_15(ShiftRows_io_state_in_15),
    .io_state_out_0(ShiftRows_io_state_out_0),
    .io_state_out_1(ShiftRows_io_state_out_1),
    .io_state_out_2(ShiftRows_io_state_out_2),
    .io_state_out_3(ShiftRows_io_state_out_3),
    .io_state_out_4(ShiftRows_io_state_out_4),
    .io_state_out_5(ShiftRows_io_state_out_5),
    .io_state_out_6(ShiftRows_io_state_out_6),
    .io_state_out_7(ShiftRows_io_state_out_7),
    .io_state_out_8(ShiftRows_io_state_out_8),
    .io_state_out_9(ShiftRows_io_state_out_9),
    .io_state_out_10(ShiftRows_io_state_out_10),
    .io_state_out_11(ShiftRows_io_state_out_11),
    .io_state_out_12(ShiftRows_io_state_out_12),
    .io_state_out_13(ShiftRows_io_state_out_13),
    .io_state_out_14(ShiftRows_io_state_out_14),
    .io_state_out_15(ShiftRows_io_state_out_15)
  );
  MixColumns MixColumns ( // @[MixColumns.scala 153:61]
    .io_state_in_0(MixColumns_io_state_in_0),
    .io_state_in_1(MixColumns_io_state_in_1),
    .io_state_in_2(MixColumns_io_state_in_2),
    .io_state_in_3(MixColumns_io_state_in_3),
    .io_state_in_4(MixColumns_io_state_in_4),
    .io_state_in_5(MixColumns_io_state_in_5),
    .io_state_in_6(MixColumns_io_state_in_6),
    .io_state_in_7(MixColumns_io_state_in_7),
    .io_state_in_8(MixColumns_io_state_in_8),
    .io_state_in_9(MixColumns_io_state_in_9),
    .io_state_in_10(MixColumns_io_state_in_10),
    .io_state_in_11(MixColumns_io_state_in_11),
    .io_state_in_12(MixColumns_io_state_in_12),
    .io_state_in_13(MixColumns_io_state_in_13),
    .io_state_in_14(MixColumns_io_state_in_14),
    .io_state_in_15(MixColumns_io_state_in_15),
    .io_state_out_0(MixColumns_io_state_out_0),
    .io_state_out_1(MixColumns_io_state_out_1),
    .io_state_out_2(MixColumns_io_state_out_2),
    .io_state_out_3(MixColumns_io_state_out_3),
    .io_state_out_4(MixColumns_io_state_out_4),
    .io_state_out_5(MixColumns_io_state_out_5),
    .io_state_out_6(MixColumns_io_state_out_6),
    .io_state_out_7(MixColumns_io_state_out_7),
    .io_state_out_8(MixColumns_io_state_out_8),
    .io_state_out_9(MixColumns_io_state_out_9),
    .io_state_out_10(MixColumns_io_state_out_10),
    .io_state_out_11(MixColumns_io_state_out_11),
    .io_state_out_12(MixColumns_io_state_out_12),
    .io_state_out_13(MixColumns_io_state_out_13),
    .io_state_out_14(MixColumns_io_state_out_14),
    .io_state_out_15(MixColumns_io_state_out_15)
  );
  assign io_state_out_2 = r__2; // @[CipherRound.scala 88:18]
  assign io_output_valid = r_1; // @[CipherRound.scala 89:21]
  assign AddRoundKey_io_state_in_0 = MixColumns_io_state_out_0; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_1 = MixColumns_io_state_out_1; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_2 = MixColumns_io_state_out_2; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_3 = MixColumns_io_state_out_3; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_4 = MixColumns_io_state_out_4; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_5 = MixColumns_io_state_out_5; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_6 = MixColumns_io_state_out_6; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_7 = MixColumns_io_state_out_7; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_8 = MixColumns_io_state_out_8; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_9 = MixColumns_io_state_out_9; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_10 = MixColumns_io_state_out_10; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_11 = MixColumns_io_state_out_11; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_12 = MixColumns_io_state_out_12; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_13 = MixColumns_io_state_out_13; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_14 = MixColumns_io_state_out_14; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_state_in_15 = MixColumns_io_state_out_15; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_roundKey_0 = io_roundKey_0 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_1 = io_roundKey_1 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_2 = io_roundKey_2 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_3 = io_roundKey_3 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_4 = io_roundKey_4 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_5 = io_roundKey_5 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_6 = io_roundKey_6 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_7 = io_roundKey_7 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_8 = io_roundKey_8 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_9 = io_roundKey_9 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_10 = io_roundKey_10 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_11 = io_roundKey_11 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_12 = io_roundKey_12 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_13 = io_roundKey_13 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_14 = io_roundKey_14 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign AddRoundKey_io_roundKey_15 = io_roundKey_15 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign ShiftRows_io_state_in_0 = SubBytes_io_state_out_0; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_1 = SubBytes_io_state_out_1; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_2 = SubBytes_io_state_out_2; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_3 = SubBytes_io_state_out_3; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_4 = SubBytes_io_state_out_4; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_5 = SubBytes_io_state_out_5; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_6 = SubBytes_io_state_out_6; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_7 = SubBytes_io_state_out_7; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_8 = SubBytes_io_state_out_8; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_9 = SubBytes_io_state_out_9; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_10 = SubBytes_io_state_out_10; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_11 = SubBytes_io_state_out_11; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_12 = SubBytes_io_state_out_12; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_13 = SubBytes_io_state_out_13; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_14 = SubBytes_io_state_out_14; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_15 = SubBytes_io_state_out_15; // @[CipherRound.scala 81:33]
  assign MixColumns_io_state_in_0 = ShiftRows_io_state_out_0; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_1 = ShiftRows_io_state_out_1; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_2 = ShiftRows_io_state_out_2; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_3 = ShiftRows_io_state_out_3; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_4 = ShiftRows_io_state_out_4; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_5 = ShiftRows_io_state_out_5; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_6 = ShiftRows_io_state_out_6; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_7 = ShiftRows_io_state_out_7; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_8 = ShiftRows_io_state_out_8; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_9 = ShiftRows_io_state_out_9; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_10 = ShiftRows_io_state_out_10; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_11 = ShiftRows_io_state_out_11; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_12 = ShiftRows_io_state_out_12; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_13 = ShiftRows_io_state_out_13; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_14 = ShiftRows_io_state_out_14; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_15 = ShiftRows_io_state_out_15; // @[CipherRound.scala 83:34]
  always @(posedge clock) begin
    r__2 <= AddRoundKey_io_state_out_2; // @[Reg.scala 15:16 16:{19,23}]
    r_1 <= io_input_valid; // @[Reg.scala 15:16 16:{19,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r__2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CipherRound_10(
  input   clock,
  input   io_input_valid,
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15,
  output  io_output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  AddRoundKey_io_state_in_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_in_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_15; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_0; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_1; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_3; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_4; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_5; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_6; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_7; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_8; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_9; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_10; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_11; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_12; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_13; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_14; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_15; // @[AddRoundKey.scala 25:62]
  wire  SubBytes_io_state_out_0; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_1; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_2; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_3; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_4; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_5; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_6; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_7; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_8; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_9; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_10; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_11; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_12; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_13; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_14; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_15; // @[SubBytes.scala 41:81]
  wire  ShiftRows_io_state_in_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_1; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_2; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_3; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_4; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_5; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_6; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_7; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_8; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_9; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_10; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_11; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_12; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_13; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_14; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_15; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_1; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_2; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_3; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_4; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_5; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_6; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_7; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_8; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_9; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_10; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_11; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_12; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_13; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_14; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_15; // @[ShiftRows.scala 35:34]
  reg  r__0; // @[Reg.scala 15:16]
  reg  r__1; // @[Reg.scala 15:16]
  reg  r__2; // @[Reg.scala 15:16]
  reg  r__3; // @[Reg.scala 15:16]
  reg  r__4; // @[Reg.scala 15:16]
  reg  r__5; // @[Reg.scala 15:16]
  reg  r__6; // @[Reg.scala 15:16]
  reg  r__7; // @[Reg.scala 15:16]
  reg  r__8; // @[Reg.scala 15:16]
  reg  r__9; // @[Reg.scala 15:16]
  reg  r__10; // @[Reg.scala 15:16]
  reg  r__11; // @[Reg.scala 15:16]
  reg  r__12; // @[Reg.scala 15:16]
  reg  r__13; // @[Reg.scala 15:16]
  reg  r__14; // @[Reg.scala 15:16]
  reg  r__15; // @[Reg.scala 15:16]
  reg  r_1; // @[Reg.scala 15:16]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_0(AddRoundKey_io_state_in_0),
    .io_state_in_1(AddRoundKey_io_state_in_1),
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_state_in_3(AddRoundKey_io_state_in_3),
    .io_state_in_4(AddRoundKey_io_state_in_4),
    .io_state_in_5(AddRoundKey_io_state_in_5),
    .io_state_in_6(AddRoundKey_io_state_in_6),
    .io_state_in_7(AddRoundKey_io_state_in_7),
    .io_state_in_8(AddRoundKey_io_state_in_8),
    .io_state_in_9(AddRoundKey_io_state_in_9),
    .io_state_in_10(AddRoundKey_io_state_in_10),
    .io_state_in_11(AddRoundKey_io_state_in_11),
    .io_state_in_12(AddRoundKey_io_state_in_12),
    .io_state_in_13(AddRoundKey_io_state_in_13),
    .io_state_in_14(AddRoundKey_io_state_in_14),
    .io_state_in_15(AddRoundKey_io_state_in_15),
    .io_roundKey_0(AddRoundKey_io_roundKey_0),
    .io_roundKey_1(AddRoundKey_io_roundKey_1),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_roundKey_3(AddRoundKey_io_roundKey_3),
    .io_roundKey_4(AddRoundKey_io_roundKey_4),
    .io_roundKey_5(AddRoundKey_io_roundKey_5),
    .io_roundKey_6(AddRoundKey_io_roundKey_6),
    .io_roundKey_7(AddRoundKey_io_roundKey_7),
    .io_roundKey_8(AddRoundKey_io_roundKey_8),
    .io_roundKey_9(AddRoundKey_io_roundKey_9),
    .io_roundKey_10(AddRoundKey_io_roundKey_10),
    .io_roundKey_11(AddRoundKey_io_roundKey_11),
    .io_roundKey_12(AddRoundKey_io_roundKey_12),
    .io_roundKey_13(AddRoundKey_io_roundKey_13),
    .io_roundKey_14(AddRoundKey_io_roundKey_14),
    .io_roundKey_15(AddRoundKey_io_roundKey_15),
    .io_state_out_0(AddRoundKey_io_state_out_0),
    .io_state_out_1(AddRoundKey_io_state_out_1),
    .io_state_out_2(AddRoundKey_io_state_out_2),
    .io_state_out_3(AddRoundKey_io_state_out_3),
    .io_state_out_4(AddRoundKey_io_state_out_4),
    .io_state_out_5(AddRoundKey_io_state_out_5),
    .io_state_out_6(AddRoundKey_io_state_out_6),
    .io_state_out_7(AddRoundKey_io_state_out_7),
    .io_state_out_8(AddRoundKey_io_state_out_8),
    .io_state_out_9(AddRoundKey_io_state_out_9),
    .io_state_out_10(AddRoundKey_io_state_out_10),
    .io_state_out_11(AddRoundKey_io_state_out_11),
    .io_state_out_12(AddRoundKey_io_state_out_12),
    .io_state_out_13(AddRoundKey_io_state_out_13),
    .io_state_out_14(AddRoundKey_io_state_out_14),
    .io_state_out_15(AddRoundKey_io_state_out_15)
  );
  SubBytes SubBytes ( // @[SubBytes.scala 41:81]
    .io_state_out_0(SubBytes_io_state_out_0),
    .io_state_out_1(SubBytes_io_state_out_1),
    .io_state_out_2(SubBytes_io_state_out_2),
    .io_state_out_3(SubBytes_io_state_out_3),
    .io_state_out_4(SubBytes_io_state_out_4),
    .io_state_out_5(SubBytes_io_state_out_5),
    .io_state_out_6(SubBytes_io_state_out_6),
    .io_state_out_7(SubBytes_io_state_out_7),
    .io_state_out_8(SubBytes_io_state_out_8),
    .io_state_out_9(SubBytes_io_state_out_9),
    .io_state_out_10(SubBytes_io_state_out_10),
    .io_state_out_11(SubBytes_io_state_out_11),
    .io_state_out_12(SubBytes_io_state_out_12),
    .io_state_out_13(SubBytes_io_state_out_13),
    .io_state_out_14(SubBytes_io_state_out_14),
    .io_state_out_15(SubBytes_io_state_out_15)
  );
  ShiftRows ShiftRows ( // @[ShiftRows.scala 35:34]
    .io_state_in_0(ShiftRows_io_state_in_0),
    .io_state_in_1(ShiftRows_io_state_in_1),
    .io_state_in_2(ShiftRows_io_state_in_2),
    .io_state_in_3(ShiftRows_io_state_in_3),
    .io_state_in_4(ShiftRows_io_state_in_4),
    .io_state_in_5(ShiftRows_io_state_in_5),
    .io_state_in_6(ShiftRows_io_state_in_6),
    .io_state_in_7(ShiftRows_io_state_in_7),
    .io_state_in_8(ShiftRows_io_state_in_8),
    .io_state_in_9(ShiftRows_io_state_in_9),
    .io_state_in_10(ShiftRows_io_state_in_10),
    .io_state_in_11(ShiftRows_io_state_in_11),
    .io_state_in_12(ShiftRows_io_state_in_12),
    .io_state_in_13(ShiftRows_io_state_in_13),
    .io_state_in_14(ShiftRows_io_state_in_14),
    .io_state_in_15(ShiftRows_io_state_in_15),
    .io_state_out_0(ShiftRows_io_state_out_0),
    .io_state_out_1(ShiftRows_io_state_out_1),
    .io_state_out_2(ShiftRows_io_state_out_2),
    .io_state_out_3(ShiftRows_io_state_out_3),
    .io_state_out_4(ShiftRows_io_state_out_4),
    .io_state_out_5(ShiftRows_io_state_out_5),
    .io_state_out_6(ShiftRows_io_state_out_6),
    .io_state_out_7(ShiftRows_io_state_out_7),
    .io_state_out_8(ShiftRows_io_state_out_8),
    .io_state_out_9(ShiftRows_io_state_out_9),
    .io_state_out_10(ShiftRows_io_state_out_10),
    .io_state_out_11(ShiftRows_io_state_out_11),
    .io_state_out_12(ShiftRows_io_state_out_12),
    .io_state_out_13(ShiftRows_io_state_out_13),
    .io_state_out_14(ShiftRows_io_state_out_14),
    .io_state_out_15(ShiftRows_io_state_out_15)
  );
  assign io_state_out_0 = r__0; // @[CipherRound.scala 61:18]
  assign io_state_out_1 = r__1; // @[CipherRound.scala 61:18]
  assign io_state_out_2 = r__2; // @[CipherRound.scala 61:18]
  assign io_state_out_3 = r__3; // @[CipherRound.scala 61:18]
  assign io_state_out_4 = r__4; // @[CipherRound.scala 61:18]
  assign io_state_out_5 = r__5; // @[CipherRound.scala 61:18]
  assign io_state_out_6 = r__6; // @[CipherRound.scala 61:18]
  assign io_state_out_7 = r__7; // @[CipherRound.scala 61:18]
  assign io_state_out_8 = r__8; // @[CipherRound.scala 61:18]
  assign io_state_out_9 = r__9; // @[CipherRound.scala 61:18]
  assign io_state_out_10 = r__10; // @[CipherRound.scala 61:18]
  assign io_state_out_11 = r__11; // @[CipherRound.scala 61:18]
  assign io_state_out_12 = r__12; // @[CipherRound.scala 61:18]
  assign io_state_out_13 = r__13; // @[CipherRound.scala 61:18]
  assign io_state_out_14 = r__14; // @[CipherRound.scala 61:18]
  assign io_state_out_15 = r__15; // @[CipherRound.scala 61:18]
  assign io_output_valid = r_1; // @[CipherRound.scala 62:21]
  assign AddRoundKey_io_state_in_0 = ShiftRows_io_state_out_0; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_1 = ShiftRows_io_state_out_1; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_2 = ShiftRows_io_state_out_2; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_3 = ShiftRows_io_state_out_3; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_4 = ShiftRows_io_state_out_4; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_5 = ShiftRows_io_state_out_5; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_6 = ShiftRows_io_state_out_6; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_7 = ShiftRows_io_state_out_7; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_8 = ShiftRows_io_state_out_8; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_9 = ShiftRows_io_state_out_9; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_10 = ShiftRows_io_state_out_10; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_11 = ShiftRows_io_state_out_11; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_12 = ShiftRows_io_state_out_12; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_13 = ShiftRows_io_state_out_13; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_14 = ShiftRows_io_state_out_14; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_state_in_15 = ShiftRows_io_state_out_15; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_roundKey_0 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_1 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_2 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_3 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_4 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_5 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_6 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_7 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_8 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_9 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_10 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_11 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_12 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_13 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_14 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign AddRoundKey_io_roundKey_15 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign ShiftRows_io_state_in_0 = SubBytes_io_state_out_0; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_1 = SubBytes_io_state_out_1; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_2 = SubBytes_io_state_out_2; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_3 = SubBytes_io_state_out_3; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_4 = SubBytes_io_state_out_4; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_5 = SubBytes_io_state_out_5; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_6 = SubBytes_io_state_out_6; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_7 = SubBytes_io_state_out_7; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_8 = SubBytes_io_state_out_8; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_9 = SubBytes_io_state_out_9; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_10 = SubBytes_io_state_out_10; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_11 = SubBytes_io_state_out_11; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_12 = SubBytes_io_state_out_12; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_13 = SubBytes_io_state_out_13; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_14 = SubBytes_io_state_out_14; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_15 = SubBytes_io_state_out_15; // @[CipherRound.scala 56:33]
  always @(posedge clock) begin
    r__0 <= AddRoundKey_io_state_out_0; // @[Reg.scala 15:16 16:{19,23}]
    r__1 <= AddRoundKey_io_state_out_1; // @[Reg.scala 15:16 16:{19,23}]
    r__2 <= AddRoundKey_io_state_out_2; // @[Reg.scala 15:16 16:{19,23}]
    r__3 <= AddRoundKey_io_state_out_3; // @[Reg.scala 15:16 16:{19,23}]
    r__4 <= AddRoundKey_io_state_out_4; // @[Reg.scala 15:16 16:{19,23}]
    r__5 <= AddRoundKey_io_state_out_5; // @[Reg.scala 15:16 16:{19,23}]
    r__6 <= AddRoundKey_io_state_out_6; // @[Reg.scala 15:16 16:{19,23}]
    r__7 <= AddRoundKey_io_state_out_7; // @[Reg.scala 15:16 16:{19,23}]
    r__8 <= AddRoundKey_io_state_out_8; // @[Reg.scala 15:16 16:{19,23}]
    r__9 <= AddRoundKey_io_state_out_9; // @[Reg.scala 15:16 16:{19,23}]
    r__10 <= AddRoundKey_io_state_out_10; // @[Reg.scala 15:16 16:{19,23}]
    r__11 <= AddRoundKey_io_state_out_11; // @[Reg.scala 15:16 16:{19,23}]
    r__12 <= AddRoundKey_io_state_out_12; // @[Reg.scala 15:16 16:{19,23}]
    r__13 <= AddRoundKey_io_state_out_13; // @[Reg.scala 15:16 16:{19,23}]
    r__14 <= AddRoundKey_io_state_out_14; // @[Reg.scala 15:16 16:{19,23}]
    r__15 <= AddRoundKey_io_state_out_15; // @[Reg.scala 15:16 16:{19,23}]
    r_1 <= io_input_valid; // @[Reg.scala 15:16 16:{19,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r__0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r__1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r__2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r__3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r__4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r__5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r__6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r__7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r__8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r__9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r__10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r__11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r__12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r__13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r__14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r__15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AESEncrypt(
  input   clock,
  input   io_input_valid,
  input   io_input_text_0,
  input   io_input_text_1,
  input   io_input_text_2,
  input   io_input_text_3,
  input   io_input_text_4,
  input   io_input_text_5,
  input   io_input_text_6,
  input   io_input_text_7,
  input   io_input_text_8,
  input   io_input_text_9,
  input   io_input_text_10,
  input   io_input_text_11,
  input   io_input_text_12,
  input   io_input_text_13,
  input   io_input_text_14,
  input   io_input_text_15,
  output  io_output_text_0,
  output  io_output_text_1,
  output  io_output_text_2,
  output  io_output_text_3,
  output  io_output_text_4,
  output  io_output_text_5,
  output  io_output_text_6,
  output  io_output_text_7,
  output  io_output_text_8,
  output  io_output_text_9,
  output  io_output_text_10,
  output  io_output_text_11,
  output  io_output_text_12,
  output  io_output_text_13,
  output  io_output_text_14,
  output  io_output_text_15,
  output  io_output_intermediate,
  output  io_output_valid
);
  wire  CipherRoundARK_clock; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_0; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_1; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_2; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_3; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_4; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_5; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_6; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_7; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_8; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_9; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_10; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_11; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_12; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_13; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_14; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_state_in_15; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_0; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_1; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_3; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_4; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_5; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_6; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_7; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_8; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_9; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_10; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_11; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_12; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_13; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_14; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_15; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_output_valid; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_clock; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_input_valid; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_0; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_1; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_3; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_4; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_5; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_6; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_7; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_8; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_9; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_10; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_11; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_12; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_13; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_14; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_15; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_output_valid; // @[CipherRound.scala 95:84]
  InvCipherRound CipherRoundARK ( // @[CipherRound.scala 95:84]
    .clock(CipherRoundARK_clock),
    .io_input_valid(CipherRoundARK_io_input_valid),
    .io_state_in_0(CipherRoundARK_io_state_in_0),
    .io_state_in_1(CipherRoundARK_io_state_in_1),
    .io_state_in_2(CipherRoundARK_io_state_in_2),
    .io_state_in_3(CipherRoundARK_io_state_in_3),
    .io_state_in_4(CipherRoundARK_io_state_in_4),
    .io_state_in_5(CipherRoundARK_io_state_in_5),
    .io_state_in_6(CipherRoundARK_io_state_in_6),
    .io_state_in_7(CipherRoundARK_io_state_in_7),
    .io_state_in_8(CipherRoundARK_io_state_in_8),
    .io_state_in_9(CipherRoundARK_io_state_in_9),
    .io_state_in_10(CipherRoundARK_io_state_in_10),
    .io_state_in_11(CipherRoundARK_io_state_in_11),
    .io_state_in_12(CipherRoundARK_io_state_in_12),
    .io_state_in_13(CipherRoundARK_io_state_in_13),
    .io_state_in_14(CipherRoundARK_io_state_in_14),
    .io_state_in_15(CipherRoundARK_io_state_in_15),
    .io_roundKey_0(CipherRoundARK_io_roundKey_0),
    .io_roundKey_1(CipherRoundARK_io_roundKey_1),
    .io_roundKey_2(CipherRoundARK_io_roundKey_2),
    .io_roundKey_3(CipherRoundARK_io_roundKey_3),
    .io_roundKey_4(CipherRoundARK_io_roundKey_4),
    .io_roundKey_5(CipherRoundARK_io_roundKey_5),
    .io_roundKey_6(CipherRoundARK_io_roundKey_6),
    .io_roundKey_7(CipherRoundARK_io_roundKey_7),
    .io_roundKey_8(CipherRoundARK_io_roundKey_8),
    .io_roundKey_9(CipherRoundARK_io_roundKey_9),
    .io_roundKey_10(CipherRoundARK_io_roundKey_10),
    .io_roundKey_11(CipherRoundARK_io_roundKey_11),
    .io_roundKey_12(CipherRoundARK_io_roundKey_12),
    .io_roundKey_13(CipherRoundARK_io_roundKey_13),
    .io_roundKey_14(CipherRoundARK_io_roundKey_14),
    .io_roundKey_15(CipherRoundARK_io_roundKey_15),
    .io_output_valid(CipherRoundARK_io_output_valid)
  );
  CipherRound_1 CipherRound ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_clock),
    .io_input_valid(CipherRound_io_input_valid),
    .io_roundKey_0(CipherRound_io_roundKey_0),
    .io_roundKey_1(CipherRound_io_roundKey_1),
    .io_roundKey_2(CipherRound_io_roundKey_2),
    .io_roundKey_3(CipherRound_io_roundKey_3),
    .io_roundKey_4(CipherRound_io_roundKey_4),
    .io_roundKey_5(CipherRound_io_roundKey_5),
    .io_roundKey_6(CipherRound_io_roundKey_6),
    .io_roundKey_7(CipherRound_io_roundKey_7),
    .io_roundKey_8(CipherRound_io_roundKey_8),
    .io_roundKey_9(CipherRound_io_roundKey_9),
    .io_roundKey_10(CipherRound_io_roundKey_10),
    .io_roundKey_11(CipherRound_io_roundKey_11),
    .io_roundKey_12(CipherRound_io_roundKey_12),
    .io_roundKey_13(CipherRound_io_roundKey_13),
    .io_roundKey_14(CipherRound_io_roundKey_14),
    .io_roundKey_15(CipherRound_io_roundKey_15),
    .io_state_out_2(CipherRound_io_state_out_2),
    .io_output_valid(CipherRound_io_output_valid)
  );
  CipherRound_1 CipherRound_1 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_1_clock),
    .io_input_valid(CipherRound_1_io_input_valid),
    .io_roundKey_0(CipherRound_1_io_roundKey_0),
    .io_roundKey_1(CipherRound_1_io_roundKey_1),
    .io_roundKey_2(CipherRound_1_io_roundKey_2),
    .io_roundKey_3(CipherRound_1_io_roundKey_3),
    .io_roundKey_4(CipherRound_1_io_roundKey_4),
    .io_roundKey_5(CipherRound_1_io_roundKey_5),
    .io_roundKey_6(CipherRound_1_io_roundKey_6),
    .io_roundKey_7(CipherRound_1_io_roundKey_7),
    .io_roundKey_8(CipherRound_1_io_roundKey_8),
    .io_roundKey_9(CipherRound_1_io_roundKey_9),
    .io_roundKey_10(CipherRound_1_io_roundKey_10),
    .io_roundKey_11(CipherRound_1_io_roundKey_11),
    .io_roundKey_12(CipherRound_1_io_roundKey_12),
    .io_roundKey_13(CipherRound_1_io_roundKey_13),
    .io_roundKey_14(CipherRound_1_io_roundKey_14),
    .io_roundKey_15(CipherRound_1_io_roundKey_15),
    .io_state_out_2(CipherRound_1_io_state_out_2),
    .io_output_valid(CipherRound_1_io_output_valid)
  );
  CipherRound_1 CipherRound_2 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_2_clock),
    .io_input_valid(CipherRound_2_io_input_valid),
    .io_roundKey_0(CipherRound_2_io_roundKey_0),
    .io_roundKey_1(CipherRound_2_io_roundKey_1),
    .io_roundKey_2(CipherRound_2_io_roundKey_2),
    .io_roundKey_3(CipherRound_2_io_roundKey_3),
    .io_roundKey_4(CipherRound_2_io_roundKey_4),
    .io_roundKey_5(CipherRound_2_io_roundKey_5),
    .io_roundKey_6(CipherRound_2_io_roundKey_6),
    .io_roundKey_7(CipherRound_2_io_roundKey_7),
    .io_roundKey_8(CipherRound_2_io_roundKey_8),
    .io_roundKey_9(CipherRound_2_io_roundKey_9),
    .io_roundKey_10(CipherRound_2_io_roundKey_10),
    .io_roundKey_11(CipherRound_2_io_roundKey_11),
    .io_roundKey_12(CipherRound_2_io_roundKey_12),
    .io_roundKey_13(CipherRound_2_io_roundKey_13),
    .io_roundKey_14(CipherRound_2_io_roundKey_14),
    .io_roundKey_15(CipherRound_2_io_roundKey_15),
    .io_state_out_2(CipherRound_2_io_state_out_2),
    .io_output_valid(CipherRound_2_io_output_valid)
  );
  CipherRound_1 CipherRound_3 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_3_clock),
    .io_input_valid(CipherRound_3_io_input_valid),
    .io_roundKey_0(CipherRound_3_io_roundKey_0),
    .io_roundKey_1(CipherRound_3_io_roundKey_1),
    .io_roundKey_2(CipherRound_3_io_roundKey_2),
    .io_roundKey_3(CipherRound_3_io_roundKey_3),
    .io_roundKey_4(CipherRound_3_io_roundKey_4),
    .io_roundKey_5(CipherRound_3_io_roundKey_5),
    .io_roundKey_6(CipherRound_3_io_roundKey_6),
    .io_roundKey_7(CipherRound_3_io_roundKey_7),
    .io_roundKey_8(CipherRound_3_io_roundKey_8),
    .io_roundKey_9(CipherRound_3_io_roundKey_9),
    .io_roundKey_10(CipherRound_3_io_roundKey_10),
    .io_roundKey_11(CipherRound_3_io_roundKey_11),
    .io_roundKey_12(CipherRound_3_io_roundKey_12),
    .io_roundKey_13(CipherRound_3_io_roundKey_13),
    .io_roundKey_14(CipherRound_3_io_roundKey_14),
    .io_roundKey_15(CipherRound_3_io_roundKey_15),
    .io_state_out_2(CipherRound_3_io_state_out_2),
    .io_output_valid(CipherRound_3_io_output_valid)
  );
  CipherRound_1 CipherRound_4 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_4_clock),
    .io_input_valid(CipherRound_4_io_input_valid),
    .io_roundKey_0(CipherRound_4_io_roundKey_0),
    .io_roundKey_1(CipherRound_4_io_roundKey_1),
    .io_roundKey_2(CipherRound_4_io_roundKey_2),
    .io_roundKey_3(CipherRound_4_io_roundKey_3),
    .io_roundKey_4(CipherRound_4_io_roundKey_4),
    .io_roundKey_5(CipherRound_4_io_roundKey_5),
    .io_roundKey_6(CipherRound_4_io_roundKey_6),
    .io_roundKey_7(CipherRound_4_io_roundKey_7),
    .io_roundKey_8(CipherRound_4_io_roundKey_8),
    .io_roundKey_9(CipherRound_4_io_roundKey_9),
    .io_roundKey_10(CipherRound_4_io_roundKey_10),
    .io_roundKey_11(CipherRound_4_io_roundKey_11),
    .io_roundKey_12(CipherRound_4_io_roundKey_12),
    .io_roundKey_13(CipherRound_4_io_roundKey_13),
    .io_roundKey_14(CipherRound_4_io_roundKey_14),
    .io_roundKey_15(CipherRound_4_io_roundKey_15),
    .io_state_out_2(CipherRound_4_io_state_out_2),
    .io_output_valid(CipherRound_4_io_output_valid)
  );
  CipherRound_1 CipherRound_5 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_5_clock),
    .io_input_valid(CipherRound_5_io_input_valid),
    .io_roundKey_0(CipherRound_5_io_roundKey_0),
    .io_roundKey_1(CipherRound_5_io_roundKey_1),
    .io_roundKey_2(CipherRound_5_io_roundKey_2),
    .io_roundKey_3(CipherRound_5_io_roundKey_3),
    .io_roundKey_4(CipherRound_5_io_roundKey_4),
    .io_roundKey_5(CipherRound_5_io_roundKey_5),
    .io_roundKey_6(CipherRound_5_io_roundKey_6),
    .io_roundKey_7(CipherRound_5_io_roundKey_7),
    .io_roundKey_8(CipherRound_5_io_roundKey_8),
    .io_roundKey_9(CipherRound_5_io_roundKey_9),
    .io_roundKey_10(CipherRound_5_io_roundKey_10),
    .io_roundKey_11(CipherRound_5_io_roundKey_11),
    .io_roundKey_12(CipherRound_5_io_roundKey_12),
    .io_roundKey_13(CipherRound_5_io_roundKey_13),
    .io_roundKey_14(CipherRound_5_io_roundKey_14),
    .io_roundKey_15(CipherRound_5_io_roundKey_15),
    .io_state_out_2(CipherRound_5_io_state_out_2),
    .io_output_valid(CipherRound_5_io_output_valid)
  );
  CipherRound_1 CipherRound_6 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_6_clock),
    .io_input_valid(CipherRound_6_io_input_valid),
    .io_roundKey_0(CipherRound_6_io_roundKey_0),
    .io_roundKey_1(CipherRound_6_io_roundKey_1),
    .io_roundKey_2(CipherRound_6_io_roundKey_2),
    .io_roundKey_3(CipherRound_6_io_roundKey_3),
    .io_roundKey_4(CipherRound_6_io_roundKey_4),
    .io_roundKey_5(CipherRound_6_io_roundKey_5),
    .io_roundKey_6(CipherRound_6_io_roundKey_6),
    .io_roundKey_7(CipherRound_6_io_roundKey_7),
    .io_roundKey_8(CipherRound_6_io_roundKey_8),
    .io_roundKey_9(CipherRound_6_io_roundKey_9),
    .io_roundKey_10(CipherRound_6_io_roundKey_10),
    .io_roundKey_11(CipherRound_6_io_roundKey_11),
    .io_roundKey_12(CipherRound_6_io_roundKey_12),
    .io_roundKey_13(CipherRound_6_io_roundKey_13),
    .io_roundKey_14(CipherRound_6_io_roundKey_14),
    .io_roundKey_15(CipherRound_6_io_roundKey_15),
    .io_state_out_2(CipherRound_6_io_state_out_2),
    .io_output_valid(CipherRound_6_io_output_valid)
  );
  CipherRound_1 CipherRound_7 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_7_clock),
    .io_input_valid(CipherRound_7_io_input_valid),
    .io_roundKey_0(CipherRound_7_io_roundKey_0),
    .io_roundKey_1(CipherRound_7_io_roundKey_1),
    .io_roundKey_2(CipherRound_7_io_roundKey_2),
    .io_roundKey_3(CipherRound_7_io_roundKey_3),
    .io_roundKey_4(CipherRound_7_io_roundKey_4),
    .io_roundKey_5(CipherRound_7_io_roundKey_5),
    .io_roundKey_6(CipherRound_7_io_roundKey_6),
    .io_roundKey_7(CipherRound_7_io_roundKey_7),
    .io_roundKey_8(CipherRound_7_io_roundKey_8),
    .io_roundKey_9(CipherRound_7_io_roundKey_9),
    .io_roundKey_10(CipherRound_7_io_roundKey_10),
    .io_roundKey_11(CipherRound_7_io_roundKey_11),
    .io_roundKey_12(CipherRound_7_io_roundKey_12),
    .io_roundKey_13(CipherRound_7_io_roundKey_13),
    .io_roundKey_14(CipherRound_7_io_roundKey_14),
    .io_roundKey_15(CipherRound_7_io_roundKey_15),
    .io_state_out_2(CipherRound_7_io_state_out_2),
    .io_output_valid(CipherRound_7_io_output_valid)
  );
  CipherRound_1 CipherRound_8 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_8_clock),
    .io_input_valid(CipherRound_8_io_input_valid),
    .io_roundKey_0(CipherRound_8_io_roundKey_0),
    .io_roundKey_1(CipherRound_8_io_roundKey_1),
    .io_roundKey_2(CipherRound_8_io_roundKey_2),
    .io_roundKey_3(CipherRound_8_io_roundKey_3),
    .io_roundKey_4(CipherRound_8_io_roundKey_4),
    .io_roundKey_5(CipherRound_8_io_roundKey_5),
    .io_roundKey_6(CipherRound_8_io_roundKey_6),
    .io_roundKey_7(CipherRound_8_io_roundKey_7),
    .io_roundKey_8(CipherRound_8_io_roundKey_8),
    .io_roundKey_9(CipherRound_8_io_roundKey_9),
    .io_roundKey_10(CipherRound_8_io_roundKey_10),
    .io_roundKey_11(CipherRound_8_io_roundKey_11),
    .io_roundKey_12(CipherRound_8_io_roundKey_12),
    .io_roundKey_13(CipherRound_8_io_roundKey_13),
    .io_roundKey_14(CipherRound_8_io_roundKey_14),
    .io_roundKey_15(CipherRound_8_io_roundKey_15),
    .io_state_out_2(CipherRound_8_io_state_out_2),
    .io_output_valid(CipherRound_8_io_output_valid)
  );
  CipherRound_10 CipherRoundNMC ( // @[CipherRound.scala 95:84]
    .clock(CipherRoundNMC_clock),
    .io_input_valid(CipherRoundNMC_io_input_valid),
    .io_state_out_0(CipherRoundNMC_io_state_out_0),
    .io_state_out_1(CipherRoundNMC_io_state_out_1),
    .io_state_out_2(CipherRoundNMC_io_state_out_2),
    .io_state_out_3(CipherRoundNMC_io_state_out_3),
    .io_state_out_4(CipherRoundNMC_io_state_out_4),
    .io_state_out_5(CipherRoundNMC_io_state_out_5),
    .io_state_out_6(CipherRoundNMC_io_state_out_6),
    .io_state_out_7(CipherRoundNMC_io_state_out_7),
    .io_state_out_8(CipherRoundNMC_io_state_out_8),
    .io_state_out_9(CipherRoundNMC_io_state_out_9),
    .io_state_out_10(CipherRoundNMC_io_state_out_10),
    .io_state_out_11(CipherRoundNMC_io_state_out_11),
    .io_state_out_12(CipherRoundNMC_io_state_out_12),
    .io_state_out_13(CipherRoundNMC_io_state_out_13),
    .io_state_out_14(CipherRoundNMC_io_state_out_14),
    .io_state_out_15(CipherRoundNMC_io_state_out_15),
    .io_output_valid(CipherRoundNMC_io_output_valid)
  );
  assign io_output_text_0 = CipherRoundNMC_io_state_out_0; // @[AESEncrypt.scala 54:18]
  assign io_output_text_1 = CipherRoundNMC_io_state_out_1; // @[AESEncrypt.scala 54:18]
  assign io_output_text_2 = CipherRoundNMC_io_state_out_2; // @[AESEncrypt.scala 54:18]
  assign io_output_text_3 = CipherRoundNMC_io_state_out_3; // @[AESEncrypt.scala 54:18]
  assign io_output_text_4 = CipherRoundNMC_io_state_out_4; // @[AESEncrypt.scala 54:18]
  assign io_output_text_5 = CipherRoundNMC_io_state_out_5; // @[AESEncrypt.scala 54:18]
  assign io_output_text_6 = CipherRoundNMC_io_state_out_6; // @[AESEncrypt.scala 54:18]
  assign io_output_text_7 = CipherRoundNMC_io_state_out_7; // @[AESEncrypt.scala 54:18]
  assign io_output_text_8 = CipherRoundNMC_io_state_out_8; // @[AESEncrypt.scala 54:18]
  assign io_output_text_9 = CipherRoundNMC_io_state_out_9; // @[AESEncrypt.scala 54:18]
  assign io_output_text_10 = CipherRoundNMC_io_state_out_10; // @[AESEncrypt.scala 54:18]
  assign io_output_text_11 = CipherRoundNMC_io_state_out_11; // @[AESEncrypt.scala 54:18]
  assign io_output_text_12 = CipherRoundNMC_io_state_out_12; // @[AESEncrypt.scala 54:18]
  assign io_output_text_13 = CipherRoundNMC_io_state_out_13; // @[AESEncrypt.scala 54:18]
  assign io_output_text_14 = CipherRoundNMC_io_state_out_14; // @[AESEncrypt.scala 54:18]
  assign io_output_text_15 = CipherRoundNMC_io_state_out_15; // @[AESEncrypt.scala 54:18]
  assign io_output_intermediate = CipherRound_3_io_state_out_2; // @[AESEncrypt.scala 52:26]
  assign io_output_valid = CipherRoundNMC_io_output_valid; // @[AESEncrypt.scala 53:19]
  assign CipherRoundARK_clock = clock;
  assign CipherRoundARK_io_input_valid = io_input_valid; // @[AESEncrypt.scala 31:33]
  assign CipherRoundARK_io_state_in_0 = io_input_text_0; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_1 = io_input_text_1; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_2 = io_input_text_2; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_3 = io_input_text_3; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_4 = io_input_text_4; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_5 = io_input_text_5; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_6 = io_input_text_6; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_7 = io_input_text_7; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_8 = io_input_text_8; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_9 = io_input_text_9; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_10 = io_input_text_10; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_11 = io_input_text_11; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_12 = io_input_text_12; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_13 = io_input_text_13; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_14 = io_input_text_14; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_state_in_15 = io_input_text_15; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRoundARK_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRound_clock = clock;
  assign CipherRound_io_input_valid = CipherRoundARK_io_output_valid; // @[AESEncrypt.scala 38:38]
  assign CipherRound_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_clock = clock;
  assign CipherRound_1_io_input_valid = CipherRound_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_1_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_clock = clock;
  assign CipherRound_2_io_input_valid = CipherRound_1_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_2_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_clock = clock;
  assign CipherRound_3_io_input_valid = CipherRound_2_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_3_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_clock = clock;
  assign CipherRound_4_io_input_valid = CipherRound_3_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_4_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_clock = clock;
  assign CipherRound_5_io_input_valid = CipherRound_4_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_5_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_clock = clock;
  assign CipherRound_6_io_input_valid = CipherRound_5_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_6_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_clock = clock;
  assign CipherRound_7_io_input_valid = CipherRound_6_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_7_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_clock = clock;
  assign CipherRound_8_io_input_valid = CipherRound_7_io_output_valid; // @[AESEncrypt.scala 42:38]
  assign CipherRound_8_io_roundKey_0 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_1 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_3 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_4 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_5 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_6 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_7 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_8 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_9 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_10 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_11 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_12 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_13 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_14 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_io_roundKey_15 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRoundNMC_clock = clock;
  assign CipherRoundNMC_io_input_valid = CipherRound_8_io_output_valid; // @[AESEncrypt.scala 49:33]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19,
  output  io_out_20,
  output  io_out_21,
  output  io_out_22,
  output  io_out_23,
  output  io_out_24,
  output  io_out_25,
  output  io_out_26,
  output  io_out_27,
  output  io_out_28,
  output  io_out_29,
  output  io_out_30,
  output  io_out_31,
  output  io_out_32,
  output  io_out_33,
  output  io_out_34,
  output  io_out_35,
  output  io_out_36,
  output  io_out_37,
  output  io_out_38,
  output  io_out_39,
  output  io_out_40,
  output  io_out_41,
  output  io_out_42,
  output  io_out_43,
  output  io_out_44,
  output  io_out_45,
  output  io_out_46,
  output  io_out_47,
  output  io_out_48,
  output  io_out_49,
  output  io_out_50,
  output  io_out_51,
  output  io_out_52,
  output  io_out_53,
  output  io_out_54,
  output  io_out_55,
  output  io_out_56,
  output  io_out_57,
  output  io_out_58,
  output  io_out_59,
  output  io_out_60,
  output  io_out_61,
  output  io_out_62,
  output  io_out_63
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 47:50]
  reg  state_1; // @[PRNG.scala 47:50]
  reg  state_2; // @[PRNG.scala 47:50]
  reg  state_3; // @[PRNG.scala 47:50]
  reg  state_4; // @[PRNG.scala 47:50]
  reg  state_5; // @[PRNG.scala 47:50]
  reg  state_6; // @[PRNG.scala 47:50]
  reg  state_7; // @[PRNG.scala 47:50]
  reg  state_8; // @[PRNG.scala 47:50]
  reg  state_9; // @[PRNG.scala 47:50]
  reg  state_10; // @[PRNG.scala 47:50]
  reg  state_11; // @[PRNG.scala 47:50]
  reg  state_12; // @[PRNG.scala 47:50]
  reg  state_13; // @[PRNG.scala 47:50]
  reg  state_14; // @[PRNG.scala 47:50]
  reg  state_15; // @[PRNG.scala 47:50]
  reg  state_16; // @[PRNG.scala 47:50]
  reg  state_17; // @[PRNG.scala 47:50]
  reg  state_18; // @[PRNG.scala 47:50]
  reg  state_19; // @[PRNG.scala 47:50]
  reg  state_20; // @[PRNG.scala 47:50]
  reg  state_21; // @[PRNG.scala 47:50]
  reg  state_22; // @[PRNG.scala 47:50]
  reg  state_23; // @[PRNG.scala 47:50]
  reg  state_24; // @[PRNG.scala 47:50]
  reg  state_25; // @[PRNG.scala 47:50]
  reg  state_26; // @[PRNG.scala 47:50]
  reg  state_27; // @[PRNG.scala 47:50]
  reg  state_28; // @[PRNG.scala 47:50]
  reg  state_29; // @[PRNG.scala 47:50]
  reg  state_30; // @[PRNG.scala 47:50]
  reg  state_31; // @[PRNG.scala 47:50]
  reg  state_32; // @[PRNG.scala 47:50]
  reg  state_33; // @[PRNG.scala 47:50]
  reg  state_34; // @[PRNG.scala 47:50]
  reg  state_35; // @[PRNG.scala 47:50]
  reg  state_36; // @[PRNG.scala 47:50]
  reg  state_37; // @[PRNG.scala 47:50]
  reg  state_38; // @[PRNG.scala 47:50]
  reg  state_39; // @[PRNG.scala 47:50]
  reg  state_40; // @[PRNG.scala 47:50]
  reg  state_41; // @[PRNG.scala 47:50]
  reg  state_42; // @[PRNG.scala 47:50]
  reg  state_43; // @[PRNG.scala 47:50]
  reg  state_44; // @[PRNG.scala 47:50]
  reg  state_45; // @[PRNG.scala 47:50]
  reg  state_46; // @[PRNG.scala 47:50]
  reg  state_47; // @[PRNG.scala 47:50]
  reg  state_48; // @[PRNG.scala 47:50]
  reg  state_49; // @[PRNG.scala 47:50]
  reg  state_50; // @[PRNG.scala 47:50]
  reg  state_51; // @[PRNG.scala 47:50]
  reg  state_52; // @[PRNG.scala 47:50]
  reg  state_53; // @[PRNG.scala 47:50]
  reg  state_54; // @[PRNG.scala 47:50]
  reg  state_55; // @[PRNG.scala 47:50]
  reg  state_56; // @[PRNG.scala 47:50]
  reg  state_57; // @[PRNG.scala 47:50]
  reg  state_58; // @[PRNG.scala 47:50]
  reg  state_59; // @[PRNG.scala 47:50]
  reg  state_60; // @[PRNG.scala 47:50]
  reg  state_61; // @[PRNG.scala 47:50]
  reg  state_62; // @[PRNG.scala 47:50]
  reg  state_63; // @[PRNG.scala 47:50]
  wire  _T_2 = state_63 & state_62 & state_60 & state_59; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  assign io_out_4 = state_4; // @[PRNG.scala 69:10]
  assign io_out_5 = state_5; // @[PRNG.scala 69:10]
  assign io_out_6 = state_6; // @[PRNG.scala 69:10]
  assign io_out_7 = state_7; // @[PRNG.scala 69:10]
  assign io_out_8 = state_8; // @[PRNG.scala 69:10]
  assign io_out_9 = state_9; // @[PRNG.scala 69:10]
  assign io_out_10 = state_10; // @[PRNG.scala 69:10]
  assign io_out_11 = state_11; // @[PRNG.scala 69:10]
  assign io_out_12 = state_12; // @[PRNG.scala 69:10]
  assign io_out_13 = state_13; // @[PRNG.scala 69:10]
  assign io_out_14 = state_14; // @[PRNG.scala 69:10]
  assign io_out_15 = state_15; // @[PRNG.scala 69:10]
  assign io_out_16 = state_16; // @[PRNG.scala 69:10]
  assign io_out_17 = state_17; // @[PRNG.scala 69:10]
  assign io_out_18 = state_18; // @[PRNG.scala 69:10]
  assign io_out_19 = state_19; // @[PRNG.scala 69:10]
  assign io_out_20 = state_20; // @[PRNG.scala 69:10]
  assign io_out_21 = state_21; // @[PRNG.scala 69:10]
  assign io_out_22 = state_22; // @[PRNG.scala 69:10]
  assign io_out_23 = state_23; // @[PRNG.scala 69:10]
  assign io_out_24 = state_24; // @[PRNG.scala 69:10]
  assign io_out_25 = state_25; // @[PRNG.scala 69:10]
  assign io_out_26 = state_26; // @[PRNG.scala 69:10]
  assign io_out_27 = state_27; // @[PRNG.scala 69:10]
  assign io_out_28 = state_28; // @[PRNG.scala 69:10]
  assign io_out_29 = state_29; // @[PRNG.scala 69:10]
  assign io_out_30 = state_30; // @[PRNG.scala 69:10]
  assign io_out_31 = state_31; // @[PRNG.scala 69:10]
  assign io_out_32 = state_32; // @[PRNG.scala 69:10]
  assign io_out_33 = state_33; // @[PRNG.scala 69:10]
  assign io_out_34 = state_34; // @[PRNG.scala 69:10]
  assign io_out_35 = state_35; // @[PRNG.scala 69:10]
  assign io_out_36 = state_36; // @[PRNG.scala 69:10]
  assign io_out_37 = state_37; // @[PRNG.scala 69:10]
  assign io_out_38 = state_38; // @[PRNG.scala 69:10]
  assign io_out_39 = state_39; // @[PRNG.scala 69:10]
  assign io_out_40 = state_40; // @[PRNG.scala 69:10]
  assign io_out_41 = state_41; // @[PRNG.scala 69:10]
  assign io_out_42 = state_42; // @[PRNG.scala 69:10]
  assign io_out_43 = state_43; // @[PRNG.scala 69:10]
  assign io_out_44 = state_44; // @[PRNG.scala 69:10]
  assign io_out_45 = state_45; // @[PRNG.scala 69:10]
  assign io_out_46 = state_46; // @[PRNG.scala 69:10]
  assign io_out_47 = state_47; // @[PRNG.scala 69:10]
  assign io_out_48 = state_48; // @[PRNG.scala 69:10]
  assign io_out_49 = state_49; // @[PRNG.scala 69:10]
  assign io_out_50 = state_50; // @[PRNG.scala 69:10]
  assign io_out_51 = state_51; // @[PRNG.scala 69:10]
  assign io_out_52 = state_52; // @[PRNG.scala 69:10]
  assign io_out_53 = state_53; // @[PRNG.scala 69:10]
  assign io_out_54 = state_54; // @[PRNG.scala 69:10]
  assign io_out_55 = state_55; // @[PRNG.scala 69:10]
  assign io_out_56 = state_56; // @[PRNG.scala 69:10]
  assign io_out_57 = state_57; // @[PRNG.scala 69:10]
  assign io_out_58 = state_58; // @[PRNG.scala 69:10]
  assign io_out_59 = state_59; // @[PRNG.scala 69:10]
  assign io_out_60 = state_60; // @[PRNG.scala 69:10]
  assign io_out_61 = state_61; // @[PRNG.scala 69:10]
  assign io_out_62 = state_62; // @[PRNG.scala 69:10]
  assign io_out_63 = state_63; // @[PRNG.scala 69:10]
  always @(posedge clock) begin
    state_0 <= 1'h1 & _T_2; // @[PRNG.scala 47:{50,50}]
    state_1 <= reset & state_0; // @[PRNG.scala 47:{50,50}]
    state_2 <= reset & state_1; // @[PRNG.scala 47:{50,50}]
    state_3 <= 1'h1 & state_2; // @[PRNG.scala 47:{50,50}]
    state_4 <= 1'h1 & state_3; // @[PRNG.scala 47:{50,50}]
    state_5 <= 1'h1 & state_4; // @[PRNG.scala 47:{50,50}]
    state_6 <= 1'h1 & state_5; // @[PRNG.scala 47:{50,50}]
    state_7 <= reset & state_6; // @[PRNG.scala 47:{50,50}]
    state_8 <= reset & state_7; // @[PRNG.scala 47:{50,50}]
    state_9 <= reset & state_8; // @[PRNG.scala 47:{50,50}]
    state_10 <= reset & state_9; // @[PRNG.scala 47:{50,50}]
    state_11 <= reset & state_10; // @[PRNG.scala 47:{50,50}]
    state_12 <= reset & state_11; // @[PRNG.scala 47:{50,50}]
    state_13 <= reset & state_12; // @[PRNG.scala 47:{50,50}]
    state_14 <= reset & state_13; // @[PRNG.scala 47:{50,50}]
    state_15 <= 1'h1 & state_14; // @[PRNG.scala 47:{50,50}]
    state_16 <= reset & state_15; // @[PRNG.scala 47:{50,50}]
    state_17 <= 1'h1 & state_16; // @[PRNG.scala 47:{50,50}]
    state_18 <= reset & state_17; // @[PRNG.scala 47:{50,50}]
    state_19 <= 1'h1 & state_18; // @[PRNG.scala 47:{50,50}]
    state_20 <= reset & state_19; // @[PRNG.scala 47:{50,50}]
    state_21 <= reset & state_20; // @[PRNG.scala 47:{50,50}]
    state_22 <= reset & state_21; // @[PRNG.scala 47:{50,50}]
    state_23 <= reset & state_22; // @[PRNG.scala 47:{50,50}]
    state_24 <= 1'h1 & state_23; // @[PRNG.scala 47:{50,50}]
    state_25 <= 1'h1 & state_24; // @[PRNG.scala 47:{50,50}]
    state_26 <= reset & state_25; // @[PRNG.scala 47:{50,50}]
    state_27 <= 1'h1 & state_26; // @[PRNG.scala 47:{50,50}]
    state_28 <= reset & state_27; // @[PRNG.scala 47:{50,50}]
    state_29 <= 1'h1 & state_28; // @[PRNG.scala 47:{50,50}]
    state_30 <= 1'h1 & state_29; // @[PRNG.scala 47:{50,50}]
    state_31 <= 1'h1 & state_30; // @[PRNG.scala 47:{50,50}]
    state_32 <= 1'h1 & state_31; // @[PRNG.scala 47:{50,50}]
    state_33 <= reset & state_32; // @[PRNG.scala 47:{50,50}]
    state_34 <= reset & state_33; // @[PRNG.scala 47:{50,50}]
    state_35 <= reset & state_34; // @[PRNG.scala 47:{50,50}]
    state_36 <= reset & state_35; // @[PRNG.scala 47:{50,50}]
    state_37 <= 1'h1 & state_36; // @[PRNG.scala 47:{50,50}]
    state_38 <= 1'h1 & state_37; // @[PRNG.scala 47:{50,50}]
    state_39 <= 1'h1 & state_38; // @[PRNG.scala 47:{50,50}]
    state_40 <= reset & state_39; // @[PRNG.scala 47:{50,50}]
    state_41 <= reset & state_40; // @[PRNG.scala 47:{50,50}]
    state_42 <= reset & state_41; // @[PRNG.scala 47:{50,50}]
    state_43 <= reset & state_42; // @[PRNG.scala 47:{50,50}]
    state_44 <= 1'h1 & state_43; // @[PRNG.scala 47:{50,50}]
    state_45 <= reset & state_44; // @[PRNG.scala 47:{50,50}]
    state_46 <= 1'h1 & state_45; // @[PRNG.scala 47:{50,50}]
    state_47 <= 1'h1 & state_46; // @[PRNG.scala 47:{50,50}]
    state_48 <= reset & state_47; // @[PRNG.scala 47:{50,50}]
    state_49 <= 1'h1 & state_48; // @[PRNG.scala 47:{50,50}]
    state_50 <= 1'h1 & state_49; // @[PRNG.scala 47:{50,50}]
    state_51 <= reset & state_50; // @[PRNG.scala 47:{50,50}]
    state_52 <= 1'h1 & state_51; // @[PRNG.scala 47:{50,50}]
    state_53 <= 1'h1 & state_52; // @[PRNG.scala 47:{50,50}]
    state_54 <= reset & state_53; // @[PRNG.scala 47:{50,50}]
    state_55 <= reset & state_54; // @[PRNG.scala 47:{50,50}]
    state_56 <= reset & state_55; // @[PRNG.scala 47:{50,50}]
    state_57 <= 1'h1 & state_56; // @[PRNG.scala 47:{50,50}]
    state_58 <= reset & state_57; // @[PRNG.scala 47:{50,50}]
    state_59 <= reset & state_58; // @[PRNG.scala 47:{50,50}]
    state_60 <= reset & state_59; // @[PRNG.scala 47:{50,50}]
    state_61 <= 1'h1 & state_60; // @[PRNG.scala 47:{50,50}]
    state_62 <= 1'h1 & state_61; // @[PRNG.scala 47:{50,50}]
    state_63 <= reset & state_62; // @[PRNG.scala 47:{50,50}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  state_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  state_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  state_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  state_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  state_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  state_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  state_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  state_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  state_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  state_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  state_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  state_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  state_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  state_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  state_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  state_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  state_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  state_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  state_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  state_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  state_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  state_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  state_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  state_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  state_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  state_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  state_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  state_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  state_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  state_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  state_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  state_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  state_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  state_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  state_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  state_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  state_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  state_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  state_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  state_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  state_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  state_63 = _RAND_63[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SE(
  input   clock,
  input   reset,
  input   io_in_inst,
  input   io_in_op1,
  input   io_in_op2,
  input   io_in_cond,
  input   io_in_valid,
  output  io_in_ready,
  output  io_out_result,
  output  io_out_valid,
  input   io_out_ready,
  output  io_out_cntr,
  output  io_out_zero_cntr,
  output  io_out_mult_cntr,
  output  io_out_intermediate
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  seoperation_io_op1_input; // @[SE.scala 83:33]
  wire  seoperation_io_op2_input; // @[SE.scala 83:33]
  wire  seoperation_io_result; // @[SE.scala 83:33]
  wire  aes_invcipher_clock; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_valid; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op1_15; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_15; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_15; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_15; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_15; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_valid; // @[SE.scala 84:35]
  wire  aes_cipher_clock; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_valid; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_0; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_1; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_2; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_3; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_4; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_5; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_6; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_7; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_8; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_9; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_10; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_11; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_12; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_13; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_14; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_15; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_0; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_1; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_2; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_3; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_4; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_5; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_6; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_7; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_8; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_9; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_10; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_11; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_12; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_13; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_14; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_15; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_intermediate; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_valid; // @[SE.scala 85:32]
  wire  prng_clock; // @[PRNG.scala 82:22]
  wire  prng_reset; // @[PRNG.scala 82:22]
  wire  prng_io_out_0; // @[PRNG.scala 82:22]
  wire  prng_io_out_1; // @[PRNG.scala 82:22]
  wire  prng_io_out_2; // @[PRNG.scala 82:22]
  wire  prng_io_out_3; // @[PRNG.scala 82:22]
  wire  prng_io_out_4; // @[PRNG.scala 82:22]
  wire  prng_io_out_5; // @[PRNG.scala 82:22]
  wire  prng_io_out_6; // @[PRNG.scala 82:22]
  wire  prng_io_out_7; // @[PRNG.scala 82:22]
  wire  prng_io_out_8; // @[PRNG.scala 82:22]
  wire  prng_io_out_9; // @[PRNG.scala 82:22]
  wire  prng_io_out_10; // @[PRNG.scala 82:22]
  wire  prng_io_out_11; // @[PRNG.scala 82:22]
  wire  prng_io_out_12; // @[PRNG.scala 82:22]
  wire  prng_io_out_13; // @[PRNG.scala 82:22]
  wire  prng_io_out_14; // @[PRNG.scala 82:22]
  wire  prng_io_out_15; // @[PRNG.scala 82:22]
  wire  prng_io_out_16; // @[PRNG.scala 82:22]
  wire  prng_io_out_17; // @[PRNG.scala 82:22]
  wire  prng_io_out_18; // @[PRNG.scala 82:22]
  wire  prng_io_out_19; // @[PRNG.scala 82:22]
  wire  prng_io_out_20; // @[PRNG.scala 82:22]
  wire  prng_io_out_21; // @[PRNG.scala 82:22]
  wire  prng_io_out_22; // @[PRNG.scala 82:22]
  wire  prng_io_out_23; // @[PRNG.scala 82:22]
  wire  prng_io_out_24; // @[PRNG.scala 82:22]
  wire  prng_io_out_25; // @[PRNG.scala 82:22]
  wire  prng_io_out_26; // @[PRNG.scala 82:22]
  wire  prng_io_out_27; // @[PRNG.scala 82:22]
  wire  prng_io_out_28; // @[PRNG.scala 82:22]
  wire  prng_io_out_29; // @[PRNG.scala 82:22]
  wire  prng_io_out_30; // @[PRNG.scala 82:22]
  wire  prng_io_out_31; // @[PRNG.scala 82:22]
  wire  prng_io_out_32; // @[PRNG.scala 82:22]
  wire  prng_io_out_33; // @[PRNG.scala 82:22]
  wire  prng_io_out_34; // @[PRNG.scala 82:22]
  wire  prng_io_out_35; // @[PRNG.scala 82:22]
  wire  prng_io_out_36; // @[PRNG.scala 82:22]
  wire  prng_io_out_37; // @[PRNG.scala 82:22]
  wire  prng_io_out_38; // @[PRNG.scala 82:22]
  wire  prng_io_out_39; // @[PRNG.scala 82:22]
  wire  prng_io_out_40; // @[PRNG.scala 82:22]
  wire  prng_io_out_41; // @[PRNG.scala 82:22]
  wire  prng_io_out_42; // @[PRNG.scala 82:22]
  wire  prng_io_out_43; // @[PRNG.scala 82:22]
  wire  prng_io_out_44; // @[PRNG.scala 82:22]
  wire  prng_io_out_45; // @[PRNG.scala 82:22]
  wire  prng_io_out_46; // @[PRNG.scala 82:22]
  wire  prng_io_out_47; // @[PRNG.scala 82:22]
  wire  prng_io_out_48; // @[PRNG.scala 82:22]
  wire  prng_io_out_49; // @[PRNG.scala 82:22]
  wire  prng_io_out_50; // @[PRNG.scala 82:22]
  wire  prng_io_out_51; // @[PRNG.scala 82:22]
  wire  prng_io_out_52; // @[PRNG.scala 82:22]
  wire  prng_io_out_53; // @[PRNG.scala 82:22]
  wire  prng_io_out_54; // @[PRNG.scala 82:22]
  wire  prng_io_out_55; // @[PRNG.scala 82:22]
  wire  prng_io_out_56; // @[PRNG.scala 82:22]
  wire  prng_io_out_57; // @[PRNG.scala 82:22]
  wire  prng_io_out_58; // @[PRNG.scala 82:22]
  wire  prng_io_out_59; // @[PRNG.scala 82:22]
  wire  prng_io_out_60; // @[PRNG.scala 82:22]
  wire  prng_io_out_61; // @[PRNG.scala 82:22]
  wire  prng_io_out_62; // @[PRNG.scala 82:22]
  wire  prng_io_out_63; // @[PRNG.scala 82:22]
  reg  value; // @[Counter.scala 60:40]
  reg  zero_cntr; // @[SE.scala 63:32]
  reg  mult_cntr; // @[SE.scala 64:32]
  wire  _GEN_0 = 1'h1 & (value & 1'h1); // @[Counter.scala 76:15 86:{20,28}]
  wire  _GEN_1 = _GEN_0 & value; // @[SE.scala 67:24 Counter.scala 60:40]
  wire  _T = io_in_valid & io_in_ready; // @[SE.scala 70:26]
  wire  _T_1 = io_out_valid & io_out_ready; // @[SE.scala 72:33]
  wire  _GEN_4 = 1'h1 & _GEN_1; // @[SE.scala 75:43 Counter.scala 97:11]
  reg  op1_buffer; // @[Reg.scala 15:16]
  reg  op2_buffer; // @[Reg.scala 15:16]
  reg  cond_buffer; // @[Reg.scala 15:16]
  reg  valid_buffer; // @[SE.scala 114:31]
  reg  ready_for_input; // @[SE.scala 117:38]
  wire  _GEN_185 = _T_1 & ready_for_input; // @[SE.scala 123:49 124:33 117:38]
  wire  _GEN_186 = 1'h1 & _GEN_185; // @[SE.scala 121:41 122:33]
  reg  mid_op1_buffer; // @[Reg.scala 15:16]
  wire  op1_reverse_1 = aes_invcipher_io_output_op1_14; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_0 = aes_invcipher_io_output_op1_15; // @[SE.scala 154:31 158:32]
  wire  lo_lo_lo = op1_reverse_1 & op1_reverse_0; // @[SE.scala 169:38]
  wire  op1_reverse_3 = aes_invcipher_io_output_op1_12; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_2 = aes_invcipher_io_output_op1_13; // @[SE.scala 154:31 158:32]
  wire  lo_lo_hi = op1_reverse_3 & op1_reverse_2; // @[SE.scala 169:38]
  wire  lo_lo = lo_lo_hi & lo_lo_lo; // @[SE.scala 169:38]
  wire  op1_reverse_5 = aes_invcipher_io_output_op1_10; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_4 = aes_invcipher_io_output_op1_11; // @[SE.scala 154:31 158:32]
  wire  lo_hi_lo = op1_reverse_5 & op1_reverse_4; // @[SE.scala 169:38]
  wire  op1_reverse_7 = aes_invcipher_io_output_op1_8; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_6 = aes_invcipher_io_output_op1_9; // @[SE.scala 154:31 158:32]
  wire  lo_hi_hi = op1_reverse_7 & op1_reverse_6; // @[SE.scala 169:38]
  wire  lo_hi = lo_hi_hi & lo_hi_lo; // @[SE.scala 169:38]
  wire  lo = lo_hi & lo_lo; // @[SE.scala 169:38]
  wire  op1_reverse_9 = aes_invcipher_io_output_op1_6; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_8 = aes_invcipher_io_output_op1_7; // @[SE.scala 154:31 158:32]
  wire  hi_lo_lo = op1_reverse_9 & op1_reverse_8; // @[SE.scala 169:38]
  wire  op1_reverse_11 = aes_invcipher_io_output_op1_4; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_10 = aes_invcipher_io_output_op1_5; // @[SE.scala 154:31 158:32]
  wire  hi_lo_hi = op1_reverse_11 & op1_reverse_10; // @[SE.scala 169:38]
  wire  hi_lo = hi_lo_hi & hi_lo_lo; // @[SE.scala 169:38]
  wire  op1_reverse_13 = aes_invcipher_io_output_op1_2; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_12 = aes_invcipher_io_output_op1_3; // @[SE.scala 154:31 158:32]
  wire  hi_hi_lo = op1_reverse_13 & op1_reverse_12; // @[SE.scala 169:38]
  wire  op1_reverse_15 = aes_invcipher_io_output_op1_0; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_14 = aes_invcipher_io_output_op1_1; // @[SE.scala 154:31 158:32]
  wire  hi_hi_hi = op1_reverse_15 & op1_reverse_14; // @[SE.scala 169:38]
  wire  hi_hi = hi_hi_hi & hi_hi_lo; // @[SE.scala 169:38]
  wire  hi = hi_hi & hi_lo; // @[SE.scala 169:38]
  wire  op1_asUInt = hi & lo; // @[SE.scala 169:38]
  wire  op2_reverse_1 = aes_invcipher_io_output_op2_14; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_0 = aes_invcipher_io_output_op2_15; // @[SE.scala 155:31 159:32]
  wire  lo_lo_lo_1 = op2_reverse_1 & op2_reverse_0; // @[SE.scala 170:38]
  wire  op2_reverse_3 = aes_invcipher_io_output_op2_12; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_2 = aes_invcipher_io_output_op2_13; // @[SE.scala 155:31 159:32]
  wire  lo_lo_hi_1 = op2_reverse_3 & op2_reverse_2; // @[SE.scala 170:38]
  wire  lo_lo_1 = lo_lo_hi_1 & lo_lo_lo_1; // @[SE.scala 170:38]
  wire  op2_reverse_5 = aes_invcipher_io_output_op2_10; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_4 = aes_invcipher_io_output_op2_11; // @[SE.scala 155:31 159:32]
  wire  lo_hi_lo_1 = op2_reverse_5 & op2_reverse_4; // @[SE.scala 170:38]
  wire  op2_reverse_7 = aes_invcipher_io_output_op2_8; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_6 = aes_invcipher_io_output_op2_9; // @[SE.scala 155:31 159:32]
  wire  lo_hi_hi_1 = op2_reverse_7 & op2_reverse_6; // @[SE.scala 170:38]
  wire  lo_hi_1 = lo_hi_hi_1 & lo_hi_lo_1; // @[SE.scala 170:38]
  wire  lo_1 = lo_hi_1 & lo_lo_1; // @[SE.scala 170:38]
  wire  op2_reverse_9 = aes_invcipher_io_output_op2_6; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_8 = aes_invcipher_io_output_op2_7; // @[SE.scala 155:31 159:32]
  wire  hi_lo_lo_1 = op2_reverse_9 & op2_reverse_8; // @[SE.scala 170:38]
  wire  op2_reverse_11 = aes_invcipher_io_output_op2_4; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_10 = aes_invcipher_io_output_op2_5; // @[SE.scala 155:31 159:32]
  wire  hi_lo_hi_1 = op2_reverse_11 & op2_reverse_10; // @[SE.scala 170:38]
  wire  hi_lo_1 = hi_lo_hi_1 & hi_lo_lo_1; // @[SE.scala 170:38]
  wire  op2_reverse_13 = aes_invcipher_io_output_op2_2; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_12 = aes_invcipher_io_output_op2_3; // @[SE.scala 155:31 159:32]
  wire  hi_hi_lo_1 = op2_reverse_13 & op2_reverse_12; // @[SE.scala 170:38]
  wire  op2_reverse_15 = aes_invcipher_io_output_op2_0; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_14 = aes_invcipher_io_output_op2_1; // @[SE.scala 155:31 159:32]
  wire  hi_hi_hi_1 = op2_reverse_15 & op2_reverse_14; // @[SE.scala 170:38]
  wire  hi_hi_1 = hi_hi_hi_1 & hi_hi_lo_1; // @[SE.scala 170:38]
  wire  hi_1 = hi_hi_1 & hi_lo_1; // @[SE.scala 170:38]
  wire  op2_asUInt = hi_1 & lo_1; // @[SE.scala 170:38]
  wire  _T_59 = mid_op1_buffer; // @[SE.scala 183:86]
  wire  _T_60 = op1_asUInt; // @[SE.scala 183:105]
  reg  result_valid_buffer; // @[SE.scala 188:42]
  wire  lo_lo_lo_lo_lo = prng_io_out_1 & prng_io_out_0; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_lo_hi = prng_io_out_3 & prng_io_out_2; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_lo = lo_lo_lo_lo_hi & lo_lo_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_hi_lo = prng_io_out_5 & prng_io_out_4; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_hi_hi = prng_io_out_7 & prng_io_out_6; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_hi = lo_lo_lo_hi_hi & lo_lo_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_3 = lo_lo_lo_hi & lo_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_lo_lo = prng_io_out_9 & prng_io_out_8; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_lo_hi = prng_io_out_11 & prng_io_out_10; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_lo = lo_lo_hi_lo_hi & lo_lo_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_hi_lo = prng_io_out_13 & prng_io_out_12; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_hi_hi = prng_io_out_15 & prng_io_out_14; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_hi = lo_lo_hi_hi_hi & lo_lo_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_3 = lo_lo_hi_hi & lo_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_3 = lo_lo_hi_3 & lo_lo_lo_3; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_lo_lo = prng_io_out_17 & prng_io_out_16; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_lo_hi = prng_io_out_19 & prng_io_out_18; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_lo = lo_hi_lo_lo_hi & lo_hi_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_hi_lo = prng_io_out_21 & prng_io_out_20; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_hi_hi = prng_io_out_23 & prng_io_out_22; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_hi = lo_hi_lo_hi_hi & lo_hi_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_3 = lo_hi_lo_hi & lo_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_lo_lo = prng_io_out_25 & prng_io_out_24; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_lo_hi = prng_io_out_27 & prng_io_out_26; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_lo = lo_hi_hi_lo_hi & lo_hi_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_hi_lo = prng_io_out_29 & prng_io_out_28; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_hi_hi = prng_io_out_31 & prng_io_out_30; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_hi = lo_hi_hi_hi_hi & lo_hi_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_3 = lo_hi_hi_hi & lo_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_3 = lo_hi_hi_3 & lo_hi_lo_3; // @[PRNG.scala 86:17]
  wire  lo_3 = lo_hi_3 & lo_lo_3; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_lo_lo = prng_io_out_33 & prng_io_out_32; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_lo_hi = prng_io_out_35 & prng_io_out_34; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_lo = hi_lo_lo_lo_hi & hi_lo_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_hi_lo = prng_io_out_37 & prng_io_out_36; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_hi_hi = prng_io_out_39 & prng_io_out_38; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_hi = hi_lo_lo_hi_hi & hi_lo_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_3 = hi_lo_lo_hi & hi_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_lo_lo = prng_io_out_41 & prng_io_out_40; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_lo_hi = prng_io_out_43 & prng_io_out_42; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_lo = hi_lo_hi_lo_hi & hi_lo_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_hi_lo = prng_io_out_45 & prng_io_out_44; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_hi_hi = prng_io_out_47 & prng_io_out_46; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_hi = hi_lo_hi_hi_hi & hi_lo_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_3 = hi_lo_hi_hi & hi_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_3 = hi_lo_hi_3 & hi_lo_lo_3; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_lo_lo = prng_io_out_49 & prng_io_out_48; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_lo_hi = prng_io_out_51 & prng_io_out_50; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_lo = hi_hi_lo_lo_hi & hi_hi_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_hi_lo = prng_io_out_53 & prng_io_out_52; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_hi_hi = prng_io_out_55 & prng_io_out_54; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_hi = hi_hi_lo_hi_hi & hi_hi_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_3 = hi_hi_lo_hi & hi_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_lo_lo = prng_io_out_57 & prng_io_out_56; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_lo_hi = prng_io_out_59 & prng_io_out_58; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_lo = hi_hi_hi_lo_hi & hi_hi_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_hi_lo = prng_io_out_61 & prng_io_out_60; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_hi_hi = prng_io_out_63 & prng_io_out_62; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_hi = hi_hi_hi_hi_hi & hi_hi_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_3 = hi_hi_hi_hi & hi_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_3 = hi_hi_hi_3 & hi_hi_lo_3; // @[PRNG.scala 86:17]
  wire  hi_3 = hi_hi_3 & hi_lo_3; // @[PRNG.scala 86:17]
  wire  bit64_randnum = hi_3 & lo_3; // @[PRNG.scala 86:17]
  wire  padded_result = seoperation_io_result & bit64_randnum; // @[Cat.scala 30:58]
  reg  result_buffer; // @[Reg.scala 15:16]
  wire  _GEN_190 = zero_cntr & 1'h1 & zero_cntr; // @[SE.scala 211:44 212:27 63:32]
  wire  _GEN_191 = mult_cntr & 1'h1 & mult_cntr; // @[SE.scala 214:56 215:27 64:32]
  wire  lo_lo_lo_4 = aes_cipher_io_output_text_1 & aes_cipher_io_output_text_0; // @[SE.scala 219:65]
  wire  lo_lo_hi_4 = aes_cipher_io_output_text_3 & aes_cipher_io_output_text_2; // @[SE.scala 219:65]
  wire  lo_lo_4 = lo_lo_hi_4 & lo_lo_lo_4; // @[SE.scala 219:65]
  wire  lo_hi_lo_4 = aes_cipher_io_output_text_5 & aes_cipher_io_output_text_4; // @[SE.scala 219:65]
  wire  lo_hi_hi_4 = aes_cipher_io_output_text_7 & aes_cipher_io_output_text_6; // @[SE.scala 219:65]
  wire  lo_hi_4 = lo_hi_hi_4 & lo_hi_lo_4; // @[SE.scala 219:65]
  wire  lo_4 = lo_hi_4 & lo_lo_4; // @[SE.scala 219:65]
  wire  hi_lo_lo_4 = aes_cipher_io_output_text_9 & aes_cipher_io_output_text_8; // @[SE.scala 219:65]
  wire  hi_lo_hi_4 = aes_cipher_io_output_text_11 & aes_cipher_io_output_text_10; // @[SE.scala 219:65]
  wire  hi_lo_4 = hi_lo_hi_4 & hi_lo_lo_4; // @[SE.scala 219:65]
  wire  hi_hi_lo_4 = aes_cipher_io_output_text_13 & aes_cipher_io_output_text_12; // @[SE.scala 219:65]
  wire  hi_hi_hi_4 = aes_cipher_io_output_text_15 & aes_cipher_io_output_text_14; // @[SE.scala 219:65]
  wire  hi_hi_4 = hi_hi_hi_4 & hi_hi_lo_4; // @[SE.scala 219:65]
  wire  hi_4 = hi_hi_4 & hi_lo_4; // @[SE.scala 219:65]
  wire  _T_89 = hi_4 & lo_4; // @[SE.scala 219:65]
  reg  output_buffer; // @[Reg.scala 15:16]
  reg  output_valid; // @[SE.scala 220:35]
  wire  _GEN_193 = 1'h1 & output_valid; // @[SE.scala 224:49 225:30 220:35]
  wire  _GEN_194 = aes_cipher_io_output_valid & _GEN_193; // @[SE.scala 222:41 223:30]
  SEOperation seoperation ( // @[SE.scala 83:33]
    .io_op1_input(seoperation_io_op1_input),
    .io_op2_input(seoperation_io_op2_input),
    .io_result(seoperation_io_result)
  );
  AESDecrypt aes_invcipher ( // @[SE.scala 84:35]
    .clock(aes_invcipher_clock),
    .io_input_valid(aes_invcipher_io_input_valid),
    .io_input_op1_0(aes_invcipher_io_input_op1_0),
    .io_input_op1_1(aes_invcipher_io_input_op1_1),
    .io_input_op1_2(aes_invcipher_io_input_op1_2),
    .io_input_op1_3(aes_invcipher_io_input_op1_3),
    .io_input_op1_4(aes_invcipher_io_input_op1_4),
    .io_input_op1_5(aes_invcipher_io_input_op1_5),
    .io_input_op1_6(aes_invcipher_io_input_op1_6),
    .io_input_op1_7(aes_invcipher_io_input_op1_7),
    .io_input_op1_8(aes_invcipher_io_input_op1_8),
    .io_input_op1_9(aes_invcipher_io_input_op1_9),
    .io_input_op1_10(aes_invcipher_io_input_op1_10),
    .io_input_op1_11(aes_invcipher_io_input_op1_11),
    .io_input_op1_12(aes_invcipher_io_input_op1_12),
    .io_input_op1_13(aes_invcipher_io_input_op1_13),
    .io_input_op1_14(aes_invcipher_io_input_op1_14),
    .io_input_op1_15(aes_invcipher_io_input_op1_15),
    .io_input_op2_0(aes_invcipher_io_input_op2_0),
    .io_input_op2_1(aes_invcipher_io_input_op2_1),
    .io_input_op2_2(aes_invcipher_io_input_op2_2),
    .io_input_op2_3(aes_invcipher_io_input_op2_3),
    .io_input_op2_4(aes_invcipher_io_input_op2_4),
    .io_input_op2_5(aes_invcipher_io_input_op2_5),
    .io_input_op2_6(aes_invcipher_io_input_op2_6),
    .io_input_op2_7(aes_invcipher_io_input_op2_7),
    .io_input_op2_8(aes_invcipher_io_input_op2_8),
    .io_input_op2_9(aes_invcipher_io_input_op2_9),
    .io_input_op2_10(aes_invcipher_io_input_op2_10),
    .io_input_op2_11(aes_invcipher_io_input_op2_11),
    .io_input_op2_12(aes_invcipher_io_input_op2_12),
    .io_input_op2_13(aes_invcipher_io_input_op2_13),
    .io_input_op2_14(aes_invcipher_io_input_op2_14),
    .io_input_op2_15(aes_invcipher_io_input_op2_15),
    .io_input_cond_0(aes_invcipher_io_input_cond_0),
    .io_input_cond_1(aes_invcipher_io_input_cond_1),
    .io_input_cond_2(aes_invcipher_io_input_cond_2),
    .io_input_cond_3(aes_invcipher_io_input_cond_3),
    .io_input_cond_4(aes_invcipher_io_input_cond_4),
    .io_input_cond_5(aes_invcipher_io_input_cond_5),
    .io_input_cond_6(aes_invcipher_io_input_cond_6),
    .io_input_cond_7(aes_invcipher_io_input_cond_7),
    .io_input_cond_8(aes_invcipher_io_input_cond_8),
    .io_input_cond_9(aes_invcipher_io_input_cond_9),
    .io_input_cond_10(aes_invcipher_io_input_cond_10),
    .io_input_cond_11(aes_invcipher_io_input_cond_11),
    .io_input_cond_12(aes_invcipher_io_input_cond_12),
    .io_input_cond_13(aes_invcipher_io_input_cond_13),
    .io_input_cond_14(aes_invcipher_io_input_cond_14),
    .io_input_cond_15(aes_invcipher_io_input_cond_15),
    .io_output_op1_0(aes_invcipher_io_output_op1_0),
    .io_output_op1_1(aes_invcipher_io_output_op1_1),
    .io_output_op1_2(aes_invcipher_io_output_op1_2),
    .io_output_op1_3(aes_invcipher_io_output_op1_3),
    .io_output_op1_4(aes_invcipher_io_output_op1_4),
    .io_output_op1_5(aes_invcipher_io_output_op1_5),
    .io_output_op1_6(aes_invcipher_io_output_op1_6),
    .io_output_op1_7(aes_invcipher_io_output_op1_7),
    .io_output_op1_8(aes_invcipher_io_output_op1_8),
    .io_output_op1_9(aes_invcipher_io_output_op1_9),
    .io_output_op1_10(aes_invcipher_io_output_op1_10),
    .io_output_op1_11(aes_invcipher_io_output_op1_11),
    .io_output_op1_12(aes_invcipher_io_output_op1_12),
    .io_output_op1_13(aes_invcipher_io_output_op1_13),
    .io_output_op1_14(aes_invcipher_io_output_op1_14),
    .io_output_op1_15(aes_invcipher_io_output_op1_15),
    .io_output_op2_0(aes_invcipher_io_output_op2_0),
    .io_output_op2_1(aes_invcipher_io_output_op2_1),
    .io_output_op2_2(aes_invcipher_io_output_op2_2),
    .io_output_op2_3(aes_invcipher_io_output_op2_3),
    .io_output_op2_4(aes_invcipher_io_output_op2_4),
    .io_output_op2_5(aes_invcipher_io_output_op2_5),
    .io_output_op2_6(aes_invcipher_io_output_op2_6),
    .io_output_op2_7(aes_invcipher_io_output_op2_7),
    .io_output_op2_8(aes_invcipher_io_output_op2_8),
    .io_output_op2_9(aes_invcipher_io_output_op2_9),
    .io_output_op2_10(aes_invcipher_io_output_op2_10),
    .io_output_op2_11(aes_invcipher_io_output_op2_11),
    .io_output_op2_12(aes_invcipher_io_output_op2_12),
    .io_output_op2_13(aes_invcipher_io_output_op2_13),
    .io_output_op2_14(aes_invcipher_io_output_op2_14),
    .io_output_op2_15(aes_invcipher_io_output_op2_15),
    .io_output_valid(aes_invcipher_io_output_valid)
  );
  AESEncrypt aes_cipher ( // @[SE.scala 85:32]
    .clock(aes_cipher_clock),
    .io_input_valid(aes_cipher_io_input_valid),
    .io_input_text_0(aes_cipher_io_input_text_0),
    .io_input_text_1(aes_cipher_io_input_text_1),
    .io_input_text_2(aes_cipher_io_input_text_2),
    .io_input_text_3(aes_cipher_io_input_text_3),
    .io_input_text_4(aes_cipher_io_input_text_4),
    .io_input_text_5(aes_cipher_io_input_text_5),
    .io_input_text_6(aes_cipher_io_input_text_6),
    .io_input_text_7(aes_cipher_io_input_text_7),
    .io_input_text_8(aes_cipher_io_input_text_8),
    .io_input_text_9(aes_cipher_io_input_text_9),
    .io_input_text_10(aes_cipher_io_input_text_10),
    .io_input_text_11(aes_cipher_io_input_text_11),
    .io_input_text_12(aes_cipher_io_input_text_12),
    .io_input_text_13(aes_cipher_io_input_text_13),
    .io_input_text_14(aes_cipher_io_input_text_14),
    .io_input_text_15(aes_cipher_io_input_text_15),
    .io_output_text_0(aes_cipher_io_output_text_0),
    .io_output_text_1(aes_cipher_io_output_text_1),
    .io_output_text_2(aes_cipher_io_output_text_2),
    .io_output_text_3(aes_cipher_io_output_text_3),
    .io_output_text_4(aes_cipher_io_output_text_4),
    .io_output_text_5(aes_cipher_io_output_text_5),
    .io_output_text_6(aes_cipher_io_output_text_6),
    .io_output_text_7(aes_cipher_io_output_text_7),
    .io_output_text_8(aes_cipher_io_output_text_8),
    .io_output_text_9(aes_cipher_io_output_text_9),
    .io_output_text_10(aes_cipher_io_output_text_10),
    .io_output_text_11(aes_cipher_io_output_text_11),
    .io_output_text_12(aes_cipher_io_output_text_12),
    .io_output_text_13(aes_cipher_io_output_text_13),
    .io_output_text_14(aes_cipher_io_output_text_14),
    .io_output_text_15(aes_cipher_io_output_text_15),
    .io_output_intermediate(aes_cipher_io_output_intermediate),
    .io_output_valid(aes_cipher_io_output_valid)
  );
  MaxPeriodFibonacciLFSR prng ( // @[PRNG.scala 82:22]
    .clock(prng_clock),
    .reset(prng_reset),
    .io_out_0(prng_io_out_0),
    .io_out_1(prng_io_out_1),
    .io_out_2(prng_io_out_2),
    .io_out_3(prng_io_out_3),
    .io_out_4(prng_io_out_4),
    .io_out_5(prng_io_out_5),
    .io_out_6(prng_io_out_6),
    .io_out_7(prng_io_out_7),
    .io_out_8(prng_io_out_8),
    .io_out_9(prng_io_out_9),
    .io_out_10(prng_io_out_10),
    .io_out_11(prng_io_out_11),
    .io_out_12(prng_io_out_12),
    .io_out_13(prng_io_out_13),
    .io_out_14(prng_io_out_14),
    .io_out_15(prng_io_out_15),
    .io_out_16(prng_io_out_16),
    .io_out_17(prng_io_out_17),
    .io_out_18(prng_io_out_18),
    .io_out_19(prng_io_out_19),
    .io_out_20(prng_io_out_20),
    .io_out_21(prng_io_out_21),
    .io_out_22(prng_io_out_22),
    .io_out_23(prng_io_out_23),
    .io_out_24(prng_io_out_24),
    .io_out_25(prng_io_out_25),
    .io_out_26(prng_io_out_26),
    .io_out_27(prng_io_out_27),
    .io_out_28(prng_io_out_28),
    .io_out_29(prng_io_out_29),
    .io_out_30(prng_io_out_30),
    .io_out_31(prng_io_out_31),
    .io_out_32(prng_io_out_32),
    .io_out_33(prng_io_out_33),
    .io_out_34(prng_io_out_34),
    .io_out_35(prng_io_out_35),
    .io_out_36(prng_io_out_36),
    .io_out_37(prng_io_out_37),
    .io_out_38(prng_io_out_38),
    .io_out_39(prng_io_out_39),
    .io_out_40(prng_io_out_40),
    .io_out_41(prng_io_out_41),
    .io_out_42(prng_io_out_42),
    .io_out_43(prng_io_out_43),
    .io_out_44(prng_io_out_44),
    .io_out_45(prng_io_out_45),
    .io_out_46(prng_io_out_46),
    .io_out_47(prng_io_out_47),
    .io_out_48(prng_io_out_48),
    .io_out_49(prng_io_out_49),
    .io_out_50(prng_io_out_50),
    .io_out_51(prng_io_out_51),
    .io_out_52(prng_io_out_52),
    .io_out_53(prng_io_out_53),
    .io_out_54(prng_io_out_54),
    .io_out_55(prng_io_out_55),
    .io_out_56(prng_io_out_56),
    .io_out_57(prng_io_out_57),
    .io_out_58(prng_io_out_58),
    .io_out_59(prng_io_out_59),
    .io_out_60(prng_io_out_60),
    .io_out_61(prng_io_out_61),
    .io_out_62(prng_io_out_62),
    .io_out_63(prng_io_out_63)
  );
  assign io_in_ready = ready_for_input; // @[SE.scala 118:21]
  assign io_out_result = output_buffer; // @[SE.scala 228:23]
  assign io_out_valid = output_valid; // @[SE.scala 227:22]
  assign io_out_cntr = value; // @[SE.scala 78:21]
  assign io_out_zero_cntr = zero_cntr; // @[SE.scala 65:26]
  assign io_out_mult_cntr = mult_cntr; // @[SE.scala 66:26]
  assign io_out_intermediate = aes_cipher_io_output_intermediate; // @[SE.scala 217:29]
  assign seoperation_io_op1_input = _T_59 & _T_60; // @[SE.scala 183:40]
  assign seoperation_io_op2_input = op2_asUInt; // @[SE.scala 184:47]
  assign aes_invcipher_clock = clock;
  assign aes_invcipher_io_input_valid = valid_buffer; // @[SE.scala 150:38]
  assign aes_invcipher_io_input_op1_0 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_1 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_2 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_3 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_4 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_5 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_6 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_7 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_8 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_9 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_10 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_11 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_12 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_13 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_14 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op1_15 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op2_0 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_1 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_2 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_3 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_4 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_5 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_6 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_7 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_8 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_9 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_10 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_11 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_12 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_13 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_14 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_op2_15 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_cond_0 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_1 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_2 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_3 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_4 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_5 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_6 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_7 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_8 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_9 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_10 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_11 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_12 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_13 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_14 = cond_buffer; // @[SE.scala 148:60]
  assign aes_invcipher_io_input_cond_15 = cond_buffer; // @[SE.scala 148:60]
  assign aes_cipher_clock = clock;
  assign aes_cipher_io_input_valid = result_valid_buffer; // @[SE.scala 209:35]
  assign aes_cipher_io_input_text_0 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_1 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_2 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_3 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_4 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_5 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_6 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_7 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_8 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_9 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_10 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_11 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_12 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_13 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_14 = result_buffer; // @[SE.scala 203:47]
  assign aes_cipher_io_input_text_15 = result_buffer; // @[SE.scala 203:47]
  assign prng_clock = clock;
  assign prng_reset = reset;
  always @(posedge clock) begin
    value <= 1'h1 & _GEN_4; // @[Counter.scala 60:{40,40}]
    zero_cntr <= 1'h1 & _GEN_190; // @[SE.scala 63:{32,32}]
    mult_cntr <= 1'h1 & _GEN_191; // @[SE.scala 64:{32,32}]
    op1_buffer <= io_in_op1 & op1_buffer; // @[Reg.scala 15:16 16:{19,23}]
    op2_buffer <= io_in_op2 & op2_buffer; // @[Reg.scala 15:16 16:{19,23}]
    cond_buffer <= io_in_cond & cond_buffer; // @[Reg.scala 15:16 16:{19,23}]
    valid_buffer <= _T & (1'h1 & valid_buffer); // @[SE.scala 120:28]
    ready_for_input <= reset & _GEN_186; // @[SE.scala 117:{38,38}]
    mid_op1_buffer <= op1_buffer & mid_op1_buffer; // @[Reg.scala 15:16 16:{19,23}]
    result_valid_buffer <= aes_invcipher_io_output_valid & (1'h1 & result_valid_buffer); // @[SE.scala 189:37]
    result_buffer <= padded_result & result_buffer; // @[Reg.scala 15:16 16:{19,23}]
    output_buffer <= _T_89 & output_buffer; // @[Reg.scala 15:16 16:{19,23}]
    output_valid <= 1'h1 & _GEN_194; // @[SE.scala 220:{35,35}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  zero_cntr = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mult_cntr = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  op1_buffer = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  op2_buffer = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cond_buffer = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_buffer = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ready_for_input = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mid_op1_buffer = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  result_valid_buffer = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  result_buffer = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_buffer = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_valid = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
