module Crc64 (
    input [63:0] crcIn,
    input [63:0] data,
    output [63:0] crcOut
);
    assign crcOut[0] = crcIn[1] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[15] ^ crcIn[18] ^ crcIn[22] ^ crcIn[23] ^ crcIn[26] ^ crcIn[27] ^ crcIn[29] ^ crcIn[30] ^ crcIn[36] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[43] ^ crcIn[45] ^ crcIn[48] ^ crcIn[50] ^ crcIn[51] ^ crcIn[55] ^ crcIn[56] ^ crcIn[57] ^ crcIn[58] ^ crcIn[60] ^ crcIn[62] ^ data[1] ^ data[4] ^ data[5] ^ data[6] ^ data[11] ^ data[12] ^ data[13] ^ data[14] ^ data[15] ^ data[18] ^ data[22] ^ data[23] ^ data[26] ^ data[27] ^ data[29] ^ data[30] ^ data[36] ^ data[38] ^ data[39] ^ data[40] ^ data[43] ^ data[45] ^ data[48] ^ data[50] ^ data[51] ^ data[55] ^ data[56] ^ data[57] ^ data[58] ^ data[60] ^ data[62];
    assign crcOut[1] = crcIn[2] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[15] ^ crcIn[16] ^ crcIn[19] ^ crcIn[23] ^ crcIn[24] ^ crcIn[27] ^ crcIn[28] ^ crcIn[30] ^ crcIn[31] ^ crcIn[37] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[44] ^ crcIn[46] ^ crcIn[49] ^ crcIn[51] ^ crcIn[52] ^ crcIn[56] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[63] ^ data[2] ^ data[5] ^ data[6] ^ data[7] ^ data[12] ^ data[13] ^ data[14] ^ data[15] ^ data[16] ^ data[19] ^ data[23] ^ data[24] ^ data[27] ^ data[28] ^ data[30] ^ data[31] ^ data[37] ^ data[39] ^ data[40] ^ data[41] ^ data[44] ^ data[46] ^ data[49] ^ data[51] ^ data[52] ^ data[56] ^ data[57] ^ data[58] ^ data[59] ^ data[61] ^ data[63];
    assign crcOut[2] = crcIn[1] ^ crcIn[3] ^ crcIn[4] ^ crcIn[5] ^ crcIn[7] ^ crcIn[8] ^ crcIn[11] ^ crcIn[12] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[20] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[36] ^ crcIn[39] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[47] ^ crcIn[48] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[55] ^ crcIn[56] ^ crcIn[59] ^ data[1] ^ data[3] ^ data[4] ^ data[5] ^ data[7] ^ data[8] ^ data[11] ^ data[12] ^ data[16] ^ data[17] ^ data[18] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[28] ^ data[30] ^ data[31] ^ data[32] ^ data[36] ^ data[39] ^ data[41] ^ data[42] ^ data[43] ^ data[47] ^ data[48] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[56] ^ data[59];
    assign crcOut[3] = crcIn[2] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[8] ^ crcIn[9] ^ crcIn[12] ^ crcIn[13] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[21] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[37] ^ crcIn[40] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[48] ^ crcIn[49] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[57] ^ crcIn[60] ^ data[2] ^ data[4] ^ data[5] ^ data[6] ^ data[8] ^ data[9] ^ data[12] ^ data[13] ^ data[17] ^ data[18] ^ data[19] ^ data[21] ^ data[23] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[31] ^ data[32] ^ data[33] ^ data[37] ^ data[40] ^ data[42] ^ data[43] ^ data[44] ^ data[48] ^ data[49] ^ data[52] ^ data[53] ^ data[54] ^ data[56] ^ data[57] ^ data[60];
    assign crcOut[4] = crcIn[3] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[9] ^ crcIn[10] ^ crcIn[13] ^ crcIn[14] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[22] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[38] ^ crcIn[41] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[49] ^ crcIn[50] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[57] ^ crcIn[58] ^ crcIn[61] ^ data[3] ^ data[5] ^ data[6] ^ data[7] ^ data[9] ^ data[10] ^ data[13] ^ data[14] ^ data[18] ^ data[19] ^ data[20] ^ data[22] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[30] ^ data[32] ^ data[33] ^ data[34] ^ data[38] ^ data[41] ^ data[43] ^ data[44] ^ data[45] ^ data[49] ^ data[50] ^ data[53] ^ data[54] ^ data[55] ^ data[57] ^ data[58] ^ data[61];
    assign crcOut[5] = crcIn[4] ^ crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[10] ^ crcIn[11] ^ crcIn[14] ^ crcIn[15] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[23] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[39] ^ crcIn[42] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[50] ^ crcIn[51] ^ crcIn[54] ^ crcIn[55] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[62] ^ data[4] ^ data[6] ^ data[7] ^ data[8] ^ data[10] ^ data[11] ^ data[14] ^ data[15] ^ data[19] ^ data[20] ^ data[21] ^ data[23] ^ data[25] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[30] ^ data[31] ^ data[33] ^ data[34] ^ data[35] ^ data[39] ^ data[42] ^ data[44] ^ data[45] ^ data[46] ^ data[50] ^ data[51] ^ data[54] ^ data[55] ^ data[56] ^ data[58] ^ data[59] ^ data[62];
    assign crcOut[6] = crcIn[0] ^ crcIn[5] ^ crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[11] ^ crcIn[12] ^ crcIn[15] ^ crcIn[16] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[24] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[40] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[51] ^ crcIn[52] ^ crcIn[55] ^ crcIn[56] ^ crcIn[57] ^ crcIn[59] ^ crcIn[60] ^ crcIn[63] ^ data[0] ^ data[5] ^ data[7] ^ data[8] ^ data[9] ^ data[11] ^ data[12] ^ data[15] ^ data[16] ^ data[20] ^ data[21] ^ data[22] ^ data[24] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[34] ^ data[35] ^ data[36] ^ data[40] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[51] ^ data[52] ^ data[55] ^ data[56] ^ data[57] ^ data[59] ^ data[60] ^ data[63];
    assign crcOut[7] = crcIn[4] ^ crcIn[5] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[14] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[21] ^ crcIn[25] ^ crcIn[26] ^ crcIn[28] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[35] ^ crcIn[37] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[55] ^ crcIn[61] ^ crcIn[62] ^ data[4] ^ data[5] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[14] ^ data[15] ^ data[16] ^ data[17] ^ data[18] ^ data[21] ^ data[25] ^ data[26] ^ data[28] ^ data[31] ^ data[32] ^ data[33] ^ data[35] ^ data[37] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[47] ^ data[50] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[61] ^ data[62];
    assign crcOut[8] = crcIn[0] ^ crcIn[5] ^ crcIn[6] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[22] ^ crcIn[26] ^ crcIn[27] ^ crcIn[29] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[36] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[5] ^ data[6] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[15] ^ data[16] ^ data[17] ^ data[18] ^ data[19] ^ data[22] ^ data[26] ^ data[27] ^ data[29] ^ data[32] ^ data[33] ^ data[34] ^ data[36] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[44] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[51] ^ data[52] ^ data[53] ^ data[54] ^ data[56] ^ data[62] ^ data[63];
    assign crcOut[9] = crcIn[0] ^ crcIn[4] ^ crcIn[5] ^ crcIn[7] ^ crcIn[10] ^ crcIn[14] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[19] ^ crcIn[20] ^ crcIn[22] ^ crcIn[26] ^ crcIn[28] ^ crcIn[29] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[37] ^ crcIn[38] ^ crcIn[41] ^ crcIn[42] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[60] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[4] ^ data[5] ^ data[7] ^ data[10] ^ data[14] ^ data[15] ^ data[16] ^ data[17] ^ data[19] ^ data[20] ^ data[22] ^ data[26] ^ data[28] ^ data[29] ^ data[33] ^ data[34] ^ data[35] ^ data[36] ^ data[37] ^ data[38] ^ data[41] ^ data[42] ^ data[46] ^ data[47] ^ data[49] ^ data[50] ^ data[51] ^ data[52] ^ data[53] ^ data[54] ^ data[56] ^ data[58] ^ data[60] ^ data[62] ^ data[63];
    assign crcOut[10] = crcIn[0] ^ crcIn[4] ^ crcIn[8] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[16] ^ crcIn[17] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[26] ^ crcIn[34] ^ crcIn[35] ^ crcIn[37] ^ crcIn[40] ^ crcIn[42] ^ crcIn[45] ^ crcIn[47] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[4] ^ data[8] ^ data[12] ^ data[13] ^ data[14] ^ data[16] ^ data[17] ^ data[20] ^ data[21] ^ data[22] ^ data[26] ^ data[34] ^ data[35] ^ data[37] ^ data[40] ^ data[42] ^ data[45] ^ data[47] ^ data[52] ^ data[53] ^ data[54] ^ data[56] ^ data[58] ^ data[59] ^ data[60] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[11] = crcIn[0] ^ crcIn[4] ^ crcIn[6] ^ crcIn[9] ^ crcIn[11] ^ crcIn[12] ^ crcIn[17] ^ crcIn[21] ^ crcIn[26] ^ crcIn[29] ^ crcIn[30] ^ crcIn[35] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[45] ^ crcIn[46] ^ crcIn[50] ^ crcIn[51] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[63] ^ data[0] ^ data[4] ^ data[6] ^ data[9] ^ data[11] ^ data[12] ^ data[17] ^ data[21] ^ data[26] ^ data[29] ^ data[30] ^ data[35] ^ data[39] ^ data[40] ^ data[41] ^ data[45] ^ data[46] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[56] ^ data[58] ^ data[59] ^ data[61] ^ data[63];
    assign crcOut[12] = crcIn[0] ^ crcIn[4] ^ crcIn[6] ^ crcIn[7] ^ crcIn[10] ^ crcIn[11] ^ crcIn[14] ^ crcIn[15] ^ crcIn[23] ^ crcIn[26] ^ crcIn[29] ^ crcIn[31] ^ crcIn[38] ^ crcIn[39] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[50] ^ crcIn[52] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ data[0] ^ data[4] ^ data[6] ^ data[7] ^ data[10] ^ data[11] ^ data[14] ^ data[15] ^ data[23] ^ data[26] ^ data[29] ^ data[31] ^ data[38] ^ data[39] ^ data[41] ^ data[42] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[50] ^ data[52] ^ data[54] ^ data[56] ^ data[58] ^ data[59];
    assign crcOut[13] = crcIn[1] ^ crcIn[5] ^ crcIn[7] ^ crcIn[8] ^ crcIn[11] ^ crcIn[12] ^ crcIn[15] ^ crcIn[16] ^ crcIn[24] ^ crcIn[27] ^ crcIn[30] ^ crcIn[32] ^ crcIn[39] ^ crcIn[40] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[51] ^ crcIn[53] ^ crcIn[55] ^ crcIn[57] ^ crcIn[59] ^ crcIn[60] ^ data[1] ^ data[5] ^ data[7] ^ data[8] ^ data[11] ^ data[12] ^ data[15] ^ data[16] ^ data[24] ^ data[27] ^ data[30] ^ data[32] ^ data[39] ^ data[40] ^ data[42] ^ data[43] ^ data[44] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[51] ^ data[53] ^ data[55] ^ data[57] ^ data[59] ^ data[60];
    assign crcOut[14] = crcIn[0] ^ crcIn[2] ^ crcIn[6] ^ crcIn[8] ^ crcIn[9] ^ crcIn[12] ^ crcIn[13] ^ crcIn[16] ^ crcIn[17] ^ crcIn[25] ^ crcIn[28] ^ crcIn[31] ^ crcIn[33] ^ crcIn[40] ^ crcIn[41] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[52] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[60] ^ crcIn[61] ^ data[0] ^ data[2] ^ data[6] ^ data[8] ^ data[9] ^ data[12] ^ data[13] ^ data[16] ^ data[17] ^ data[25] ^ data[28] ^ data[31] ^ data[33] ^ data[40] ^ data[41] ^ data[43] ^ data[44] ^ data[45] ^ data[47] ^ data[48] ^ data[49] ^ data[50] ^ data[52] ^ data[54] ^ data[56] ^ data[58] ^ data[60] ^ data[61];
    assign crcOut[15] = crcIn[1] ^ crcIn[3] ^ crcIn[7] ^ crcIn[9] ^ crcIn[10] ^ crcIn[13] ^ crcIn[14] ^ crcIn[17] ^ crcIn[18] ^ crcIn[26] ^ crcIn[29] ^ crcIn[32] ^ crcIn[34] ^ crcIn[41] ^ crcIn[42] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[51] ^ crcIn[53] ^ crcIn[55] ^ crcIn[57] ^ crcIn[59] ^ crcIn[61] ^ crcIn[62] ^ data[1] ^ data[3] ^ data[7] ^ data[9] ^ data[10] ^ data[13] ^ data[14] ^ data[17] ^ data[18] ^ data[26] ^ data[29] ^ data[32] ^ data[34] ^ data[41] ^ data[42] ^ data[44] ^ data[45] ^ data[46] ^ data[48] ^ data[49] ^ data[50] ^ data[51] ^ data[53] ^ data[55] ^ data[57] ^ data[59] ^ data[61] ^ data[62];
    assign crcOut[16] = crcIn[0] ^ crcIn[2] ^ crcIn[4] ^ crcIn[8] ^ crcIn[10] ^ crcIn[11] ^ crcIn[14] ^ crcIn[15] ^ crcIn[18] ^ crcIn[19] ^ crcIn[27] ^ crcIn[30] ^ crcIn[33] ^ crcIn[35] ^ crcIn[42] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[60] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[2] ^ data[4] ^ data[8] ^ data[10] ^ data[11] ^ data[14] ^ data[15] ^ data[18] ^ data[19] ^ data[27] ^ data[30] ^ data[33] ^ data[35] ^ data[42] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[49] ^ data[50] ^ data[51] ^ data[52] ^ data[54] ^ data[56] ^ data[58] ^ data[60] ^ data[62] ^ data[63];
    assign crcOut[17] = crcIn[0] ^ crcIn[3] ^ crcIn[4] ^ crcIn[6] ^ crcIn[9] ^ crcIn[13] ^ crcIn[14] ^ crcIn[16] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[22] ^ crcIn[23] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[34] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[52] ^ crcIn[53] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[3] ^ data[4] ^ data[6] ^ data[9] ^ data[13] ^ data[14] ^ data[16] ^ data[18] ^ data[19] ^ data[20] ^ data[22] ^ data[23] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[30] ^ data[31] ^ data[34] ^ data[38] ^ data[39] ^ data[40] ^ data[44] ^ data[45] ^ data[46] ^ data[47] ^ data[52] ^ data[53] ^ data[56] ^ data[58] ^ data[59] ^ data[60] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[18] = crcIn[0] ^ crcIn[6] ^ crcIn[7] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[24] ^ crcIn[26] ^ crcIn[28] ^ crcIn[31] ^ crcIn[32] ^ crcIn[35] ^ crcIn[36] ^ crcIn[38] ^ crcIn[41] ^ crcIn[43] ^ crcIn[46] ^ crcIn[47] ^ crcIn[50] ^ crcIn[51] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[63] ^ data[0] ^ data[6] ^ data[7] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[17] ^ data[18] ^ data[19] ^ data[20] ^ data[21] ^ data[22] ^ data[24] ^ data[26] ^ data[28] ^ data[31] ^ data[32] ^ data[35] ^ data[36] ^ data[38] ^ data[41] ^ data[43] ^ data[46] ^ data[47] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[55] ^ data[56] ^ data[58] ^ data[59] ^ data[61] ^ data[63];
    assign crcOut[19] = crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[15] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[25] ^ crcIn[26] ^ crcIn[30] ^ crcIn[32] ^ crcIn[33] ^ crcIn[37] ^ crcIn[38] ^ crcIn[40] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[47] ^ crcIn[50] ^ crcIn[52] ^ crcIn[54] ^ crcIn[58] ^ crcIn[59] ^ data[4] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[15] ^ data[19] ^ data[20] ^ data[21] ^ data[25] ^ data[26] ^ data[30] ^ data[32] ^ data[33] ^ data[37] ^ data[38] ^ data[40] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[47] ^ data[50] ^ data[52] ^ data[54] ^ data[58] ^ data[59];
    assign crcOut[20] = crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[16] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[26] ^ crcIn[27] ^ crcIn[31] ^ crcIn[33] ^ crcIn[34] ^ crcIn[38] ^ crcIn[39] ^ crcIn[41] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[51] ^ crcIn[53] ^ crcIn[55] ^ crcIn[59] ^ crcIn[60] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[16] ^ data[20] ^ data[21] ^ data[22] ^ data[26] ^ data[27] ^ data[31] ^ data[33] ^ data[34] ^ data[38] ^ data[39] ^ data[41] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[48] ^ data[51] ^ data[53] ^ data[55] ^ data[59] ^ data[60];
    assign crcOut[21] = crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[17] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[27] ^ crcIn[28] ^ crcIn[32] ^ crcIn[34] ^ crcIn[35] ^ crcIn[39] ^ crcIn[40] ^ crcIn[42] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[52] ^ crcIn[54] ^ crcIn[56] ^ crcIn[60] ^ crcIn[61] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[17] ^ data[21] ^ data[22] ^ data[23] ^ data[27] ^ data[28] ^ data[32] ^ data[34] ^ data[35] ^ data[39] ^ data[40] ^ data[42] ^ data[44] ^ data[45] ^ data[46] ^ data[47] ^ data[49] ^ data[52] ^ data[54] ^ data[56] ^ data[60] ^ data[61];
    assign crcOut[22] = crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[18] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[28] ^ crcIn[29] ^ crcIn[33] ^ crcIn[35] ^ crcIn[36] ^ crcIn[40] ^ crcIn[41] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[50] ^ crcIn[53] ^ crcIn[55] ^ crcIn[57] ^ crcIn[61] ^ crcIn[62] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[18] ^ data[22] ^ data[23] ^ data[24] ^ data[28] ^ data[29] ^ data[33] ^ data[35] ^ data[36] ^ data[40] ^ data[41] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[50] ^ data[53] ^ data[55] ^ data[57] ^ data[61] ^ data[62];
    assign crcOut[23] = crcIn[0] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[19] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[29] ^ crcIn[30] ^ crcIn[34] ^ crcIn[36] ^ crcIn[37] ^ crcIn[41] ^ crcIn[42] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[51] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[19] ^ data[23] ^ data[24] ^ data[25] ^ data[29] ^ data[30] ^ data[34] ^ data[36] ^ data[37] ^ data[41] ^ data[42] ^ data[44] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[51] ^ data[54] ^ data[56] ^ data[58] ^ data[62] ^ data[63];
    assign crcOut[24] = crcIn[0] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[9] ^ crcIn[10] ^ crcIn[14] ^ crcIn[15] ^ crcIn[18] ^ crcIn[20] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[27] ^ crcIn[29] ^ crcIn[31] ^ crcIn[35] ^ crcIn[36] ^ crcIn[37] ^ crcIn[39] ^ crcIn[40] ^ crcIn[42] ^ crcIn[47] ^ crcIn[49] ^ crcIn[51] ^ crcIn[52] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[4] ^ data[5] ^ data[6] ^ data[9] ^ data[10] ^ data[14] ^ data[15] ^ data[18] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[25] ^ data[27] ^ data[29] ^ data[31] ^ data[35] ^ data[36] ^ data[37] ^ data[39] ^ data[40] ^ data[42] ^ data[47] ^ data[49] ^ data[51] ^ data[52] ^ data[56] ^ data[58] ^ data[59] ^ data[60] ^ data[62] ^ data[63];
    assign crcOut[25] = crcIn[0] ^ crcIn[4] ^ crcIn[7] ^ crcIn[10] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[16] ^ crcIn[18] ^ crcIn[19] ^ crcIn[21] ^ crcIn[22] ^ crcIn[24] ^ crcIn[25] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[32] ^ crcIn[37] ^ crcIn[39] ^ crcIn[41] ^ crcIn[45] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[55] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[4] ^ data[7] ^ data[10] ^ data[12] ^ data[13] ^ data[14] ^ data[16] ^ data[18] ^ data[19] ^ data[21] ^ data[22] ^ data[24] ^ data[25] ^ data[27] ^ data[28] ^ data[29] ^ data[32] ^ data[37] ^ data[39] ^ data[41] ^ data[45] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[56] ^ data[58] ^ data[59] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[26] = crcIn[0] ^ crcIn[4] ^ crcIn[6] ^ crcIn[8] ^ crcIn[12] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[25] ^ crcIn[27] ^ crcIn[28] ^ crcIn[33] ^ crcIn[36] ^ crcIn[39] ^ crcIn[42] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[58] ^ crcIn[59] ^ crcIn[63] ^ data[0] ^ data[4] ^ data[6] ^ data[8] ^ data[12] ^ data[17] ^ data[18] ^ data[19] ^ data[20] ^ data[25] ^ data[27] ^ data[28] ^ data[33] ^ data[36] ^ data[39] ^ data[42] ^ data[43] ^ data[45] ^ data[46] ^ data[48] ^ data[50] ^ data[51] ^ data[52] ^ data[53] ^ data[54] ^ data[55] ^ data[58] ^ data[59] ^ data[63];
    assign crcOut[27] = crcIn[4] ^ crcIn[6] ^ crcIn[7] ^ crcIn[9] ^ crcIn[11] ^ crcIn[12] ^ crcIn[14] ^ crcIn[15] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[27] ^ crcIn[28] ^ crcIn[30] ^ crcIn[34] ^ crcIn[36] ^ crcIn[37] ^ crcIn[38] ^ crcIn[39] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[62] ^ data[4] ^ data[6] ^ data[7] ^ data[9] ^ data[11] ^ data[12] ^ data[14] ^ data[15] ^ data[19] ^ data[20] ^ data[21] ^ data[22] ^ data[23] ^ data[27] ^ data[28] ^ data[30] ^ data[34] ^ data[36] ^ data[37] ^ data[38] ^ data[39] ^ data[44] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[50] ^ data[52] ^ data[53] ^ data[54] ^ data[57] ^ data[58] ^ data[59] ^ data[62];
    assign crcOut[28] = crcIn[5] ^ crcIn[7] ^ crcIn[8] ^ crcIn[10] ^ crcIn[12] ^ crcIn[13] ^ crcIn[15] ^ crcIn[16] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[28] ^ crcIn[29] ^ crcIn[31] ^ crcIn[35] ^ crcIn[37] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[51] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[63] ^ data[5] ^ data[7] ^ data[8] ^ data[10] ^ data[12] ^ data[13] ^ data[15] ^ data[16] ^ data[20] ^ data[21] ^ data[22] ^ data[23] ^ data[24] ^ data[28] ^ data[29] ^ data[31] ^ data[35] ^ data[37] ^ data[38] ^ data[39] ^ data[40] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[55] ^ data[58] ^ data[59] ^ data[60] ^ data[63];
    assign crcOut[29] = crcIn[1] ^ crcIn[4] ^ crcIn[5] ^ crcIn[8] ^ crcIn[9] ^ crcIn[12] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[21] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[32] ^ crcIn[41] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[52] ^ crcIn[54] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[62] ^ data[1] ^ data[4] ^ data[5] ^ data[8] ^ data[9] ^ data[12] ^ data[15] ^ data[16] ^ data[17] ^ data[18] ^ data[21] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[32] ^ data[41] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[49] ^ data[52] ^ data[54] ^ data[57] ^ data[58] ^ data[59] ^ data[61] ^ data[62];
    assign crcOut[30] = crcIn[0] ^ crcIn[2] ^ crcIn[5] ^ crcIn[6] ^ crcIn[9] ^ crcIn[10] ^ crcIn[13] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[22] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[33] ^ crcIn[42] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[50] ^ crcIn[53] ^ crcIn[55] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[2] ^ data[5] ^ data[6] ^ data[9] ^ data[10] ^ data[13] ^ data[16] ^ data[17] ^ data[18] ^ data[19] ^ data[22] ^ data[25] ^ data[26] ^ data[27] ^ data[28] ^ data[33] ^ data[42] ^ data[44] ^ data[46] ^ data[47] ^ data[48] ^ data[50] ^ data[53] ^ data[55] ^ data[58] ^ data[59] ^ data[60] ^ data[62] ^ data[63];
    assign crcOut[31] = crcIn[0] ^ crcIn[3] ^ crcIn[4] ^ crcIn[5] ^ crcIn[7] ^ crcIn[10] ^ crcIn[12] ^ crcIn[13] ^ crcIn[15] ^ crcIn[17] ^ crcIn[19] ^ crcIn[20] ^ crcIn[22] ^ crcIn[28] ^ crcIn[30] ^ crcIn[34] ^ crcIn[36] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[47] ^ crcIn[49] ^ crcIn[50] ^ crcIn[54] ^ crcIn[55] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[3] ^ data[4] ^ data[5] ^ data[7] ^ data[10] ^ data[12] ^ data[13] ^ data[15] ^ data[17] ^ data[19] ^ data[20] ^ data[22] ^ data[28] ^ data[30] ^ data[34] ^ data[36] ^ data[38] ^ data[39] ^ data[40] ^ data[47] ^ data[49] ^ data[50] ^ data[54] ^ data[55] ^ data[57] ^ data[58] ^ data[59] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[32] = crcIn[0] ^ crcIn[8] ^ crcIn[12] ^ crcIn[15] ^ crcIn[16] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[26] ^ crcIn[27] ^ crcIn[30] ^ crcIn[31] ^ crcIn[35] ^ crcIn[36] ^ crcIn[37] ^ crcIn[38] ^ crcIn[41] ^ crcIn[43] ^ crcIn[45] ^ crcIn[57] ^ crcIn[59] ^ crcIn[63] ^ data[0] ^ data[8] ^ data[12] ^ data[15] ^ data[16] ^ data[20] ^ data[21] ^ data[22] ^ data[26] ^ data[27] ^ data[30] ^ data[31] ^ data[35] ^ data[36] ^ data[37] ^ data[38] ^ data[41] ^ data[43] ^ data[45] ^ data[57] ^ data[59] ^ data[63];
    assign crcOut[33] = crcIn[0] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[9] ^ crcIn[11] ^ crcIn[12] ^ crcIn[14] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[21] ^ crcIn[26] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[37] ^ crcIn[40] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[50] ^ crcIn[51] ^ crcIn[55] ^ crcIn[56] ^ crcIn[57] ^ crcIn[62] ^ data[0] ^ data[4] ^ data[5] ^ data[6] ^ data[9] ^ data[11] ^ data[12] ^ data[14] ^ data[15] ^ data[16] ^ data[17] ^ data[18] ^ data[21] ^ data[26] ^ data[28] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[37] ^ data[40] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[48] ^ data[50] ^ data[51] ^ data[55] ^ data[56] ^ data[57] ^ data[62];
    assign crcOut[34] = crcIn[0] ^ crcIn[1] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[10] ^ crcIn[12] ^ crcIn[13] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[22] ^ crcIn[27] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[38] ^ crcIn[41] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[51] ^ crcIn[52] ^ crcIn[56] ^ crcIn[57] ^ crcIn[58] ^ crcIn[63] ^ data[0] ^ data[1] ^ data[5] ^ data[6] ^ data[7] ^ data[10] ^ data[12] ^ data[13] ^ data[15] ^ data[16] ^ data[17] ^ data[18] ^ data[19] ^ data[22] ^ data[27] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[33] ^ data[38] ^ data[41] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[47] ^ data[49] ^ data[51] ^ data[52] ^ data[56] ^ data[57] ^ data[58] ^ data[63];
    assign crcOut[35] = crcIn[0] ^ crcIn[2] ^ crcIn[4] ^ crcIn[5] ^ crcIn[7] ^ crcIn[8] ^ crcIn[12] ^ crcIn[15] ^ crcIn[16] ^ crcIn[17] ^ crcIn[19] ^ crcIn[20] ^ crcIn[22] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[36] ^ crcIn[38] ^ crcIn[40] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[55] ^ crcIn[56] ^ crcIn[59] ^ crcIn[60] ^ crcIn[62] ^ data[0] ^ data[2] ^ data[4] ^ data[5] ^ data[7] ^ data[8] ^ data[12] ^ data[15] ^ data[16] ^ data[17] ^ data[19] ^ data[20] ^ data[22] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[31] ^ data[32] ^ data[33] ^ data[34] ^ data[36] ^ data[38] ^ data[40] ^ data[42] ^ data[43] ^ data[44] ^ data[46] ^ data[47] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[56] ^ data[59] ^ data[60] ^ data[62];
    assign crcOut[36] = crcIn[1] ^ crcIn[3] ^ crcIn[5] ^ crcIn[6] ^ crcIn[8] ^ crcIn[9] ^ crcIn[13] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[20] ^ crcIn[21] ^ crcIn[23] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[37] ^ crcIn[39] ^ crcIn[41] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[47] ^ crcIn[48] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[57] ^ crcIn[60] ^ crcIn[61] ^ crcIn[63] ^ data[1] ^ data[3] ^ data[5] ^ data[6] ^ data[8] ^ data[9] ^ data[13] ^ data[16] ^ data[17] ^ data[18] ^ data[20] ^ data[21] ^ data[23] ^ data[27] ^ data[28] ^ data[29] ^ data[30] ^ data[32] ^ data[33] ^ data[34] ^ data[35] ^ data[37] ^ data[39] ^ data[41] ^ data[43] ^ data[44] ^ data[45] ^ data[47] ^ data[48] ^ data[52] ^ data[53] ^ data[54] ^ data[56] ^ data[57] ^ data[60] ^ data[61] ^ data[63];
    assign crcOut[37] = crcIn[0] ^ crcIn[1] ^ crcIn[2] ^ crcIn[5] ^ crcIn[7] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[15] ^ crcIn[17] ^ crcIn[19] ^ crcIn[21] ^ crcIn[23] ^ crcIn[24] ^ crcIn[26] ^ crcIn[27] ^ crcIn[28] ^ crcIn[31] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[39] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[46] ^ crcIn[49] ^ crcIn[50] ^ crcIn[51] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[60] ^ crcIn[61] ^ data[0] ^ data[1] ^ data[2] ^ data[5] ^ data[7] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[15] ^ data[17] ^ data[19] ^ data[21] ^ data[23] ^ data[24] ^ data[26] ^ data[27] ^ data[28] ^ data[31] ^ data[33] ^ data[34] ^ data[35] ^ data[39] ^ data[42] ^ data[43] ^ data[44] ^ data[46] ^ data[49] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[56] ^ data[60] ^ data[61];
    assign crcOut[38] = crcIn[1] ^ crcIn[2] ^ crcIn[3] ^ crcIn[6] ^ crcIn[8] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[16] ^ crcIn[18] ^ crcIn[20] ^ crcIn[22] ^ crcIn[24] ^ crcIn[25] ^ crcIn[27] ^ crcIn[28] ^ crcIn[29] ^ crcIn[32] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[40] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[47] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[54] ^ crcIn[55] ^ crcIn[57] ^ crcIn[61] ^ crcIn[62] ^ data[1] ^ data[2] ^ data[3] ^ data[6] ^ data[8] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[14] ^ data[16] ^ data[18] ^ data[20] ^ data[22] ^ data[24] ^ data[25] ^ data[27] ^ data[28] ^ data[29] ^ data[32] ^ data[34] ^ data[35] ^ data[36] ^ data[40] ^ data[43] ^ data[44] ^ data[45] ^ data[47] ^ data[50] ^ data[51] ^ data[52] ^ data[54] ^ data[55] ^ data[57] ^ data[61] ^ data[62];
    assign crcOut[39] = crcIn[0] ^ crcIn[2] ^ crcIn[3] ^ crcIn[4] ^ crcIn[7] ^ crcIn[9] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[15] ^ crcIn[17] ^ crcIn[19] ^ crcIn[21] ^ crcIn[23] ^ crcIn[25] ^ crcIn[26] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[33] ^ crcIn[35] ^ crcIn[36] ^ crcIn[37] ^ crcIn[41] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[55] ^ crcIn[56] ^ crcIn[58] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[2] ^ data[3] ^ data[4] ^ data[7] ^ data[9] ^ data[11] ^ data[12] ^ data[13] ^ data[14] ^ data[15] ^ data[17] ^ data[19] ^ data[21] ^ data[23] ^ data[25] ^ data[26] ^ data[28] ^ data[29] ^ data[30] ^ data[33] ^ data[35] ^ data[36] ^ data[37] ^ data[41] ^ data[44] ^ data[45] ^ data[46] ^ data[48] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[56] ^ data[58] ^ data[62] ^ data[63];
    assign crcOut[40] = crcIn[0] ^ crcIn[3] ^ crcIn[6] ^ crcIn[8] ^ crcIn[10] ^ crcIn[11] ^ crcIn[16] ^ crcIn[20] ^ crcIn[23] ^ crcIn[24] ^ crcIn[31] ^ crcIn[34] ^ crcIn[37] ^ crcIn[39] ^ crcIn[40] ^ crcIn[42] ^ crcIn[43] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[3] ^ data[6] ^ data[8] ^ data[10] ^ data[11] ^ data[16] ^ data[20] ^ data[23] ^ data[24] ^ data[31] ^ data[34] ^ data[37] ^ data[39] ^ data[40] ^ data[42] ^ data[43] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[50] ^ data[51] ^ data[52] ^ data[53] ^ data[54] ^ data[55] ^ data[58] ^ data[59] ^ data[60] ^ data[62] ^ data[63];
    assign crcOut[41] = crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[9] ^ crcIn[13] ^ crcIn[14] ^ crcIn[15] ^ crcIn[17] ^ crcIn[18] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[29] ^ crcIn[30] ^ crcIn[32] ^ crcIn[35] ^ crcIn[36] ^ crcIn[39] ^ crcIn[41] ^ crcIn[44] ^ crcIn[45] ^ crcIn[47] ^ crcIn[49] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[5] ^ data[6] ^ data[7] ^ data[9] ^ data[13] ^ data[14] ^ data[15] ^ data[17] ^ data[18] ^ data[21] ^ data[22] ^ data[23] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[29] ^ data[30] ^ data[32] ^ data[35] ^ data[36] ^ data[39] ^ data[41] ^ data[44] ^ data[45] ^ data[47] ^ data[49] ^ data[52] ^ data[53] ^ data[54] ^ data[57] ^ data[58] ^ data[59] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[42] = crcIn[0] ^ crcIn[1] ^ crcIn[4] ^ crcIn[5] ^ crcIn[7] ^ crcIn[8] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[16] ^ crcIn[19] ^ crcIn[24] ^ crcIn[25] ^ crcIn[28] ^ crcIn[29] ^ crcIn[31] ^ crcIn[33] ^ crcIn[37] ^ crcIn[38] ^ crcIn[39] ^ crcIn[42] ^ crcIn[43] ^ crcIn[46] ^ crcIn[51] ^ crcIn[53] ^ crcIn[54] ^ crcIn[56] ^ crcIn[57] ^ crcIn[59] ^ crcIn[63] ^ data[0] ^ data[1] ^ data[4] ^ data[5] ^ data[7] ^ data[8] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[16] ^ data[19] ^ data[24] ^ data[25] ^ data[28] ^ data[29] ^ data[31] ^ data[33] ^ data[37] ^ data[38] ^ data[39] ^ data[42] ^ data[43] ^ data[46] ^ data[51] ^ data[53] ^ data[54] ^ data[56] ^ data[57] ^ data[59] ^ data[63];
    assign crcOut[43] = crcIn[2] ^ crcIn[4] ^ crcIn[8] ^ crcIn[9] ^ crcIn[15] ^ crcIn[17] ^ crcIn[18] ^ crcIn[20] ^ crcIn[22] ^ crcIn[23] ^ crcIn[25] ^ crcIn[27] ^ crcIn[32] ^ crcIn[34] ^ crcIn[36] ^ crcIn[44] ^ crcIn[45] ^ crcIn[47] ^ crcIn[48] ^ crcIn[50] ^ crcIn[51] ^ crcIn[52] ^ crcIn[54] ^ crcIn[56] ^ crcIn[62] ^ data[2] ^ data[4] ^ data[8] ^ data[9] ^ data[15] ^ data[17] ^ data[18] ^ data[20] ^ data[22] ^ data[23] ^ data[25] ^ data[27] ^ data[32] ^ data[34] ^ data[36] ^ data[44] ^ data[45] ^ data[47] ^ data[48] ^ data[50] ^ data[51] ^ data[52] ^ data[54] ^ data[56] ^ data[62];
    assign crcOut[44] = crcIn[0] ^ crcIn[3] ^ crcIn[5] ^ crcIn[9] ^ crcIn[10] ^ crcIn[16] ^ crcIn[18] ^ crcIn[19] ^ crcIn[21] ^ crcIn[23] ^ crcIn[24] ^ crcIn[26] ^ crcIn[28] ^ crcIn[33] ^ crcIn[35] ^ crcIn[37] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[49] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[55] ^ crcIn[57] ^ crcIn[63] ^ data[0] ^ data[3] ^ data[5] ^ data[9] ^ data[10] ^ data[16] ^ data[18] ^ data[19] ^ data[21] ^ data[23] ^ data[24] ^ data[26] ^ data[28] ^ data[33] ^ data[35] ^ data[37] ^ data[45] ^ data[46] ^ data[48] ^ data[49] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[57] ^ data[63];
    assign crcOut[45] = crcIn[5] ^ crcIn[10] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[15] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[30] ^ crcIn[34] ^ crcIn[39] ^ crcIn[40] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[51] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[57] ^ crcIn[60] ^ crcIn[62] ^ data[5] ^ data[10] ^ data[12] ^ data[13] ^ data[14] ^ data[15] ^ data[17] ^ data[18] ^ data[19] ^ data[20] ^ data[23] ^ data[24] ^ data[25] ^ data[26] ^ data[30] ^ data[34] ^ data[39] ^ data[40] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[51] ^ data[52] ^ data[53] ^ data[54] ^ data[55] ^ data[57] ^ data[60] ^ data[62];
    assign crcOut[46] = crcIn[6] ^ crcIn[11] ^ crcIn[13] ^ crcIn[14] ^ crcIn[15] ^ crcIn[16] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[27] ^ crcIn[31] ^ crcIn[35] ^ crcIn[40] ^ crcIn[41] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[52] ^ crcIn[53] ^ crcIn[54] ^ crcIn[55] ^ crcIn[56] ^ crcIn[58] ^ crcIn[61] ^ crcIn[63] ^ data[6] ^ data[11] ^ data[13] ^ data[14] ^ data[15] ^ data[16] ^ data[18] ^ data[19] ^ data[20] ^ data[21] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[31] ^ data[35] ^ data[40] ^ data[41] ^ data[44] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[50] ^ data[52] ^ data[53] ^ data[54] ^ data[55] ^ data[56] ^ data[58] ^ data[61] ^ data[63];
    assign crcOut[47] = crcIn[0] ^ crcIn[1] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[11] ^ crcIn[13] ^ crcIn[16] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[23] ^ crcIn[25] ^ crcIn[28] ^ crcIn[29] ^ crcIn[30] ^ crcIn[32] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[47] ^ crcIn[49] ^ crcIn[53] ^ crcIn[54] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ data[0] ^ data[1] ^ data[4] ^ data[5] ^ data[6] ^ data[7] ^ data[11] ^ data[13] ^ data[16] ^ data[17] ^ data[18] ^ data[19] ^ data[20] ^ data[21] ^ data[23] ^ data[25] ^ data[28] ^ data[29] ^ data[30] ^ data[32] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[47] ^ data[49] ^ data[53] ^ data[54] ^ data[58] ^ data[59] ^ data[60];
    assign crcOut[48] = crcIn[1] ^ crcIn[2] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[12] ^ crcIn[14] ^ crcIn[17] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[24] ^ crcIn[26] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[33] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[48] ^ crcIn[50] ^ crcIn[54] ^ crcIn[55] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ data[1] ^ data[2] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[12] ^ data[14] ^ data[17] ^ data[18] ^ data[19] ^ data[20] ^ data[21] ^ data[22] ^ data[24] ^ data[26] ^ data[29] ^ data[30] ^ data[31] ^ data[33] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[48] ^ data[50] ^ data[54] ^ data[55] ^ data[59] ^ data[60] ^ data[61];
    assign crcOut[49] = crcIn[0] ^ crcIn[2] ^ crcIn[3] ^ crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[13] ^ crcIn[15] ^ crcIn[18] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[25] ^ crcIn[27] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[34] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[49] ^ crcIn[51] ^ crcIn[55] ^ crcIn[56] ^ crcIn[60] ^ crcIn[61] ^ crcIn[62] ^ data[0] ^ data[2] ^ data[3] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[13] ^ data[15] ^ data[18] ^ data[19] ^ data[20] ^ data[21] ^ data[22] ^ data[23] ^ data[25] ^ data[27] ^ data[30] ^ data[31] ^ data[32] ^ data[34] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[49] ^ data[51] ^ data[55] ^ data[56] ^ data[60] ^ data[61] ^ data[62];
    assign crcOut[50] = crcIn[0] ^ crcIn[1] ^ crcIn[3] ^ crcIn[4] ^ crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[14] ^ crcIn[16] ^ crcIn[19] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[26] ^ crcIn[28] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[35] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[50] ^ crcIn[52] ^ crcIn[56] ^ crcIn[57] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[1] ^ data[3] ^ data[4] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[14] ^ data[16] ^ data[19] ^ data[20] ^ data[21] ^ data[22] ^ data[23] ^ data[24] ^ data[26] ^ data[28] ^ data[31] ^ data[32] ^ data[33] ^ data[35] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[50] ^ data[52] ^ data[56] ^ data[57] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[51] = crcIn[0] ^ crcIn[2] ^ crcIn[6] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[17] ^ crcIn[18] ^ crcIn[20] ^ crcIn[21] ^ crcIn[24] ^ crcIn[25] ^ crcIn[26] ^ crcIn[30] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[42] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[50] ^ crcIn[53] ^ crcIn[55] ^ crcIn[56] ^ crcIn[60] ^ crcIn[63] ^ data[0] ^ data[2] ^ data[6] ^ data[8] ^ data[9] ^ data[10] ^ data[12] ^ data[13] ^ data[14] ^ data[17] ^ data[18] ^ data[20] ^ data[21] ^ data[24] ^ data[25] ^ data[26] ^ data[30] ^ data[32] ^ data[33] ^ data[34] ^ data[38] ^ data[39] ^ data[40] ^ data[42] ^ data[44] ^ data[46] ^ data[47] ^ data[48] ^ data[50] ^ data[53] ^ data[55] ^ data[56] ^ data[60] ^ data[63];
    assign crcOut[52] = crcIn[0] ^ crcIn[3] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[9] ^ crcIn[10] ^ crcIn[12] ^ crcIn[19] ^ crcIn[21] ^ crcIn[23] ^ crcIn[25] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[38] ^ crcIn[41] ^ crcIn[47] ^ crcIn[49] ^ crcIn[50] ^ crcIn[54] ^ crcIn[55] ^ crcIn[58] ^ crcIn[60] ^ crcIn[61] ^ crcIn[62] ^ data[0] ^ data[3] ^ data[4] ^ data[5] ^ data[6] ^ data[7] ^ data[9] ^ data[10] ^ data[12] ^ data[19] ^ data[21] ^ data[23] ^ data[25] ^ data[29] ^ data[30] ^ data[31] ^ data[33] ^ data[34] ^ data[35] ^ data[36] ^ data[38] ^ data[41] ^ data[47] ^ data[49] ^ data[50] ^ data[54] ^ data[55] ^ data[58] ^ data[60] ^ data[61] ^ data[62];
    assign crcOut[53] = crcIn[0] ^ crcIn[1] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[7] ^ crcIn[8] ^ crcIn[10] ^ crcIn[11] ^ crcIn[13] ^ crcIn[20] ^ crcIn[22] ^ crcIn[24] ^ crcIn[26] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[37] ^ crcIn[39] ^ crcIn[42] ^ crcIn[48] ^ crcIn[50] ^ crcIn[51] ^ crcIn[55] ^ crcIn[56] ^ crcIn[59] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[1] ^ data[4] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[10] ^ data[11] ^ data[13] ^ data[20] ^ data[22] ^ data[24] ^ data[26] ^ data[30] ^ data[31] ^ data[32] ^ data[34] ^ data[35] ^ data[36] ^ data[37] ^ data[39] ^ data[42] ^ data[48] ^ data[50] ^ data[51] ^ data[55] ^ data[56] ^ data[59] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[54] = crcIn[2] ^ crcIn[4] ^ crcIn[7] ^ crcIn[8] ^ crcIn[9] ^ crcIn[13] ^ crcIn[15] ^ crcIn[18] ^ crcIn[21] ^ crcIn[22] ^ crcIn[25] ^ crcIn[26] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[35] ^ crcIn[37] ^ crcIn[39] ^ crcIn[45] ^ crcIn[48] ^ crcIn[49] ^ crcIn[50] ^ crcIn[52] ^ crcIn[55] ^ crcIn[58] ^ crcIn[63] ^ data[2] ^ data[4] ^ data[7] ^ data[8] ^ data[9] ^ data[13] ^ data[15] ^ data[18] ^ data[21] ^ data[22] ^ data[25] ^ data[26] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[33] ^ data[35] ^ data[37] ^ data[39] ^ data[45] ^ data[48] ^ data[49] ^ data[50] ^ data[52] ^ data[55] ^ data[58] ^ data[63];
    assign crcOut[55] = crcIn[0] ^ crcIn[1] ^ crcIn[3] ^ crcIn[4] ^ crcIn[6] ^ crcIn[8] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[15] ^ crcIn[16] ^ crcIn[18] ^ crcIn[19] ^ crcIn[29] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[39] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[49] ^ crcIn[53] ^ crcIn[55] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[62] ^ data[0] ^ data[1] ^ data[3] ^ data[4] ^ data[6] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[15] ^ data[16] ^ data[18] ^ data[19] ^ data[29] ^ data[31] ^ data[32] ^ data[33] ^ data[34] ^ data[39] ^ data[43] ^ data[45] ^ data[46] ^ data[48] ^ data[49] ^ data[53] ^ data[55] ^ data[57] ^ data[58] ^ data[59] ^ data[60] ^ data[62];
    assign crcOut[56] = crcIn[1] ^ crcIn[2] ^ crcIn[4] ^ crcIn[5] ^ crcIn[7] ^ crcIn[9] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[16] ^ crcIn[17] ^ crcIn[19] ^ crcIn[20] ^ crcIn[30] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[40] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[50] ^ crcIn[54] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ crcIn[63] ^ data[1] ^ data[2] ^ data[4] ^ data[5] ^ data[7] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[14] ^ data[16] ^ data[17] ^ data[19] ^ data[20] ^ data[30] ^ data[32] ^ data[33] ^ data[34] ^ data[35] ^ data[40] ^ data[44] ^ data[46] ^ data[47] ^ data[49] ^ data[50] ^ data[54] ^ data[56] ^ data[58] ^ data[59] ^ data[60] ^ data[61] ^ data[63];
    assign crcOut[57] = crcIn[0] ^ crcIn[1] ^ crcIn[2] ^ crcIn[3] ^ crcIn[4] ^ crcIn[8] ^ crcIn[10] ^ crcIn[17] ^ crcIn[20] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[26] ^ crcIn[27] ^ crcIn[29] ^ crcIn[30] ^ crcIn[31] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[38] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[43] ^ crcIn[47] ^ crcIn[56] ^ crcIn[58] ^ crcIn[59] ^ crcIn[61] ^ data[0] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[8] ^ data[10] ^ data[17] ^ data[20] ^ data[21] ^ data[22] ^ data[23] ^ data[26] ^ data[27] ^ data[29] ^ data[30] ^ data[31] ^ data[33] ^ data[34] ^ data[35] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[43] ^ data[47] ^ data[56] ^ data[58] ^ data[59] ^ data[61];
    assign crcOut[58] = crcIn[1] ^ crcIn[2] ^ crcIn[3] ^ crcIn[4] ^ crcIn[5] ^ crcIn[9] ^ crcIn[11] ^ crcIn[18] ^ crcIn[21] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[27] ^ crcIn[28] ^ crcIn[30] ^ crcIn[31] ^ crcIn[32] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[44] ^ crcIn[48] ^ crcIn[57] ^ crcIn[59] ^ crcIn[60] ^ crcIn[62] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[5] ^ data[9] ^ data[11] ^ data[18] ^ data[21] ^ data[22] ^ data[23] ^ data[24] ^ data[27] ^ data[28] ^ data[30] ^ data[31] ^ data[32] ^ data[34] ^ data[35] ^ data[36] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[44] ^ data[48] ^ data[57] ^ data[59] ^ data[60] ^ data[62];
    assign crcOut[59] = crcIn[0] ^ crcIn[2] ^ crcIn[3] ^ crcIn[4] ^ crcIn[5] ^ crcIn[6] ^ crcIn[10] ^ crcIn[12] ^ crcIn[19] ^ crcIn[22] ^ crcIn[23] ^ crcIn[24] ^ crcIn[25] ^ crcIn[28] ^ crcIn[29] ^ crcIn[31] ^ crcIn[32] ^ crcIn[33] ^ crcIn[35] ^ crcIn[36] ^ crcIn[37] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[45] ^ crcIn[49] ^ crcIn[58] ^ crcIn[60] ^ crcIn[61] ^ crcIn[63] ^ data[0] ^ data[2] ^ data[3] ^ data[4] ^ data[5] ^ data[6] ^ data[10] ^ data[12] ^ data[19] ^ data[22] ^ data[23] ^ data[24] ^ data[25] ^ data[28] ^ data[29] ^ data[31] ^ data[32] ^ data[33] ^ data[35] ^ data[36] ^ data[37] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[45] ^ data[49] ^ data[58] ^ data[60] ^ data[61] ^ data[63];
    assign crcOut[60] = crcIn[0] ^ crcIn[3] ^ crcIn[7] ^ crcIn[12] ^ crcIn[14] ^ crcIn[15] ^ crcIn[18] ^ crcIn[20] ^ crcIn[22] ^ crcIn[24] ^ crcIn[25] ^ crcIn[27] ^ crcIn[32] ^ crcIn[33] ^ crcIn[34] ^ crcIn[37] ^ crcIn[39] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[44] ^ crcIn[45] ^ crcIn[46] ^ crcIn[48] ^ crcIn[51] ^ crcIn[55] ^ crcIn[56] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ data[0] ^ data[3] ^ data[7] ^ data[12] ^ data[14] ^ data[15] ^ data[18] ^ data[20] ^ data[22] ^ data[24] ^ data[25] ^ data[27] ^ data[32] ^ data[33] ^ data[34] ^ data[37] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[44] ^ data[45] ^ data[46] ^ data[48] ^ data[51] ^ data[55] ^ data[56] ^ data[57] ^ data[58] ^ data[59] ^ data[60] ^ data[61];
    assign crcOut[61] = crcIn[1] ^ crcIn[4] ^ crcIn[8] ^ crcIn[13] ^ crcIn[15] ^ crcIn[16] ^ crcIn[19] ^ crcIn[21] ^ crcIn[23] ^ crcIn[25] ^ crcIn[26] ^ crcIn[28] ^ crcIn[33] ^ crcIn[34] ^ crcIn[35] ^ crcIn[38] ^ crcIn[40] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[45] ^ crcIn[46] ^ crcIn[47] ^ crcIn[49] ^ crcIn[52] ^ crcIn[56] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ crcIn[62] ^ data[1] ^ data[4] ^ data[8] ^ data[13] ^ data[15] ^ data[16] ^ data[19] ^ data[21] ^ data[23] ^ data[25] ^ data[26] ^ data[28] ^ data[33] ^ data[34] ^ data[35] ^ data[38] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[45] ^ data[46] ^ data[47] ^ data[49] ^ data[52] ^ data[56] ^ data[57] ^ data[58] ^ data[59] ^ data[60] ^ data[61] ^ data[62];
    assign crcOut[62] = crcIn[0] ^ crcIn[2] ^ crcIn[5] ^ crcIn[9] ^ crcIn[14] ^ crcIn[16] ^ crcIn[17] ^ crcIn[20] ^ crcIn[22] ^ crcIn[24] ^ crcIn[26] ^ crcIn[27] ^ crcIn[29] ^ crcIn[34] ^ crcIn[35] ^ crcIn[36] ^ crcIn[39] ^ crcIn[41] ^ crcIn[42] ^ crcIn[43] ^ crcIn[44] ^ crcIn[46] ^ crcIn[47] ^ crcIn[48] ^ crcIn[50] ^ crcIn[53] ^ crcIn[57] ^ crcIn[58] ^ crcIn[59] ^ crcIn[60] ^ crcIn[61] ^ crcIn[62] ^ crcIn[63] ^ data[0] ^ data[2] ^ data[5] ^ data[9] ^ data[14] ^ data[16] ^ data[17] ^ data[20] ^ data[22] ^ data[24] ^ data[26] ^ data[27] ^ data[29] ^ data[34] ^ data[35] ^ data[36] ^ data[39] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[46] ^ data[47] ^ data[48] ^ data[50] ^ data[53] ^ data[57] ^ data[58] ^ data[59] ^ data[60] ^ data[61] ^ data[62] ^ data[63];
    assign crcOut[63] = crcIn[0] ^ crcIn[3] ^ crcIn[4] ^ crcIn[5] ^ crcIn[10] ^ crcIn[11] ^ crcIn[12] ^ crcIn[13] ^ crcIn[14] ^ crcIn[17] ^ crcIn[21] ^ crcIn[22] ^ crcIn[25] ^ crcIn[26] ^ crcIn[28] ^ crcIn[29] ^ crcIn[35] ^ crcIn[37] ^ crcIn[38] ^ crcIn[39] ^ crcIn[42] ^ crcIn[44] ^ crcIn[47] ^ crcIn[49] ^ crcIn[50] ^ crcIn[54] ^ crcIn[55] ^ crcIn[56] ^ crcIn[57] ^ crcIn[59] ^ crcIn[61] ^ crcIn[63] ^ data[0] ^ data[3] ^ data[4] ^ data[5] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[14] ^ data[17] ^ data[21] ^ data[22] ^ data[25] ^ data[26] ^ data[28] ^ data[29] ^ data[35] ^ data[37] ^ data[38] ^ data[39] ^ data[42] ^ data[44] ^ data[47] ^ data[49] ^ data[50] ^ data[54] ^ data[55] ^ data[56] ^ data[57] ^ data[59] ^ data[61] ^ data[63];
endmodule