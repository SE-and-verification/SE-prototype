module FU(
  input   io_A,
  input   io_B,
  output  io_out
);
  wire  _T_2 = io_B; // @[FU.scala 48:29]
  wire  _T_7 = io_A; // @[FU.scala 54:25]
  wire  _T_8 = io_A; // @[FU.scala 54:36]
  wire  _T_11 = _T_8 & _T_2; // @[FU.scala 54:56]
  wire  _T_12 = _T_7 & _T_11; // @[Cat.scala 30:58]
  wire  _GEN_0 = io_A & _T_2 & _T_12; // @[FU.scala 49:41 51:14 54:14]
  wire  _GEN_1 = io_A & _T_2 & _GEN_0; // @[FU.scala 46:35 48:14]
  wire  _T_15 = io_B; // @[FU.scala 59:39]
  wire  _GEN_2 = io_A & io_B & (io_A & io_B); // @[FU.scala 64:43 66:16 69:16]
  wire  _GEN_3 = io_A & io_B & _GEN_2; // @[FU.scala 61:37 63:16]
  wire  _GEN_4 = _T_8 & _T_15 & _GEN_3; // @[FU.scala 57:20 59:16]
  wire  _GEN_5 = io_A & io_B & (io_A & io_B); // @[FU.scala 76:44 78:16 81:16]
  wire  _GEN_6 = io_A & io_B & _GEN_5; // @[FU.scala 73:39 75:16]
  wire  _GEN_7 = _T_8 & _T_15 & (io_A & io_B); // @[FU.scala 84:20 86:14 89:14]
  wire  _GEN_8 = io_A & io_B; // @[FU.scala 92:26 94:14 97:14]
  wire  _GEN_9 = _GEN_8 & io_A; // @[FU.scala 101:14 91:37]
  wire  _GEN_10 = _GEN_7 & _GEN_9; // @[FU.scala 83:35]
  wire  _GEN_11 = _GEN_6 & _GEN_10; // @[FU.scala 72:38]
  wire  _GEN_12 = _GEN_4 & _GEN_11; // @[FU.scala 56:36]
  wire  _GEN_13 = _GEN_1 & _GEN_12; // @[FU.scala 45:30]
  assign io_out = _GEN_13; // @[FU.scala 43:20]
endmodule
module SEOperation(
  input   io_op1_input,
  input   io_op2_input,
  output  io_result
);
  wire  fu_io_A; // @[SEOperation.scala 32:24]
  wire  fu_io_B; // @[SEOperation.scala 32:24]
  wire  fu_io_out; // @[SEOperation.scala 32:24]
  FU fu ( // @[SEOperation.scala 32:24]
    .io_A(fu_io_A),
    .io_B(fu_io_B),
    .io_out(fu_io_out)
  );
  assign io_result = fu_io_out; // @[SEOperation.scala 47:19]
  assign fu_io_A = io_op1_input; // @[SEOperation.scala 41:11]
  assign fu_io_B = io_op2_input; // @[SEOperation.scala 42:11]
endmodule
module AddRoundKey(
  input   io_state_in_2,
  input   io_roundKey_2,
  output  io_state_out_2
);
  assign io_state_out_2 = io_state_in_2 & io_roundKey_2; // @[AddRoundKey.scala 19:41]
endmodule
module InvCipherRound(
  input   io_state_in_2,
  input   io_roundKey_2
);
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_state_out_2(AddRoundKey_io_state_out_2)
  );
  assign AddRoundKey_io_state_in_2 = io_state_in_2 & 1'h1; // @[InvCipherRound.scala 28:26 29:37 32:37]
  assign AddRoundKey_io_roundKey_2 = io_roundKey_2 & 1'h1; // @[InvCipherRound.scala 28:26 30:37 33:37]
endmodule
module InvSubBytes(
  output  io_state_out_2
);
  wire  _GEN_542 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_572 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_542))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_602 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_572))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_632 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_602))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_662 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_632))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_692 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_662))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_722 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_692))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  wire  _GEN_752 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_722))))))))))))))))))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
  assign io_state_out_2 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_752)))))))))))))); // @[InvSubBytes.scala 36:{23,23}]
endmodule
module InvCipherRound_3(
  input   io_roundKey_2
);
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  InvSubBytes_io_state_out_2; // @[InvSubBytes.scala 43:84]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_state_out_2(AddRoundKey_io_state_out_2)
  );
  InvSubBytes InvSubBytes ( // @[InvSubBytes.scala 43:84]
    .io_state_out_2(InvSubBytes_io_state_out_2)
  );
  assign AddRoundKey_io_state_in_2 = InvSubBytes_io_state_out_2; // @[InvCipherRound.scala 83:35]
  assign AddRoundKey_io_roundKey_2 = io_roundKey_2 & 1'h1; // @[InvCipherRound.scala 73:26 75:37 78:37]
endmodule
module InvCipherRound_30(
);
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  InvSubBytes_io_state_out_2; // @[InvSubBytes.scala 43:84]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_state_out_2(AddRoundKey_io_state_out_2)
  );
  InvSubBytes InvSubBytes ( // @[InvSubBytes.scala 43:84]
    .io_state_out_2(InvSubBytes_io_state_out_2)
  );
  assign AddRoundKey_io_state_in_2 = InvSubBytes_io_state_out_2; // @[InvCipherRound.scala 58:35]
  assign AddRoundKey_io_roundKey_2 = 1'h1 & 1'h1; // @[InvCipherRound.scala 48:26 50:37 53:37]
endmodule
module AESDecrypt(
  input   io_input_op1_2,
  input   io_input_op2_2,
  input   io_input_cond_2,
  output  io_output_op1_0,
  output  io_output_op1_1,
  output  io_output_op1_2,
  output  io_output_op1_3,
  output  io_output_op1_4,
  output  io_output_op1_5,
  output  io_output_op1_6,
  output  io_output_op1_7,
  output  io_output_op1_8,
  output  io_output_op1_9,
  output  io_output_op1_10,
  output  io_output_op1_11,
  output  io_output_op1_12,
  output  io_output_op1_13,
  output  io_output_op1_14,
  output  io_output_op1_15,
  output  io_output_op2_0,
  output  io_output_op2_1,
  output  io_output_op2_2,
  output  io_output_op2_3,
  output  io_output_op2_4,
  output  io_output_op2_5,
  output  io_output_op2_6,
  output  io_output_op2_7,
  output  io_output_op2_8,
  output  io_output_op2_9,
  output  io_output_op2_10,
  output  io_output_op2_11,
  output  io_output_op2_12,
  output  io_output_op2_13,
  output  io_output_op2_14,
  output  io_output_op2_15
);
  wire  InvCipherRound_io_state_in_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_state_in_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_1_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_state_in_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_2_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_3_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_4_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_5_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_6_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_7_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_8_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_9_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_10_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_11_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_12_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_13_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_14_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_15_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_16_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_17_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_18_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_19_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_20_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_21_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_22_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_23_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_24_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_25_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_26_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_27_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_28_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  wire  InvCipherRound_29_io_roundKey_2; // @[InvCipherRound.scala 96:79]
  InvCipherRound InvCipherRound ( // @[InvCipherRound.scala 96:79]
    .io_state_in_2(InvCipherRound_io_state_in_2),
    .io_roundKey_2(InvCipherRound_io_roundKey_2)
  );
  InvCipherRound InvCipherRound_1 ( // @[InvCipherRound.scala 96:79]
    .io_state_in_2(InvCipherRound_1_io_state_in_2),
    .io_roundKey_2(InvCipherRound_1_io_roundKey_2)
  );
  InvCipherRound InvCipherRound_2 ( // @[InvCipherRound.scala 96:79]
    .io_state_in_2(InvCipherRound_2_io_state_in_2),
    .io_roundKey_2(InvCipherRound_2_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_3 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_3_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_4 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_4_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_5 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_5_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_6 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_6_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_7 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_7_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_8 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_8_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_9 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_9_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_10 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_10_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_11 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_11_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_12 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_12_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_13 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_13_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_14 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_14_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_15 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_15_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_16 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_16_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_17 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_17_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_18 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_18_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_19 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_19_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_20 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_20_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_21 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_21_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_22 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_22_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_23 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_23_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_24 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_24_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_25 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_25_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_26 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_26_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_27 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_27_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_28 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_28_io_roundKey_2)
  );
  InvCipherRound_3 InvCipherRound_29 ( // @[InvCipherRound.scala 96:79]
    .io_roundKey_2(InvCipherRound_29_io_roundKey_2)
  );
  InvCipherRound_30 InvCipherRound_30 ( // @[InvCipherRound.scala 96:79]
  );
  InvCipherRound_30 InvCipherRound_31 ( // @[InvCipherRound.scala 96:79]
  );
  InvCipherRound_30 InvCipherRound_32 ( // @[InvCipherRound.scala 96:79]
  );
  assign io_output_op1_0 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_1 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_2 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_3 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_4 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_5 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_6 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_7 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_8 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_9 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_10 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_11 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_12 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_13 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_14 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op1_15 = 1'h0; // @[AESDecrypt.scala 74:17]
  assign io_output_op2_0 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_1 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_2 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_3 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_4 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_5 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_6 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_7 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_8 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_9 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_10 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_11 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_12 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_13 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_14 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign io_output_op2_15 = 1'h0; // @[AESDecrypt.scala 75:17]
  assign InvCipherRound_io_state_in_2 = io_input_op1_2; // @[AESDecrypt.scala 43:36]
  assign InvCipherRound_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 44:36]
  assign InvCipherRound_1_io_state_in_2 = io_input_op2_2; // @[AESDecrypt.scala 47:36]
  assign InvCipherRound_1_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 48:36]
  assign InvCipherRound_2_io_state_in_2 = io_input_cond_2; // @[AESDecrypt.scala 51:36]
  assign InvCipherRound_2_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 52:36]
  assign InvCipherRound_3_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_4_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_5_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_6_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_7_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_8_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_9_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_10_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_11_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_12_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_13_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_14_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_15_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_16_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_17_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_18_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_19_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_20_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_21_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_22_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_23_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_24_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_25_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_26_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_27_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_28_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
  assign InvCipherRound_29_io_roundKey_2 = 1'h1; // @[AESDecrypt.scala 64:41]
endmodule
module SubBytes(
  output  io_state_out_0,
  output  io_state_out_5,
  output  io_state_out_10
);
  wire  _GEN_30 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_60 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_30))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_90 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_60))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_120 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_90))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_150 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_120))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_180 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_150))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_210 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_180))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_240 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_210))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1310 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1340 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1310))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1370 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1340))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1400 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1370))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1430 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1400))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1460 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1430))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1490 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1460))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_1520 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1490))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2590 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2620 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2590))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2650 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2620))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2680 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2650))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2710 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2680))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2740 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2710))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2770 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2740))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  wire  _GEN_2800 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_2770))))))))))))))))))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_0 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_240)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_5 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_1520)))))))))))))); // @[SubBytes.scala 35:{23,23}]
  assign io_state_out_10 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & _GEN_2800)))))))))))))); // @[SubBytes.scala 35:{23,23}]
endmodule
module ShiftRows(
  input   io_state_in_0,
  input   io_state_in_5,
  input   io_state_in_10,
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2
);
  assign io_state_out_0 = io_state_in_0; // @[ShiftRows.scala 13:19]
  assign io_state_out_1 = io_state_in_5; // @[ShiftRows.scala 14:19]
  assign io_state_out_2 = io_state_in_10; // @[ShiftRows.scala 15:19]
endmodule
module MixColumns(
  input   io_state_in_0,
  input   io_state_in_1,
  output  io_state_out_2
);
  wire  _GEN_1054 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1084 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1054))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1114 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1084))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1144 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1114))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1174 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1144))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1204 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1174))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1234 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1204))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1264 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1234))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{51,51}]
  wire  _GEN_1310 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & 1'h1))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1340 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1310))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1370 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1340))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1400 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1370))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1430 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1400))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1460 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1430))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1490 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1460))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1520 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1490))))))))))))))))))))))))))))); // @[MixColumns.scala 127:{75,75}]
  wire  _GEN_1535 = 1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & _GEN_1520)))))))))))))); // @[MixColumns.scala 127:{75,75}]
  assign io_state_out_2 = io_state_in_0 & io_state_in_1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1
     & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & (1'h1 & _GEN_1264))))))))))))))) & _GEN_1535; // @[MixColumns.scala 127:75]
endmodule
module CipherRound_1(
  input   clock,
  input   io_roundKey_2,
  output  io_state_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  SubBytes_io_state_out_0; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_5; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_10; // @[SubBytes.scala 41:81]
  wire  ShiftRows_io_state_in_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_5; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_10; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_1; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_2; // @[ShiftRows.scala 35:34]
  wire  MixColumns_io_state_in_0; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_in_1; // @[MixColumns.scala 153:61]
  wire  MixColumns_io_state_out_2; // @[MixColumns.scala 153:61]
  reg  r__2; // @[Reg.scala 15:16]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_state_out_2(AddRoundKey_io_state_out_2)
  );
  SubBytes SubBytes ( // @[SubBytes.scala 41:81]
    .io_state_out_0(SubBytes_io_state_out_0),
    .io_state_out_5(SubBytes_io_state_out_5),
    .io_state_out_10(SubBytes_io_state_out_10)
  );
  ShiftRows ShiftRows ( // @[ShiftRows.scala 35:34]
    .io_state_in_0(ShiftRows_io_state_in_0),
    .io_state_in_5(ShiftRows_io_state_in_5),
    .io_state_in_10(ShiftRows_io_state_in_10),
    .io_state_out_0(ShiftRows_io_state_out_0),
    .io_state_out_1(ShiftRows_io_state_out_1),
    .io_state_out_2(ShiftRows_io_state_out_2)
  );
  MixColumns MixColumns ( // @[MixColumns.scala 153:61]
    .io_state_in_0(MixColumns_io_state_in_0),
    .io_state_in_1(MixColumns_io_state_in_1),
    .io_state_out_2(MixColumns_io_state_out_2)
  );
  assign io_state_out_2 = r__2; // @[CipherRound.scala 88:18]
  assign AddRoundKey_io_state_in_2 = MixColumns_io_state_out_2; // @[CipherRound.scala 85:35]
  assign AddRoundKey_io_roundKey_2 = io_roundKey_2 & 1'h1; // @[CipherRound.scala 73:26 75:37 78:37]
  assign ShiftRows_io_state_in_0 = SubBytes_io_state_out_0; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_5 = SubBytes_io_state_out_5; // @[CipherRound.scala 81:33]
  assign ShiftRows_io_state_in_10 = SubBytes_io_state_out_10; // @[CipherRound.scala 81:33]
  assign MixColumns_io_state_in_0 = ShiftRows_io_state_out_0; // @[CipherRound.scala 83:34]
  assign MixColumns_io_state_in_1 = ShiftRows_io_state_out_1; // @[CipherRound.scala 83:34]
  always @(posedge clock) begin
    r__2 <= AddRoundKey_io_state_out_2; // @[Reg.scala 15:16 16:{19,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r__2 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CipherRound_10(
  output  io_state_out_0,
  output  io_state_out_1,
  output  io_state_out_2,
  output  io_state_out_3,
  output  io_state_out_4,
  output  io_state_out_5,
  output  io_state_out_6,
  output  io_state_out_7,
  output  io_state_out_8,
  output  io_state_out_9,
  output  io_state_out_10,
  output  io_state_out_11,
  output  io_state_out_12,
  output  io_state_out_13,
  output  io_state_out_14,
  output  io_state_out_15,
  output  io_output_valid
);
  wire  AddRoundKey_io_state_in_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_roundKey_2; // @[AddRoundKey.scala 25:62]
  wire  AddRoundKey_io_state_out_2; // @[AddRoundKey.scala 25:62]
  wire  SubBytes_io_state_out_0; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_5; // @[SubBytes.scala 41:81]
  wire  SubBytes_io_state_out_10; // @[SubBytes.scala 41:81]
  wire  ShiftRows_io_state_in_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_5; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_in_10; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_0; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_1; // @[ShiftRows.scala 35:34]
  wire  ShiftRows_io_state_out_2; // @[ShiftRows.scala 35:34]
  AddRoundKey AddRoundKey ( // @[AddRoundKey.scala 25:62]
    .io_state_in_2(AddRoundKey_io_state_in_2),
    .io_roundKey_2(AddRoundKey_io_roundKey_2),
    .io_state_out_2(AddRoundKey_io_state_out_2)
  );
  SubBytes SubBytes ( // @[SubBytes.scala 41:81]
    .io_state_out_0(SubBytes_io_state_out_0),
    .io_state_out_5(SubBytes_io_state_out_5),
    .io_state_out_10(SubBytes_io_state_out_10)
  );
  ShiftRows ShiftRows ( // @[ShiftRows.scala 35:34]
    .io_state_in_0(ShiftRows_io_state_in_0),
    .io_state_in_5(ShiftRows_io_state_in_5),
    .io_state_in_10(ShiftRows_io_state_in_10),
    .io_state_out_0(ShiftRows_io_state_out_0),
    .io_state_out_1(ShiftRows_io_state_out_1),
    .io_state_out_2(ShiftRows_io_state_out_2)
  );
  assign io_state_out_0 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_1 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_2 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_3 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_4 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_5 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_6 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_7 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_8 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_9 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_10 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_11 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_12 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_13 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_14 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_state_out_15 = 1'h1; // @[CipherRound.scala 61:18]
  assign io_output_valid = 1'h1; // @[CipherRound.scala 62:21]
  assign AddRoundKey_io_state_in_2 = ShiftRows_io_state_out_2; // @[CipherRound.scala 58:35]
  assign AddRoundKey_io_roundKey_2 = 1'h1 & 1'h1; // @[CipherRound.scala 48:26 50:37 53:37]
  assign ShiftRows_io_state_in_0 = SubBytes_io_state_out_0; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_5 = SubBytes_io_state_out_5; // @[CipherRound.scala 56:33]
  assign ShiftRows_io_state_in_10 = SubBytes_io_state_out_10; // @[CipherRound.scala 56:33]
endmodule
module AESEncrypt(
  input   clock,
  input   io_input_text_2,
  output  io_output_text_0,
  output  io_output_text_1,
  output  io_output_text_2,
  output  io_output_text_3,
  output  io_output_text_4,
  output  io_output_text_5,
  output  io_output_text_6,
  output  io_output_text_7,
  output  io_output_text_8,
  output  io_output_text_9,
  output  io_output_text_10,
  output  io_output_text_11,
  output  io_output_text_12,
  output  io_output_text_13,
  output  io_output_text_14,
  output  io_output_text_15,
  output  io_output_intermediate,
  output  io_output_valid
);
  wire  CipherRoundARK_io_state_in_2; // @[CipherRound.scala 95:84]
  wire  CipherRoundARK_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_1_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_2_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_3_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_4_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_5_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_6_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_7_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_clock; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_roundKey_2; // @[CipherRound.scala 95:84]
  wire  CipherRound_8_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_0; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_1; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_2; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_3; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_4; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_5; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_6; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_7; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_8; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_9; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_10; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_11; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_12; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_13; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_14; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_state_out_15; // @[CipherRound.scala 95:84]
  wire  CipherRoundNMC_io_output_valid; // @[CipherRound.scala 95:84]
  InvCipherRound CipherRoundARK ( // @[CipherRound.scala 95:84]
    .io_state_in_2(CipherRoundARK_io_state_in_2),
    .io_roundKey_2(CipherRoundARK_io_roundKey_2)
  );
  CipherRound_1 CipherRound ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_clock),
    .io_roundKey_2(CipherRound_io_roundKey_2),
    .io_state_out_2(CipherRound_io_state_out_2)
  );
  CipherRound_1 CipherRound_1 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_1_clock),
    .io_roundKey_2(CipherRound_1_io_roundKey_2),
    .io_state_out_2(CipherRound_1_io_state_out_2)
  );
  CipherRound_1 CipherRound_2 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_2_clock),
    .io_roundKey_2(CipherRound_2_io_roundKey_2),
    .io_state_out_2(CipherRound_2_io_state_out_2)
  );
  CipherRound_1 CipherRound_3 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_3_clock),
    .io_roundKey_2(CipherRound_3_io_roundKey_2),
    .io_state_out_2(CipherRound_3_io_state_out_2)
  );
  CipherRound_1 CipherRound_4 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_4_clock),
    .io_roundKey_2(CipherRound_4_io_roundKey_2),
    .io_state_out_2(CipherRound_4_io_state_out_2)
  );
  CipherRound_1 CipherRound_5 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_5_clock),
    .io_roundKey_2(CipherRound_5_io_roundKey_2),
    .io_state_out_2(CipherRound_5_io_state_out_2)
  );
  CipherRound_1 CipherRound_6 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_6_clock),
    .io_roundKey_2(CipherRound_6_io_roundKey_2),
    .io_state_out_2(CipherRound_6_io_state_out_2)
  );
  CipherRound_1 CipherRound_7 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_7_clock),
    .io_roundKey_2(CipherRound_7_io_roundKey_2),
    .io_state_out_2(CipherRound_7_io_state_out_2)
  );
  CipherRound_1 CipherRound_8 ( // @[CipherRound.scala 95:84]
    .clock(CipherRound_8_clock),
    .io_roundKey_2(CipherRound_8_io_roundKey_2),
    .io_state_out_2(CipherRound_8_io_state_out_2)
  );
  CipherRound_10 CipherRoundNMC ( // @[CipherRound.scala 95:84]
    .io_state_out_0(CipherRoundNMC_io_state_out_0),
    .io_state_out_1(CipherRoundNMC_io_state_out_1),
    .io_state_out_2(CipherRoundNMC_io_state_out_2),
    .io_state_out_3(CipherRoundNMC_io_state_out_3),
    .io_state_out_4(CipherRoundNMC_io_state_out_4),
    .io_state_out_5(CipherRoundNMC_io_state_out_5),
    .io_state_out_6(CipherRoundNMC_io_state_out_6),
    .io_state_out_7(CipherRoundNMC_io_state_out_7),
    .io_state_out_8(CipherRoundNMC_io_state_out_8),
    .io_state_out_9(CipherRoundNMC_io_state_out_9),
    .io_state_out_10(CipherRoundNMC_io_state_out_10),
    .io_state_out_11(CipherRoundNMC_io_state_out_11),
    .io_state_out_12(CipherRoundNMC_io_state_out_12),
    .io_state_out_13(CipherRoundNMC_io_state_out_13),
    .io_state_out_14(CipherRoundNMC_io_state_out_14),
    .io_state_out_15(CipherRoundNMC_io_state_out_15),
    .io_output_valid(CipherRoundNMC_io_output_valid)
  );
  assign io_output_text_0 = CipherRoundNMC_io_state_out_0; // @[AESEncrypt.scala 54:18]
  assign io_output_text_1 = CipherRoundNMC_io_state_out_1; // @[AESEncrypt.scala 54:18]
  assign io_output_text_2 = CipherRoundNMC_io_state_out_2; // @[AESEncrypt.scala 54:18]
  assign io_output_text_3 = CipherRoundNMC_io_state_out_3; // @[AESEncrypt.scala 54:18]
  assign io_output_text_4 = CipherRoundNMC_io_state_out_4; // @[AESEncrypt.scala 54:18]
  assign io_output_text_5 = CipherRoundNMC_io_state_out_5; // @[AESEncrypt.scala 54:18]
  assign io_output_text_6 = CipherRoundNMC_io_state_out_6; // @[AESEncrypt.scala 54:18]
  assign io_output_text_7 = CipherRoundNMC_io_state_out_7; // @[AESEncrypt.scala 54:18]
  assign io_output_text_8 = CipherRoundNMC_io_state_out_8; // @[AESEncrypt.scala 54:18]
  assign io_output_text_9 = CipherRoundNMC_io_state_out_9; // @[AESEncrypt.scala 54:18]
  assign io_output_text_10 = CipherRoundNMC_io_state_out_10; // @[AESEncrypt.scala 54:18]
  assign io_output_text_11 = CipherRoundNMC_io_state_out_11; // @[AESEncrypt.scala 54:18]
  assign io_output_text_12 = CipherRoundNMC_io_state_out_12; // @[AESEncrypt.scala 54:18]
  assign io_output_text_13 = CipherRoundNMC_io_state_out_13; // @[AESEncrypt.scala 54:18]
  assign io_output_text_14 = CipherRoundNMC_io_state_out_14; // @[AESEncrypt.scala 54:18]
  assign io_output_text_15 = CipherRoundNMC_io_state_out_15; // @[AESEncrypt.scala 54:18]
  assign io_output_intermediate = CipherRound_3_io_state_out_2; // @[AESEncrypt.scala 52:26]
  assign io_output_valid = CipherRoundNMC_io_output_valid; // @[AESEncrypt.scala 53:19]
  assign CipherRoundARK_io_state_in_2 = io_input_text_2; // @[AESEncrypt.scala 32:30]
  assign CipherRoundARK_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 33:30]
  assign CipherRound_clock = clock;
  assign CipherRound_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_1_clock = clock;
  assign CipherRound_1_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_2_clock = clock;
  assign CipherRound_2_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_3_clock = clock;
  assign CipherRound_3_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_4_clock = clock;
  assign CipherRound_4_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_5_clock = clock;
  assign CipherRound_5_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_6_clock = clock;
  assign CipherRound_6_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_7_clock = clock;
  assign CipherRound_7_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
  assign CipherRound_8_clock = clock;
  assign CipherRound_8_io_roundKey_2 = 1'h1; // @[AESEncrypt.scala 45:33]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19,
  output  io_out_20,
  output  io_out_21,
  output  io_out_22,
  output  io_out_23,
  output  io_out_24,
  output  io_out_25,
  output  io_out_26,
  output  io_out_27,
  output  io_out_28,
  output  io_out_29,
  output  io_out_30,
  output  io_out_31,
  output  io_out_32,
  output  io_out_33,
  output  io_out_34,
  output  io_out_35,
  output  io_out_36,
  output  io_out_37,
  output  io_out_38,
  output  io_out_39,
  output  io_out_40,
  output  io_out_41,
  output  io_out_42,
  output  io_out_43,
  output  io_out_44,
  output  io_out_45,
  output  io_out_46,
  output  io_out_47,
  output  io_out_48,
  output  io_out_49,
  output  io_out_50,
  output  io_out_51,
  output  io_out_52,
  output  io_out_53,
  output  io_out_54,
  output  io_out_55,
  output  io_out_56,
  output  io_out_57,
  output  io_out_58,
  output  io_out_59,
  output  io_out_60,
  output  io_out_61,
  output  io_out_62,
  output  io_out_63
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 47:50]
  reg  state_1; // @[PRNG.scala 47:50]
  reg  state_2; // @[PRNG.scala 47:50]
  reg  state_3; // @[PRNG.scala 47:50]
  reg  state_4; // @[PRNG.scala 47:50]
  reg  state_5; // @[PRNG.scala 47:50]
  reg  state_6; // @[PRNG.scala 47:50]
  reg  state_7; // @[PRNG.scala 47:50]
  reg  state_8; // @[PRNG.scala 47:50]
  reg  state_9; // @[PRNG.scala 47:50]
  reg  state_10; // @[PRNG.scala 47:50]
  reg  state_11; // @[PRNG.scala 47:50]
  reg  state_12; // @[PRNG.scala 47:50]
  reg  state_13; // @[PRNG.scala 47:50]
  reg  state_14; // @[PRNG.scala 47:50]
  reg  state_15; // @[PRNG.scala 47:50]
  reg  state_16; // @[PRNG.scala 47:50]
  reg  state_17; // @[PRNG.scala 47:50]
  reg  state_18; // @[PRNG.scala 47:50]
  reg  state_19; // @[PRNG.scala 47:50]
  reg  state_20; // @[PRNG.scala 47:50]
  reg  state_21; // @[PRNG.scala 47:50]
  reg  state_22; // @[PRNG.scala 47:50]
  reg  state_23; // @[PRNG.scala 47:50]
  reg  state_24; // @[PRNG.scala 47:50]
  reg  state_25; // @[PRNG.scala 47:50]
  reg  state_26; // @[PRNG.scala 47:50]
  reg  state_27; // @[PRNG.scala 47:50]
  reg  state_28; // @[PRNG.scala 47:50]
  reg  state_29; // @[PRNG.scala 47:50]
  reg  state_30; // @[PRNG.scala 47:50]
  reg  state_31; // @[PRNG.scala 47:50]
  reg  state_32; // @[PRNG.scala 47:50]
  reg  state_33; // @[PRNG.scala 47:50]
  reg  state_34; // @[PRNG.scala 47:50]
  reg  state_35; // @[PRNG.scala 47:50]
  reg  state_36; // @[PRNG.scala 47:50]
  reg  state_37; // @[PRNG.scala 47:50]
  reg  state_38; // @[PRNG.scala 47:50]
  reg  state_39; // @[PRNG.scala 47:50]
  reg  state_40; // @[PRNG.scala 47:50]
  reg  state_41; // @[PRNG.scala 47:50]
  reg  state_42; // @[PRNG.scala 47:50]
  reg  state_43; // @[PRNG.scala 47:50]
  reg  state_44; // @[PRNG.scala 47:50]
  reg  state_45; // @[PRNG.scala 47:50]
  reg  state_46; // @[PRNG.scala 47:50]
  reg  state_47; // @[PRNG.scala 47:50]
  reg  state_48; // @[PRNG.scala 47:50]
  reg  state_49; // @[PRNG.scala 47:50]
  reg  state_50; // @[PRNG.scala 47:50]
  reg  state_51; // @[PRNG.scala 47:50]
  reg  state_52; // @[PRNG.scala 47:50]
  reg  state_53; // @[PRNG.scala 47:50]
  reg  state_54; // @[PRNG.scala 47:50]
  reg  state_55; // @[PRNG.scala 47:50]
  reg  state_56; // @[PRNG.scala 47:50]
  reg  state_57; // @[PRNG.scala 47:50]
  reg  state_58; // @[PRNG.scala 47:50]
  reg  state_59; // @[PRNG.scala 47:50]
  reg  state_60; // @[PRNG.scala 47:50]
  reg  state_61; // @[PRNG.scala 47:50]
  reg  state_62; // @[PRNG.scala 47:50]
  reg  state_63; // @[PRNG.scala 47:50]
  wire  _T_2 = state_63 & state_62 & state_60 & state_59; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  assign io_out_4 = state_4; // @[PRNG.scala 69:10]
  assign io_out_5 = state_5; // @[PRNG.scala 69:10]
  assign io_out_6 = state_6; // @[PRNG.scala 69:10]
  assign io_out_7 = state_7; // @[PRNG.scala 69:10]
  assign io_out_8 = state_8; // @[PRNG.scala 69:10]
  assign io_out_9 = state_9; // @[PRNG.scala 69:10]
  assign io_out_10 = state_10; // @[PRNG.scala 69:10]
  assign io_out_11 = state_11; // @[PRNG.scala 69:10]
  assign io_out_12 = state_12; // @[PRNG.scala 69:10]
  assign io_out_13 = state_13; // @[PRNG.scala 69:10]
  assign io_out_14 = state_14; // @[PRNG.scala 69:10]
  assign io_out_15 = state_15; // @[PRNG.scala 69:10]
  assign io_out_16 = state_16; // @[PRNG.scala 69:10]
  assign io_out_17 = state_17; // @[PRNG.scala 69:10]
  assign io_out_18 = state_18; // @[PRNG.scala 69:10]
  assign io_out_19 = state_19; // @[PRNG.scala 69:10]
  assign io_out_20 = state_20; // @[PRNG.scala 69:10]
  assign io_out_21 = state_21; // @[PRNG.scala 69:10]
  assign io_out_22 = state_22; // @[PRNG.scala 69:10]
  assign io_out_23 = state_23; // @[PRNG.scala 69:10]
  assign io_out_24 = state_24; // @[PRNG.scala 69:10]
  assign io_out_25 = state_25; // @[PRNG.scala 69:10]
  assign io_out_26 = state_26; // @[PRNG.scala 69:10]
  assign io_out_27 = state_27; // @[PRNG.scala 69:10]
  assign io_out_28 = state_28; // @[PRNG.scala 69:10]
  assign io_out_29 = state_29; // @[PRNG.scala 69:10]
  assign io_out_30 = state_30; // @[PRNG.scala 69:10]
  assign io_out_31 = state_31; // @[PRNG.scala 69:10]
  assign io_out_32 = state_32; // @[PRNG.scala 69:10]
  assign io_out_33 = state_33; // @[PRNG.scala 69:10]
  assign io_out_34 = state_34; // @[PRNG.scala 69:10]
  assign io_out_35 = state_35; // @[PRNG.scala 69:10]
  assign io_out_36 = state_36; // @[PRNG.scala 69:10]
  assign io_out_37 = state_37; // @[PRNG.scala 69:10]
  assign io_out_38 = state_38; // @[PRNG.scala 69:10]
  assign io_out_39 = state_39; // @[PRNG.scala 69:10]
  assign io_out_40 = state_40; // @[PRNG.scala 69:10]
  assign io_out_41 = state_41; // @[PRNG.scala 69:10]
  assign io_out_42 = state_42; // @[PRNG.scala 69:10]
  assign io_out_43 = state_43; // @[PRNG.scala 69:10]
  assign io_out_44 = state_44; // @[PRNG.scala 69:10]
  assign io_out_45 = state_45; // @[PRNG.scala 69:10]
  assign io_out_46 = state_46; // @[PRNG.scala 69:10]
  assign io_out_47 = state_47; // @[PRNG.scala 69:10]
  assign io_out_48 = state_48; // @[PRNG.scala 69:10]
  assign io_out_49 = state_49; // @[PRNG.scala 69:10]
  assign io_out_50 = state_50; // @[PRNG.scala 69:10]
  assign io_out_51 = state_51; // @[PRNG.scala 69:10]
  assign io_out_52 = state_52; // @[PRNG.scala 69:10]
  assign io_out_53 = state_53; // @[PRNG.scala 69:10]
  assign io_out_54 = state_54; // @[PRNG.scala 69:10]
  assign io_out_55 = state_55; // @[PRNG.scala 69:10]
  assign io_out_56 = state_56; // @[PRNG.scala 69:10]
  assign io_out_57 = state_57; // @[PRNG.scala 69:10]
  assign io_out_58 = state_58; // @[PRNG.scala 69:10]
  assign io_out_59 = state_59; // @[PRNG.scala 69:10]
  assign io_out_60 = state_60; // @[PRNG.scala 69:10]
  assign io_out_61 = state_61; // @[PRNG.scala 69:10]
  assign io_out_62 = state_62; // @[PRNG.scala 69:10]
  assign io_out_63 = state_63; // @[PRNG.scala 69:10]
  always @(posedge clock) begin
    state_0 <= 1'h1 & _T_2; // @[PRNG.scala 47:{50,50}]
    state_1 <= reset & state_0; // @[PRNG.scala 47:{50,50}]
    state_2 <= reset & state_1; // @[PRNG.scala 47:{50,50}]
    state_3 <= 1'h1 & state_2; // @[PRNG.scala 47:{50,50}]
    state_4 <= 1'h1 & state_3; // @[PRNG.scala 47:{50,50}]
    state_5 <= 1'h1 & state_4; // @[PRNG.scala 47:{50,50}]
    state_6 <= 1'h1 & state_5; // @[PRNG.scala 47:{50,50}]
    state_7 <= reset & state_6; // @[PRNG.scala 47:{50,50}]
    state_8 <= reset & state_7; // @[PRNG.scala 47:{50,50}]
    state_9 <= reset & state_8; // @[PRNG.scala 47:{50,50}]
    state_10 <= reset & state_9; // @[PRNG.scala 47:{50,50}]
    state_11 <= reset & state_10; // @[PRNG.scala 47:{50,50}]
    state_12 <= reset & state_11; // @[PRNG.scala 47:{50,50}]
    state_13 <= reset & state_12; // @[PRNG.scala 47:{50,50}]
    state_14 <= reset & state_13; // @[PRNG.scala 47:{50,50}]
    state_15 <= 1'h1 & state_14; // @[PRNG.scala 47:{50,50}]
    state_16 <= reset & state_15; // @[PRNG.scala 47:{50,50}]
    state_17 <= 1'h1 & state_16; // @[PRNG.scala 47:{50,50}]
    state_18 <= reset & state_17; // @[PRNG.scala 47:{50,50}]
    state_19 <= 1'h1 & state_18; // @[PRNG.scala 47:{50,50}]
    state_20 <= reset & state_19; // @[PRNG.scala 47:{50,50}]
    state_21 <= reset & state_20; // @[PRNG.scala 47:{50,50}]
    state_22 <= reset & state_21; // @[PRNG.scala 47:{50,50}]
    state_23 <= reset & state_22; // @[PRNG.scala 47:{50,50}]
    state_24 <= 1'h1 & state_23; // @[PRNG.scala 47:{50,50}]
    state_25 <= 1'h1 & state_24; // @[PRNG.scala 47:{50,50}]
    state_26 <= reset & state_25; // @[PRNG.scala 47:{50,50}]
    state_27 <= 1'h1 & state_26; // @[PRNG.scala 47:{50,50}]
    state_28 <= reset & state_27; // @[PRNG.scala 47:{50,50}]
    state_29 <= 1'h1 & state_28; // @[PRNG.scala 47:{50,50}]
    state_30 <= 1'h1 & state_29; // @[PRNG.scala 47:{50,50}]
    state_31 <= 1'h1 & state_30; // @[PRNG.scala 47:{50,50}]
    state_32 <= 1'h1 & state_31; // @[PRNG.scala 47:{50,50}]
    state_33 <= reset & state_32; // @[PRNG.scala 47:{50,50}]
    state_34 <= reset & state_33; // @[PRNG.scala 47:{50,50}]
    state_35 <= reset & state_34; // @[PRNG.scala 47:{50,50}]
    state_36 <= reset & state_35; // @[PRNG.scala 47:{50,50}]
    state_37 <= 1'h1 & state_36; // @[PRNG.scala 47:{50,50}]
    state_38 <= 1'h1 & state_37; // @[PRNG.scala 47:{50,50}]
    state_39 <= 1'h1 & state_38; // @[PRNG.scala 47:{50,50}]
    state_40 <= reset & state_39; // @[PRNG.scala 47:{50,50}]
    state_41 <= reset & state_40; // @[PRNG.scala 47:{50,50}]
    state_42 <= reset & state_41; // @[PRNG.scala 47:{50,50}]
    state_43 <= reset & state_42; // @[PRNG.scala 47:{50,50}]
    state_44 <= 1'h1 & state_43; // @[PRNG.scala 47:{50,50}]
    state_45 <= reset & state_44; // @[PRNG.scala 47:{50,50}]
    state_46 <= 1'h1 & state_45; // @[PRNG.scala 47:{50,50}]
    state_47 <= 1'h1 & state_46; // @[PRNG.scala 47:{50,50}]
    state_48 <= reset & state_47; // @[PRNG.scala 47:{50,50}]
    state_49 <= 1'h1 & state_48; // @[PRNG.scala 47:{50,50}]
    state_50 <= 1'h1 & state_49; // @[PRNG.scala 47:{50,50}]
    state_51 <= reset & state_50; // @[PRNG.scala 47:{50,50}]
    state_52 <= 1'h1 & state_51; // @[PRNG.scala 47:{50,50}]
    state_53 <= 1'h1 & state_52; // @[PRNG.scala 47:{50,50}]
    state_54 <= reset & state_53; // @[PRNG.scala 47:{50,50}]
    state_55 <= reset & state_54; // @[PRNG.scala 47:{50,50}]
    state_56 <= reset & state_55; // @[PRNG.scala 47:{50,50}]
    state_57 <= 1'h1 & state_56; // @[PRNG.scala 47:{50,50}]
    state_58 <= reset & state_57; // @[PRNG.scala 47:{50,50}]
    state_59 <= reset & state_58; // @[PRNG.scala 47:{50,50}]
    state_60 <= reset & state_59; // @[PRNG.scala 47:{50,50}]
    state_61 <= 1'h1 & state_60; // @[PRNG.scala 47:{50,50}]
    state_62 <= 1'h1 & state_61; // @[PRNG.scala 47:{50,50}]
    state_63 <= reset & state_62; // @[PRNG.scala 47:{50,50}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  state_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  state_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  state_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  state_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  state_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  state_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  state_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  state_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  state_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  state_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  state_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  state_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  state_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  state_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  state_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  state_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  state_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  state_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  state_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  state_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  state_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  state_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  state_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  state_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  state_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  state_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  state_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  state_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  state_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  state_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  state_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  state_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  state_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  state_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  state_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  state_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  state_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  state_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  state_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  state_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  state_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  state_63 = _RAND_63[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SE(
  input   clock,
  input   reset,
  input   io_in_inst,
  input   io_in_op1,
  input   io_in_op2,
  input   io_in_cond,
  input   io_in_valid,
  output  io_in_ready,
  output  io_out_result,
  output  io_out_valid,
  input   io_out_ready,
  output  io_out_cntr,
  output  io_out_zero_cntr,
  output  io_out_mult_cntr,
  output  io_out_intermediate
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  seoperation_io_op1_input; // @[SE.scala 83:33]
  wire  seoperation_io_op2_input; // @[SE.scala 83:33]
  wire  seoperation_io_result; // @[SE.scala 83:33]
  wire  aes_invcipher_io_input_op1_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_op2_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_input_cond_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op1_15; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_0; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_1; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_2; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_3; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_4; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_5; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_6; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_7; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_8; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_9; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_10; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_11; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_12; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_13; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_14; // @[SE.scala 84:35]
  wire  aes_invcipher_io_output_op2_15; // @[SE.scala 84:35]
  wire  aes_cipher_clock; // @[SE.scala 85:32]
  wire  aes_cipher_io_input_text_2; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_0; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_1; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_2; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_3; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_4; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_5; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_6; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_7; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_8; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_9; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_10; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_11; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_12; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_13; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_14; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_text_15; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_intermediate; // @[SE.scala 85:32]
  wire  aes_cipher_io_output_valid; // @[SE.scala 85:32]
  wire  prng_clock; // @[PRNG.scala 82:22]
  wire  prng_reset; // @[PRNG.scala 82:22]
  wire  prng_io_out_0; // @[PRNG.scala 82:22]
  wire  prng_io_out_1; // @[PRNG.scala 82:22]
  wire  prng_io_out_2; // @[PRNG.scala 82:22]
  wire  prng_io_out_3; // @[PRNG.scala 82:22]
  wire  prng_io_out_4; // @[PRNG.scala 82:22]
  wire  prng_io_out_5; // @[PRNG.scala 82:22]
  wire  prng_io_out_6; // @[PRNG.scala 82:22]
  wire  prng_io_out_7; // @[PRNG.scala 82:22]
  wire  prng_io_out_8; // @[PRNG.scala 82:22]
  wire  prng_io_out_9; // @[PRNG.scala 82:22]
  wire  prng_io_out_10; // @[PRNG.scala 82:22]
  wire  prng_io_out_11; // @[PRNG.scala 82:22]
  wire  prng_io_out_12; // @[PRNG.scala 82:22]
  wire  prng_io_out_13; // @[PRNG.scala 82:22]
  wire  prng_io_out_14; // @[PRNG.scala 82:22]
  wire  prng_io_out_15; // @[PRNG.scala 82:22]
  wire  prng_io_out_16; // @[PRNG.scala 82:22]
  wire  prng_io_out_17; // @[PRNG.scala 82:22]
  wire  prng_io_out_18; // @[PRNG.scala 82:22]
  wire  prng_io_out_19; // @[PRNG.scala 82:22]
  wire  prng_io_out_20; // @[PRNG.scala 82:22]
  wire  prng_io_out_21; // @[PRNG.scala 82:22]
  wire  prng_io_out_22; // @[PRNG.scala 82:22]
  wire  prng_io_out_23; // @[PRNG.scala 82:22]
  wire  prng_io_out_24; // @[PRNG.scala 82:22]
  wire  prng_io_out_25; // @[PRNG.scala 82:22]
  wire  prng_io_out_26; // @[PRNG.scala 82:22]
  wire  prng_io_out_27; // @[PRNG.scala 82:22]
  wire  prng_io_out_28; // @[PRNG.scala 82:22]
  wire  prng_io_out_29; // @[PRNG.scala 82:22]
  wire  prng_io_out_30; // @[PRNG.scala 82:22]
  wire  prng_io_out_31; // @[PRNG.scala 82:22]
  wire  prng_io_out_32; // @[PRNG.scala 82:22]
  wire  prng_io_out_33; // @[PRNG.scala 82:22]
  wire  prng_io_out_34; // @[PRNG.scala 82:22]
  wire  prng_io_out_35; // @[PRNG.scala 82:22]
  wire  prng_io_out_36; // @[PRNG.scala 82:22]
  wire  prng_io_out_37; // @[PRNG.scala 82:22]
  wire  prng_io_out_38; // @[PRNG.scala 82:22]
  wire  prng_io_out_39; // @[PRNG.scala 82:22]
  wire  prng_io_out_40; // @[PRNG.scala 82:22]
  wire  prng_io_out_41; // @[PRNG.scala 82:22]
  wire  prng_io_out_42; // @[PRNG.scala 82:22]
  wire  prng_io_out_43; // @[PRNG.scala 82:22]
  wire  prng_io_out_44; // @[PRNG.scala 82:22]
  wire  prng_io_out_45; // @[PRNG.scala 82:22]
  wire  prng_io_out_46; // @[PRNG.scala 82:22]
  wire  prng_io_out_47; // @[PRNG.scala 82:22]
  wire  prng_io_out_48; // @[PRNG.scala 82:22]
  wire  prng_io_out_49; // @[PRNG.scala 82:22]
  wire  prng_io_out_50; // @[PRNG.scala 82:22]
  wire  prng_io_out_51; // @[PRNG.scala 82:22]
  wire  prng_io_out_52; // @[PRNG.scala 82:22]
  wire  prng_io_out_53; // @[PRNG.scala 82:22]
  wire  prng_io_out_54; // @[PRNG.scala 82:22]
  wire  prng_io_out_55; // @[PRNG.scala 82:22]
  wire  prng_io_out_56; // @[PRNG.scala 82:22]
  wire  prng_io_out_57; // @[PRNG.scala 82:22]
  wire  prng_io_out_58; // @[PRNG.scala 82:22]
  wire  prng_io_out_59; // @[PRNG.scala 82:22]
  wire  prng_io_out_60; // @[PRNG.scala 82:22]
  wire  prng_io_out_61; // @[PRNG.scala 82:22]
  wire  prng_io_out_62; // @[PRNG.scala 82:22]
  wire  prng_io_out_63; // @[PRNG.scala 82:22]
  reg  value; // @[Counter.scala 60:40]
  reg  zero_cntr; // @[SE.scala 63:32]
  reg  mult_cntr; // @[SE.scala 64:32]
  wire  _GEN_0 = 1'h1 & (value & 1'h1); // @[Counter.scala 76:15 86:{20,28}]
  wire  _GEN_1 = _GEN_0 & value; // @[SE.scala 67:24 Counter.scala 60:40]
  wire  _T_1 = io_out_valid & io_out_ready; // @[SE.scala 72:33]
  wire  _GEN_4 = 1'h1 & _GEN_1; // @[SE.scala 75:43 Counter.scala 97:11]
  reg  op1_buffer; // @[Reg.scala 15:16]
  reg  op2_buffer; // @[Reg.scala 15:16]
  reg  cond_buffer; // @[Reg.scala 15:16]
  reg  ready_for_input; // @[SE.scala 117:38]
  wire  _GEN_185 = _T_1 & ready_for_input; // @[SE.scala 123:49 124:33 117:38]
  wire  _GEN_186 = 1'h1 & _GEN_185; // @[SE.scala 121:41 122:33]
  reg  mid_op1_buffer; // @[Reg.scala 15:16]
  wire  op1_reverse_1 = aes_invcipher_io_output_op1_14; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_0 = aes_invcipher_io_output_op1_15; // @[SE.scala 154:31 158:32]
  wire  lo_lo_lo = op1_reverse_1 & op1_reverse_0; // @[SE.scala 169:38]
  wire  op1_reverse_3 = aes_invcipher_io_output_op1_12; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_2 = aes_invcipher_io_output_op1_13; // @[SE.scala 154:31 158:32]
  wire  lo_lo_hi = op1_reverse_3 & op1_reverse_2; // @[SE.scala 169:38]
  wire  lo_lo = lo_lo_hi & lo_lo_lo; // @[SE.scala 169:38]
  wire  op1_reverse_5 = aes_invcipher_io_output_op1_10; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_4 = aes_invcipher_io_output_op1_11; // @[SE.scala 154:31 158:32]
  wire  lo_hi_lo = op1_reverse_5 & op1_reverse_4; // @[SE.scala 169:38]
  wire  op1_reverse_7 = aes_invcipher_io_output_op1_8; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_6 = aes_invcipher_io_output_op1_9; // @[SE.scala 154:31 158:32]
  wire  lo_hi_hi = op1_reverse_7 & op1_reverse_6; // @[SE.scala 169:38]
  wire  lo_hi = lo_hi_hi & lo_hi_lo; // @[SE.scala 169:38]
  wire  lo = lo_hi & lo_lo; // @[SE.scala 169:38]
  wire  op1_reverse_9 = aes_invcipher_io_output_op1_6; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_8 = aes_invcipher_io_output_op1_7; // @[SE.scala 154:31 158:32]
  wire  hi_lo_lo = op1_reverse_9 & op1_reverse_8; // @[SE.scala 169:38]
  wire  op1_reverse_11 = aes_invcipher_io_output_op1_4; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_10 = aes_invcipher_io_output_op1_5; // @[SE.scala 154:31 158:32]
  wire  hi_lo_hi = op1_reverse_11 & op1_reverse_10; // @[SE.scala 169:38]
  wire  hi_lo = hi_lo_hi & hi_lo_lo; // @[SE.scala 169:38]
  wire  op1_reverse_13 = aes_invcipher_io_output_op1_2; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_12 = aes_invcipher_io_output_op1_3; // @[SE.scala 154:31 158:32]
  wire  hi_hi_lo = op1_reverse_13 & op1_reverse_12; // @[SE.scala 169:38]
  wire  op1_reverse_15 = aes_invcipher_io_output_op1_0; // @[SE.scala 154:31 158:32]
  wire  op1_reverse_14 = aes_invcipher_io_output_op1_1; // @[SE.scala 154:31 158:32]
  wire  hi_hi_hi = op1_reverse_15 & op1_reverse_14; // @[SE.scala 169:38]
  wire  hi_hi = hi_hi_hi & hi_hi_lo; // @[SE.scala 169:38]
  wire  hi = hi_hi & hi_lo; // @[SE.scala 169:38]
  wire  op1_asUInt = hi & lo; // @[SE.scala 169:38]
  wire  op2_reverse_1 = aes_invcipher_io_output_op2_14; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_0 = aes_invcipher_io_output_op2_15; // @[SE.scala 155:31 159:32]
  wire  lo_lo_lo_1 = op2_reverse_1 & op2_reverse_0; // @[SE.scala 170:38]
  wire  op2_reverse_3 = aes_invcipher_io_output_op2_12; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_2 = aes_invcipher_io_output_op2_13; // @[SE.scala 155:31 159:32]
  wire  lo_lo_hi_1 = op2_reverse_3 & op2_reverse_2; // @[SE.scala 170:38]
  wire  lo_lo_1 = lo_lo_hi_1 & lo_lo_lo_1; // @[SE.scala 170:38]
  wire  op2_reverse_5 = aes_invcipher_io_output_op2_10; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_4 = aes_invcipher_io_output_op2_11; // @[SE.scala 155:31 159:32]
  wire  lo_hi_lo_1 = op2_reverse_5 & op2_reverse_4; // @[SE.scala 170:38]
  wire  op2_reverse_7 = aes_invcipher_io_output_op2_8; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_6 = aes_invcipher_io_output_op2_9; // @[SE.scala 155:31 159:32]
  wire  lo_hi_hi_1 = op2_reverse_7 & op2_reverse_6; // @[SE.scala 170:38]
  wire  lo_hi_1 = lo_hi_hi_1 & lo_hi_lo_1; // @[SE.scala 170:38]
  wire  lo_1 = lo_hi_1 & lo_lo_1; // @[SE.scala 170:38]
  wire  op2_reverse_9 = aes_invcipher_io_output_op2_6; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_8 = aes_invcipher_io_output_op2_7; // @[SE.scala 155:31 159:32]
  wire  hi_lo_lo_1 = op2_reverse_9 & op2_reverse_8; // @[SE.scala 170:38]
  wire  op2_reverse_11 = aes_invcipher_io_output_op2_4; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_10 = aes_invcipher_io_output_op2_5; // @[SE.scala 155:31 159:32]
  wire  hi_lo_hi_1 = op2_reverse_11 & op2_reverse_10; // @[SE.scala 170:38]
  wire  hi_lo_1 = hi_lo_hi_1 & hi_lo_lo_1; // @[SE.scala 170:38]
  wire  op2_reverse_13 = aes_invcipher_io_output_op2_2; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_12 = aes_invcipher_io_output_op2_3; // @[SE.scala 155:31 159:32]
  wire  hi_hi_lo_1 = op2_reverse_13 & op2_reverse_12; // @[SE.scala 170:38]
  wire  op2_reverse_15 = aes_invcipher_io_output_op2_0; // @[SE.scala 155:31 159:32]
  wire  op2_reverse_14 = aes_invcipher_io_output_op2_1; // @[SE.scala 155:31 159:32]
  wire  hi_hi_hi_1 = op2_reverse_15 & op2_reverse_14; // @[SE.scala 170:38]
  wire  hi_hi_1 = hi_hi_hi_1 & hi_hi_lo_1; // @[SE.scala 170:38]
  wire  hi_1 = hi_hi_1 & hi_lo_1; // @[SE.scala 170:38]
  wire  op2_asUInt = hi_1 & lo_1; // @[SE.scala 170:38]
  wire  _T_59 = mid_op1_buffer; // @[SE.scala 183:86]
  wire  _T_60 = op1_asUInt; // @[SE.scala 183:105]
  wire  lo_lo_lo_lo_lo = prng_io_out_1 & prng_io_out_0; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_lo_hi = prng_io_out_3 & prng_io_out_2; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_lo = lo_lo_lo_lo_hi & lo_lo_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_hi_lo = prng_io_out_5 & prng_io_out_4; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_hi_hi = prng_io_out_7 & prng_io_out_6; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_hi = lo_lo_lo_hi_hi & lo_lo_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_lo_3 = lo_lo_lo_hi & lo_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_lo_lo = prng_io_out_9 & prng_io_out_8; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_lo_hi = prng_io_out_11 & prng_io_out_10; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_lo = lo_lo_hi_lo_hi & lo_lo_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_hi_lo = prng_io_out_13 & prng_io_out_12; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_hi_hi = prng_io_out_15 & prng_io_out_14; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_hi = lo_lo_hi_hi_hi & lo_lo_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_hi_3 = lo_lo_hi_hi & lo_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_lo_3 = lo_lo_hi_3 & lo_lo_lo_3; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_lo_lo = prng_io_out_17 & prng_io_out_16; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_lo_hi = prng_io_out_19 & prng_io_out_18; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_lo = lo_hi_lo_lo_hi & lo_hi_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_hi_lo = prng_io_out_21 & prng_io_out_20; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_hi_hi = prng_io_out_23 & prng_io_out_22; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_hi = lo_hi_lo_hi_hi & lo_hi_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_lo_3 = lo_hi_lo_hi & lo_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_lo_lo = prng_io_out_25 & prng_io_out_24; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_lo_hi = prng_io_out_27 & prng_io_out_26; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_lo = lo_hi_hi_lo_hi & lo_hi_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_hi_lo = prng_io_out_29 & prng_io_out_28; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_hi_hi = prng_io_out_31 & prng_io_out_30; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_hi = lo_hi_hi_hi_hi & lo_hi_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_hi_3 = lo_hi_hi_hi & lo_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  lo_hi_3 = lo_hi_hi_3 & lo_hi_lo_3; // @[PRNG.scala 86:17]
  wire  lo_3 = lo_hi_3 & lo_lo_3; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_lo_lo = prng_io_out_33 & prng_io_out_32; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_lo_hi = prng_io_out_35 & prng_io_out_34; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_lo = hi_lo_lo_lo_hi & hi_lo_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_hi_lo = prng_io_out_37 & prng_io_out_36; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_hi_hi = prng_io_out_39 & prng_io_out_38; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_hi = hi_lo_lo_hi_hi & hi_lo_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_lo_3 = hi_lo_lo_hi & hi_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_lo_lo = prng_io_out_41 & prng_io_out_40; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_lo_hi = prng_io_out_43 & prng_io_out_42; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_lo = hi_lo_hi_lo_hi & hi_lo_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_hi_lo = prng_io_out_45 & prng_io_out_44; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_hi_hi = prng_io_out_47 & prng_io_out_46; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_hi = hi_lo_hi_hi_hi & hi_lo_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_hi_3 = hi_lo_hi_hi & hi_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_lo_3 = hi_lo_hi_3 & hi_lo_lo_3; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_lo_lo = prng_io_out_49 & prng_io_out_48; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_lo_hi = prng_io_out_51 & prng_io_out_50; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_lo = hi_hi_lo_lo_hi & hi_hi_lo_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_hi_lo = prng_io_out_53 & prng_io_out_52; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_hi_hi = prng_io_out_55 & prng_io_out_54; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_hi = hi_hi_lo_hi_hi & hi_hi_lo_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_lo_3 = hi_hi_lo_hi & hi_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_lo_lo = prng_io_out_57 & prng_io_out_56; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_lo_hi = prng_io_out_59 & prng_io_out_58; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_lo = hi_hi_hi_lo_hi & hi_hi_hi_lo_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_hi_lo = prng_io_out_61 & prng_io_out_60; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_hi_hi = prng_io_out_63 & prng_io_out_62; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_hi = hi_hi_hi_hi_hi & hi_hi_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_hi_3 = hi_hi_hi_hi & hi_hi_hi_lo; // @[PRNG.scala 86:17]
  wire  hi_hi_3 = hi_hi_hi_3 & hi_hi_lo_3; // @[PRNG.scala 86:17]
  wire  hi_3 = hi_hi_3 & hi_lo_3; // @[PRNG.scala 86:17]
  wire  bit64_randnum = hi_3 & lo_3; // @[PRNG.scala 86:17]
  wire  padded_result = seoperation_io_result & bit64_randnum; // @[Cat.scala 30:58]
  reg  result_buffer; // @[Reg.scala 15:16]
  wire  _GEN_190 = zero_cntr & 1'h1 & zero_cntr; // @[SE.scala 211:44 212:27 63:32]
  wire  _GEN_191 = mult_cntr & 1'h1 & mult_cntr; // @[SE.scala 214:56 215:27 64:32]
  wire  lo_lo_lo_4 = aes_cipher_io_output_text_1 & aes_cipher_io_output_text_0; // @[SE.scala 219:65]
  wire  lo_lo_hi_4 = aes_cipher_io_output_text_3 & aes_cipher_io_output_text_2; // @[SE.scala 219:65]
  wire  lo_lo_4 = lo_lo_hi_4 & lo_lo_lo_4; // @[SE.scala 219:65]
  wire  lo_hi_lo_4 = aes_cipher_io_output_text_5 & aes_cipher_io_output_text_4; // @[SE.scala 219:65]
  wire  lo_hi_hi_4 = aes_cipher_io_output_text_7 & aes_cipher_io_output_text_6; // @[SE.scala 219:65]
  wire  lo_hi_4 = lo_hi_hi_4 & lo_hi_lo_4; // @[SE.scala 219:65]
  wire  lo_4 = lo_hi_4 & lo_lo_4; // @[SE.scala 219:65]
  wire  hi_lo_lo_4 = aes_cipher_io_output_text_9 & aes_cipher_io_output_text_8; // @[SE.scala 219:65]
  wire  hi_lo_hi_4 = aes_cipher_io_output_text_11 & aes_cipher_io_output_text_10; // @[SE.scala 219:65]
  wire  hi_lo_4 = hi_lo_hi_4 & hi_lo_lo_4; // @[SE.scala 219:65]
  wire  hi_hi_lo_4 = aes_cipher_io_output_text_13 & aes_cipher_io_output_text_12; // @[SE.scala 219:65]
  wire  hi_hi_hi_4 = aes_cipher_io_output_text_15 & aes_cipher_io_output_text_14; // @[SE.scala 219:65]
  wire  hi_hi_4 = hi_hi_hi_4 & hi_hi_lo_4; // @[SE.scala 219:65]
  wire  hi_4 = hi_hi_4 & hi_lo_4; // @[SE.scala 219:65]
  wire  _T_89 = hi_4 & lo_4; // @[SE.scala 219:65]
  reg  output_buffer; // @[Reg.scala 15:16]
  reg  output_valid; // @[SE.scala 220:35]
  wire  _GEN_193 = 1'h1 & output_valid; // @[SE.scala 224:49 225:30 220:35]
  wire  _GEN_194 = aes_cipher_io_output_valid & _GEN_193; // @[SE.scala 222:41 223:30]
  SEOperation seoperation ( // @[SE.scala 83:33]
    .io_op1_input(seoperation_io_op1_input),
    .io_op2_input(seoperation_io_op2_input),
    .io_result(seoperation_io_result)
  );
  AESDecrypt aes_invcipher ( // @[SE.scala 84:35]
    .io_input_op1_2(aes_invcipher_io_input_op1_2),
    .io_input_op2_2(aes_invcipher_io_input_op2_2),
    .io_input_cond_2(aes_invcipher_io_input_cond_2),
    .io_output_op1_0(aes_invcipher_io_output_op1_0),
    .io_output_op1_1(aes_invcipher_io_output_op1_1),
    .io_output_op1_2(aes_invcipher_io_output_op1_2),
    .io_output_op1_3(aes_invcipher_io_output_op1_3),
    .io_output_op1_4(aes_invcipher_io_output_op1_4),
    .io_output_op1_5(aes_invcipher_io_output_op1_5),
    .io_output_op1_6(aes_invcipher_io_output_op1_6),
    .io_output_op1_7(aes_invcipher_io_output_op1_7),
    .io_output_op1_8(aes_invcipher_io_output_op1_8),
    .io_output_op1_9(aes_invcipher_io_output_op1_9),
    .io_output_op1_10(aes_invcipher_io_output_op1_10),
    .io_output_op1_11(aes_invcipher_io_output_op1_11),
    .io_output_op1_12(aes_invcipher_io_output_op1_12),
    .io_output_op1_13(aes_invcipher_io_output_op1_13),
    .io_output_op1_14(aes_invcipher_io_output_op1_14),
    .io_output_op1_15(aes_invcipher_io_output_op1_15),
    .io_output_op2_0(aes_invcipher_io_output_op2_0),
    .io_output_op2_1(aes_invcipher_io_output_op2_1),
    .io_output_op2_2(aes_invcipher_io_output_op2_2),
    .io_output_op2_3(aes_invcipher_io_output_op2_3),
    .io_output_op2_4(aes_invcipher_io_output_op2_4),
    .io_output_op2_5(aes_invcipher_io_output_op2_5),
    .io_output_op2_6(aes_invcipher_io_output_op2_6),
    .io_output_op2_7(aes_invcipher_io_output_op2_7),
    .io_output_op2_8(aes_invcipher_io_output_op2_8),
    .io_output_op2_9(aes_invcipher_io_output_op2_9),
    .io_output_op2_10(aes_invcipher_io_output_op2_10),
    .io_output_op2_11(aes_invcipher_io_output_op2_11),
    .io_output_op2_12(aes_invcipher_io_output_op2_12),
    .io_output_op2_13(aes_invcipher_io_output_op2_13),
    .io_output_op2_14(aes_invcipher_io_output_op2_14),
    .io_output_op2_15(aes_invcipher_io_output_op2_15)
  );
  AESEncrypt aes_cipher ( // @[SE.scala 85:32]
    .clock(aes_cipher_clock),
    .io_input_text_2(aes_cipher_io_input_text_2),
    .io_output_text_0(aes_cipher_io_output_text_0),
    .io_output_text_1(aes_cipher_io_output_text_1),
    .io_output_text_2(aes_cipher_io_output_text_2),
    .io_output_text_3(aes_cipher_io_output_text_3),
    .io_output_text_4(aes_cipher_io_output_text_4),
    .io_output_text_5(aes_cipher_io_output_text_5),
    .io_output_text_6(aes_cipher_io_output_text_6),
    .io_output_text_7(aes_cipher_io_output_text_7),
    .io_output_text_8(aes_cipher_io_output_text_8),
    .io_output_text_9(aes_cipher_io_output_text_9),
    .io_output_text_10(aes_cipher_io_output_text_10),
    .io_output_text_11(aes_cipher_io_output_text_11),
    .io_output_text_12(aes_cipher_io_output_text_12),
    .io_output_text_13(aes_cipher_io_output_text_13),
    .io_output_text_14(aes_cipher_io_output_text_14),
    .io_output_text_15(aes_cipher_io_output_text_15),
    .io_output_intermediate(aes_cipher_io_output_intermediate),
    .io_output_valid(aes_cipher_io_output_valid)
  );
  MaxPeriodFibonacciLFSR prng ( // @[PRNG.scala 82:22]
    .clock(prng_clock),
    .reset(prng_reset),
    .io_out_0(prng_io_out_0),
    .io_out_1(prng_io_out_1),
    .io_out_2(prng_io_out_2),
    .io_out_3(prng_io_out_3),
    .io_out_4(prng_io_out_4),
    .io_out_5(prng_io_out_5),
    .io_out_6(prng_io_out_6),
    .io_out_7(prng_io_out_7),
    .io_out_8(prng_io_out_8),
    .io_out_9(prng_io_out_9),
    .io_out_10(prng_io_out_10),
    .io_out_11(prng_io_out_11),
    .io_out_12(prng_io_out_12),
    .io_out_13(prng_io_out_13),
    .io_out_14(prng_io_out_14),
    .io_out_15(prng_io_out_15),
    .io_out_16(prng_io_out_16),
    .io_out_17(prng_io_out_17),
    .io_out_18(prng_io_out_18),
    .io_out_19(prng_io_out_19),
    .io_out_20(prng_io_out_20),
    .io_out_21(prng_io_out_21),
    .io_out_22(prng_io_out_22),
    .io_out_23(prng_io_out_23),
    .io_out_24(prng_io_out_24),
    .io_out_25(prng_io_out_25),
    .io_out_26(prng_io_out_26),
    .io_out_27(prng_io_out_27),
    .io_out_28(prng_io_out_28),
    .io_out_29(prng_io_out_29),
    .io_out_30(prng_io_out_30),
    .io_out_31(prng_io_out_31),
    .io_out_32(prng_io_out_32),
    .io_out_33(prng_io_out_33),
    .io_out_34(prng_io_out_34),
    .io_out_35(prng_io_out_35),
    .io_out_36(prng_io_out_36),
    .io_out_37(prng_io_out_37),
    .io_out_38(prng_io_out_38),
    .io_out_39(prng_io_out_39),
    .io_out_40(prng_io_out_40),
    .io_out_41(prng_io_out_41),
    .io_out_42(prng_io_out_42),
    .io_out_43(prng_io_out_43),
    .io_out_44(prng_io_out_44),
    .io_out_45(prng_io_out_45),
    .io_out_46(prng_io_out_46),
    .io_out_47(prng_io_out_47),
    .io_out_48(prng_io_out_48),
    .io_out_49(prng_io_out_49),
    .io_out_50(prng_io_out_50),
    .io_out_51(prng_io_out_51),
    .io_out_52(prng_io_out_52),
    .io_out_53(prng_io_out_53),
    .io_out_54(prng_io_out_54),
    .io_out_55(prng_io_out_55),
    .io_out_56(prng_io_out_56),
    .io_out_57(prng_io_out_57),
    .io_out_58(prng_io_out_58),
    .io_out_59(prng_io_out_59),
    .io_out_60(prng_io_out_60),
    .io_out_61(prng_io_out_61),
    .io_out_62(prng_io_out_62),
    .io_out_63(prng_io_out_63)
  );
  assign io_in_ready = ready_for_input; // @[SE.scala 118:21]
  assign io_out_result = output_buffer; // @[SE.scala 228:23]
  assign io_out_valid = output_valid; // @[SE.scala 227:22]
  assign io_out_cntr = value; // @[SE.scala 78:21]
  assign io_out_zero_cntr = zero_cntr; // @[SE.scala 65:26]
  assign io_out_mult_cntr = mult_cntr; // @[SE.scala 66:26]
  assign io_out_intermediate = aes_cipher_io_output_intermediate; // @[SE.scala 217:29]
  assign seoperation_io_op1_input = _T_59 & _T_60; // @[SE.scala 183:40]
  assign seoperation_io_op2_input = op2_asUInt; // @[SE.scala 184:47]
  assign aes_invcipher_io_input_op1_2 = op1_buffer; // @[SE.scala 146:58]
  assign aes_invcipher_io_input_op2_2 = op2_buffer; // @[SE.scala 147:58]
  assign aes_invcipher_io_input_cond_2 = cond_buffer; // @[SE.scala 148:60]
  assign aes_cipher_clock = clock;
  assign aes_cipher_io_input_text_2 = result_buffer; // @[SE.scala 203:47]
  assign prng_clock = clock;
  assign prng_reset = reset;
  always @(posedge clock) begin
    value <= 1'h1 & _GEN_4; // @[Counter.scala 60:{40,40}]
    zero_cntr <= 1'h1 & _GEN_190; // @[SE.scala 63:{32,32}]
    mult_cntr <= 1'h1 & _GEN_191; // @[SE.scala 64:{32,32}]
    op1_buffer <= io_in_op1 & op1_buffer; // @[Reg.scala 15:16 16:{19,23}]
    op2_buffer <= io_in_op2 & op2_buffer; // @[Reg.scala 15:16 16:{19,23}]
    cond_buffer <= io_in_cond & cond_buffer; // @[Reg.scala 15:16 16:{19,23}]
    ready_for_input <= reset & _GEN_186; // @[SE.scala 117:{38,38}]
    mid_op1_buffer <= op1_buffer & mid_op1_buffer; // @[Reg.scala 15:16 16:{19,23}]
    result_buffer <= padded_result & result_buffer; // @[Reg.scala 15:16 16:{19,23}]
    output_buffer <= _T_89 & output_buffer; // @[Reg.scala 15:16 16:{19,23}]
    output_valid <= 1'h1 & _GEN_194; // @[SE.scala 220:{35,35}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  zero_cntr = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mult_cntr = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  op1_buffer = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  op2_buffer = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cond_buffer = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ready_for_input = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  mid_op1_buffer = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  result_buffer = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_buffer = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_valid = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
